magic
tech sky130A
magscale 1 2
timestamp 1651159710
<< viali >>
rect 4261 37417 4295 37451
rect 9689 37417 9723 37451
rect 15945 37417 15979 37451
rect 7113 37349 7147 37383
rect 13185 37349 13219 37383
rect 2973 37281 3007 37315
rect 4905 37281 4939 37315
rect 14749 37281 14783 37315
rect 15485 37281 15519 37315
rect 17049 37281 17083 37315
rect 18429 37281 18463 37315
rect 22201 37281 22235 37315
rect 23673 37281 23707 37315
rect 30665 37281 30699 37315
rect 32505 37281 32539 37315
rect 33977 37281 34011 37315
rect 38025 37281 38059 37315
rect 1869 37213 1903 37247
rect 2789 37213 2823 37247
rect 4353 37213 4387 37247
rect 5825 37213 5859 37247
rect 6837 37213 6871 37247
rect 7665 37213 7699 37247
rect 9413 37213 9447 37247
rect 10241 37213 10275 37247
rect 11989 37213 12023 37247
rect 14565 37213 14599 37247
rect 15301 37213 15335 37247
rect 18153 37213 18187 37247
rect 19257 37213 19291 37247
rect 20177 37213 20211 37247
rect 20913 37213 20947 37247
rect 22385 37213 22419 37247
rect 22937 37213 22971 37247
rect 24409 37213 24443 37247
rect 25421 37213 25455 37247
rect 26157 37213 26191 37247
rect 26985 37213 27019 37247
rect 27905 37213 27939 37247
rect 28825 37213 28859 37247
rect 29561 37213 29595 37247
rect 30849 37213 30883 37247
rect 31585 37213 31619 37247
rect 32689 37213 32723 37247
rect 33517 37213 33551 37247
rect 34989 37213 35023 37247
rect 35725 37213 35759 37247
rect 36461 37213 36495 37247
rect 37289 37213 37323 37247
rect 5089 37145 5123 37179
rect 12909 37145 12943 37179
rect 17233 37145 17267 37179
rect 1961 37077 1995 37111
rect 5641 37077 5675 37111
rect 7849 37077 7883 37111
rect 10425 37077 10459 37111
rect 12081 37077 12115 37111
rect 19441 37077 19475 37111
rect 20361 37077 20395 37111
rect 21097 37077 21131 37111
rect 23121 37077 23155 37111
rect 24593 37077 24627 37111
rect 25605 37077 25639 37111
rect 26341 37077 26375 37111
rect 27169 37077 27203 37111
rect 28089 37077 28123 37111
rect 28733 37077 28767 37111
rect 29745 37077 29779 37111
rect 31401 37077 31435 37111
rect 33333 37077 33367 37111
rect 34805 37077 34839 37111
rect 35541 37077 35575 37111
rect 36277 37077 36311 37111
rect 37473 37077 37507 37111
rect 3433 36873 3467 36907
rect 4077 36873 4111 36907
rect 4813 36873 4847 36907
rect 5641 36873 5675 36907
rect 7297 36873 7331 36907
rect 8769 36873 8803 36907
rect 9413 36873 9447 36907
rect 10885 36873 10919 36907
rect 12173 36873 12207 36907
rect 13645 36873 13679 36907
rect 14473 36873 14507 36907
rect 15761 36873 15795 36907
rect 17877 36873 17911 36907
rect 18613 36873 18647 36907
rect 19533 36873 19567 36907
rect 20269 36873 20303 36907
rect 21097 36873 21131 36907
rect 22017 36873 22051 36907
rect 22753 36873 22787 36907
rect 24225 36873 24259 36907
rect 24961 36873 24995 36907
rect 25697 36873 25731 36907
rect 27169 36873 27203 36907
rect 27905 36873 27939 36907
rect 28549 36873 28583 36907
rect 29469 36873 29503 36907
rect 30205 36873 30239 36907
rect 31217 36873 31251 36907
rect 32321 36873 32355 36907
rect 33333 36873 33367 36907
rect 34437 36873 34471 36907
rect 35449 36873 35483 36907
rect 36553 36873 36587 36907
rect 1869 36805 1903 36839
rect 10057 36805 10091 36839
rect 12909 36805 12943 36839
rect 15025 36805 15059 36839
rect 17141 36805 17175 36839
rect 37289 36805 37323 36839
rect 37933 36805 37967 36839
rect 2789 36737 2823 36771
rect 3249 36737 3283 36771
rect 4261 36737 4295 36771
rect 4997 36737 5031 36771
rect 5457 36737 5491 36771
rect 6469 36737 6503 36771
rect 7113 36737 7147 36771
rect 8125 36737 8159 36771
rect 8585 36737 8619 36771
rect 9597 36737 9631 36771
rect 10701 36737 10735 36771
rect 12357 36737 12391 36771
rect 13829 36737 13863 36771
rect 14289 36737 14323 36771
rect 15945 36737 15979 36771
rect 18061 36737 18095 36771
rect 18797 36737 18831 36771
rect 19717 36737 19751 36771
rect 20453 36737 20487 36771
rect 20913 36737 20947 36771
rect 21833 36737 21867 36771
rect 22569 36737 22603 36771
rect 23581 36737 23615 36771
rect 24041 36737 24075 36771
rect 24777 36737 24811 36771
rect 25513 36737 25547 36771
rect 26433 36737 26467 36771
rect 26985 36737 27019 36771
rect 27721 36737 27755 36771
rect 28733 36737 28767 36771
rect 29285 36737 29319 36771
rect 30021 36737 30055 36771
rect 31033 36737 31067 36771
rect 32137 36737 32171 36771
rect 33149 36737 33183 36771
rect 34253 36737 34287 36771
rect 35265 36737 35299 36771
rect 36369 36737 36403 36771
rect 11529 36669 11563 36703
rect 2053 36601 2087 36635
rect 6653 36601 6687 36635
rect 7941 36601 7975 36635
rect 13093 36601 13127 36635
rect 38117 36601 38151 36635
rect 2605 36533 2639 36567
rect 17233 36533 17267 36567
rect 23397 36533 23431 36567
rect 26249 36533 26283 36567
rect 1501 36329 1535 36363
rect 2237 36329 2271 36363
rect 3065 36329 3099 36363
rect 4077 36329 4111 36363
rect 5365 36329 5399 36363
rect 6193 36329 6227 36363
rect 7297 36329 7331 36363
rect 7941 36329 7975 36363
rect 9045 36329 9079 36363
rect 10057 36329 10091 36363
rect 10793 36329 10827 36363
rect 11529 36329 11563 36363
rect 12541 36329 12575 36363
rect 14289 36329 14323 36363
rect 15209 36329 15243 36363
rect 15945 36329 15979 36363
rect 16773 36329 16807 36363
rect 17785 36329 17819 36363
rect 19349 36329 19383 36363
rect 20177 36329 20211 36363
rect 20821 36329 20855 36363
rect 21741 36329 21775 36363
rect 24501 36329 24535 36363
rect 25329 36329 25363 36363
rect 25973 36329 26007 36363
rect 26617 36329 26651 36363
rect 27261 36329 27295 36363
rect 28181 36329 28215 36363
rect 28641 36329 28675 36363
rect 29561 36329 29595 36363
rect 31861 36329 31895 36363
rect 34897 36329 34931 36363
rect 35449 36329 35483 36363
rect 13553 36261 13587 36295
rect 22753 36261 22787 36295
rect 23673 36261 23707 36295
rect 18429 36193 18463 36227
rect 30941 36193 30975 36227
rect 33333 36193 33367 36227
rect 36553 36193 36587 36227
rect 36829 36193 36863 36227
rect 37565 36193 37599 36227
rect 1685 36125 1719 36159
rect 2421 36125 2455 36159
rect 3249 36125 3283 36159
rect 4261 36125 4295 36159
rect 5549 36125 5583 36159
rect 6377 36125 6411 36159
rect 7481 36125 7515 36159
rect 8125 36125 8159 36159
rect 9229 36125 9263 36159
rect 10241 36125 10275 36159
rect 10977 36125 11011 36159
rect 11713 36125 11747 36159
rect 12725 36125 12759 36159
rect 13369 36125 13403 36159
rect 14105 36125 14139 36159
rect 15025 36125 15059 36159
rect 16129 36125 16163 36159
rect 16957 36125 16991 36159
rect 17969 36125 18003 36159
rect 19533 36125 19567 36159
rect 19993 36125 20027 36159
rect 20637 36125 20671 36159
rect 21925 36125 21959 36159
rect 24685 36125 24719 36159
rect 26457 36125 26491 36159
rect 27077 36125 27111 36159
rect 27997 36125 28031 36159
rect 28825 36125 28859 36159
rect 30205 36125 30239 36159
rect 31677 36125 31711 36159
rect 34713 36125 34747 36159
rect 37289 36125 37323 36159
rect 4905 36057 4939 36091
rect 22385 36057 22419 36091
rect 23305 36057 23339 36091
rect 30389 36057 30423 36091
rect 31125 36057 31159 36091
rect 32597 36057 32631 36091
rect 33517 36057 33551 36091
rect 34069 36057 34103 36091
rect 22845 35989 22879 36023
rect 23765 35989 23799 36023
rect 32505 35989 32539 36023
rect 1501 35785 1535 35819
rect 2697 35785 2731 35819
rect 3341 35785 3375 35819
rect 4537 35785 4571 35819
rect 5181 35785 5215 35819
rect 6653 35785 6687 35819
rect 8585 35785 8619 35819
rect 9781 35785 9815 35819
rect 10793 35785 10827 35819
rect 12265 35785 12299 35819
rect 14197 35785 14231 35819
rect 14841 35785 14875 35819
rect 15669 35785 15703 35819
rect 16681 35785 16715 35819
rect 17325 35785 17359 35819
rect 19717 35785 19751 35819
rect 22477 35785 22511 35819
rect 23213 35785 23247 35819
rect 23765 35785 23799 35819
rect 24317 35785 24351 35819
rect 26433 35785 26467 35819
rect 30481 35785 30515 35819
rect 31217 35785 31251 35819
rect 33425 35785 33459 35819
rect 35817 35785 35851 35819
rect 37289 35785 37323 35819
rect 29929 35717 29963 35751
rect 1685 35649 1719 35683
rect 2881 35649 2915 35683
rect 3525 35649 3559 35683
rect 6469 35649 6503 35683
rect 8769 35649 8803 35683
rect 9965 35649 9999 35683
rect 10977 35649 11011 35683
rect 11529 35649 11563 35683
rect 12449 35649 12483 35683
rect 14381 35649 14415 35683
rect 15025 35649 15059 35683
rect 15853 35649 15887 35683
rect 16865 35649 16899 35683
rect 17509 35649 17543 35683
rect 19533 35649 19567 35683
rect 23029 35649 23063 35683
rect 26249 35649 26283 35683
rect 26985 35649 27019 35683
rect 27537 35649 27571 35683
rect 28365 35649 28399 35683
rect 28825 35649 28859 35683
rect 30665 35649 30699 35683
rect 32781 35649 32815 35683
rect 33609 35649 33643 35683
rect 34069 35649 34103 35683
rect 35173 35649 35207 35683
rect 35633 35649 35667 35683
rect 36461 35649 36495 35683
rect 38025 35649 38059 35683
rect 2237 35581 2271 35615
rect 18981 35581 19015 35615
rect 7205 35513 7239 35547
rect 11713 35513 11747 35547
rect 27721 35513 27755 35547
rect 34253 35513 34287 35547
rect 34989 35513 35023 35547
rect 36645 35513 36679 35547
rect 3985 35445 4019 35479
rect 5733 35445 5767 35479
rect 8033 35445 8067 35479
rect 12909 35445 12943 35479
rect 13461 35445 13495 35479
rect 17969 35445 18003 35479
rect 20177 35445 20211 35479
rect 20729 35445 20763 35479
rect 21925 35445 21959 35479
rect 24869 35445 24903 35479
rect 25421 35445 25455 35479
rect 28181 35445 28215 35479
rect 32689 35445 32723 35479
rect 37933 35445 37967 35479
rect 1593 35241 1627 35275
rect 2145 35241 2179 35275
rect 6193 35241 6227 35275
rect 6745 35241 6779 35275
rect 7849 35241 7883 35275
rect 9965 35241 9999 35275
rect 10425 35241 10459 35275
rect 12173 35241 12207 35275
rect 12725 35241 12759 35275
rect 15301 35241 15335 35275
rect 17509 35241 17543 35275
rect 18061 35241 18095 35275
rect 18613 35241 18647 35275
rect 19257 35241 19291 35275
rect 20085 35241 20119 35275
rect 29561 35241 29595 35275
rect 33517 35241 33551 35275
rect 35357 35241 35391 35275
rect 38025 35241 38059 35275
rect 2697 35173 2731 35207
rect 15945 35173 15979 35207
rect 26341 35173 26375 35207
rect 30113 35105 30147 35139
rect 2881 35037 2915 35071
rect 10609 35037 10643 35071
rect 15117 35037 15151 35071
rect 15761 35037 15795 35071
rect 16405 35037 16439 35071
rect 30021 35037 30055 35071
rect 35541 35037 35575 35071
rect 36001 35037 36035 35071
rect 37841 35037 37875 35071
rect 13369 34969 13403 35003
rect 25973 34969 26007 35003
rect 31401 34969 31435 35003
rect 36268 34969 36302 35003
rect 3893 34901 3927 34935
rect 4445 34901 4479 34935
rect 4997 34901 5031 34935
rect 5549 34901 5583 34935
rect 7297 34901 7331 34935
rect 8953 34901 8987 34935
rect 11069 34901 11103 34935
rect 11713 34901 11747 34935
rect 14473 34901 14507 34935
rect 16957 34901 16991 34935
rect 20545 34901 20579 34935
rect 21097 34901 21131 34935
rect 22845 34901 22879 34935
rect 26433 34901 26467 34935
rect 29009 34901 29043 34935
rect 29929 34901 29963 34935
rect 30849 34901 30883 34935
rect 31953 34901 31987 34935
rect 32965 34901 32999 34935
rect 34069 34901 34103 34935
rect 34713 34901 34747 34935
rect 37381 34901 37415 34935
rect 2605 34697 2639 34731
rect 9229 34697 9263 34731
rect 12173 34697 12207 34731
rect 12909 34697 12943 34731
rect 15669 34697 15703 34731
rect 16957 34697 16991 34731
rect 23305 34697 23339 34731
rect 24225 34697 24259 34731
rect 36553 34697 36587 34731
rect 37381 34697 37415 34731
rect 38025 34697 38059 34731
rect 3617 34629 3651 34663
rect 6377 34629 6411 34663
rect 22845 34629 22879 34663
rect 23765 34629 23799 34663
rect 34805 34629 34839 34663
rect 4712 34561 4746 34595
rect 13921 34561 13955 34595
rect 14565 34561 14599 34595
rect 15117 34561 15151 34595
rect 18328 34561 18362 34595
rect 35265 34561 35299 34595
rect 36737 34561 36771 34595
rect 37841 34561 37875 34595
rect 3065 34493 3099 34527
rect 4445 34493 4479 34527
rect 9781 34493 9815 34527
rect 10701 34493 10735 34527
rect 11529 34493 11563 34527
rect 17509 34493 17543 34527
rect 18061 34493 18095 34527
rect 19993 34493 20027 34527
rect 20545 34493 20579 34527
rect 32965 34493 32999 34527
rect 33793 34493 33827 34527
rect 23121 34425 23155 34459
rect 24041 34425 24075 34459
rect 5825 34357 5859 34391
rect 19441 34357 19475 34391
rect 22385 34357 22419 34391
rect 36001 34357 36035 34391
rect 18061 34153 18095 34187
rect 31309 34153 31343 34187
rect 35909 34153 35943 34187
rect 36369 34153 36403 34187
rect 37197 34153 37231 34187
rect 37933 34153 37967 34187
rect 9413 33949 9447 33983
rect 31493 33949 31527 33983
rect 36553 33949 36587 33983
rect 37013 33949 37047 33983
rect 37749 33949 37783 33983
rect 9680 33881 9714 33915
rect 10793 33813 10827 33847
rect 11345 33813 11379 33847
rect 15945 33813 15979 33847
rect 17141 33813 17175 33847
rect 23673 33813 23707 33847
rect 33885 33813 33919 33847
rect 34713 33813 34747 33847
rect 35357 33813 35391 33847
rect 5273 33609 5307 33643
rect 10149 33609 10183 33643
rect 11621 33609 11655 33643
rect 18429 33609 18463 33643
rect 29377 33609 29411 33643
rect 36737 33609 36771 33643
rect 37381 33609 37415 33643
rect 38025 33609 38059 33643
rect 5457 33473 5491 33507
rect 10333 33473 10367 33507
rect 10609 33473 10643 33507
rect 11529 33473 11563 33507
rect 11805 33473 11839 33507
rect 18613 33473 18647 33507
rect 27537 33473 27571 33507
rect 29193 33473 29227 33507
rect 37841 33473 37875 33507
rect 5733 33405 5767 33439
rect 18889 33405 18923 33439
rect 27813 33405 27847 33439
rect 11805 33337 11839 33371
rect 12357 33337 12391 33371
rect 5641 33269 5675 33303
rect 10517 33269 10551 33303
rect 18797 33269 18831 33303
rect 35357 33269 35391 33303
rect 36185 33269 36219 33303
rect 19533 33065 19567 33099
rect 28457 32997 28491 33031
rect 19257 32861 19291 32895
rect 19349 32861 19383 32895
rect 28273 32861 28307 32895
rect 37841 32861 37875 32895
rect 38117 32861 38151 32895
rect 19533 32793 19567 32827
rect 19993 32725 20027 32759
rect 36277 32725 36311 32759
rect 36829 32725 36863 32759
rect 6837 32521 6871 32555
rect 26157 32521 26191 32555
rect 32137 32521 32171 32555
rect 38117 32453 38151 32487
rect 6745 32385 6779 32419
rect 6929 32385 6963 32419
rect 13645 32385 13679 32419
rect 14105 32385 14139 32419
rect 14372 32385 14406 32419
rect 25789 32385 25823 32419
rect 25973 32385 26007 32419
rect 32505 32385 32539 32419
rect 32597 32385 32631 32419
rect 32781 32317 32815 32351
rect 31493 32249 31527 32283
rect 7481 32181 7515 32215
rect 15485 32181 15519 32215
rect 25329 32181 25363 32215
rect 37565 32181 37599 32215
rect 26525 31977 26559 32011
rect 28365 31977 28399 32011
rect 25697 31773 25731 31807
rect 26157 31773 26191 31807
rect 26341 31773 26375 31807
rect 27445 31773 27479 31807
rect 27997 31773 28031 31807
rect 28181 31773 28215 31807
rect 34897 31433 34931 31467
rect 34713 31297 34747 31331
rect 36470 31297 36504 31331
rect 36737 31297 36771 31331
rect 37473 31297 37507 31331
rect 38117 31297 38151 31331
rect 35357 31093 35391 31127
rect 37933 31093 37967 31127
rect 27077 30889 27111 30923
rect 33057 30889 33091 30923
rect 35265 30889 35299 30923
rect 32873 30821 32907 30855
rect 27629 30753 27663 30787
rect 1869 30685 1903 30719
rect 3801 30685 3835 30719
rect 4813 30685 4847 30719
rect 4997 30685 5031 30719
rect 23673 30685 23707 30719
rect 27537 30685 27571 30719
rect 2136 30617 2170 30651
rect 23406 30617 23440 30651
rect 24501 30617 24535 30651
rect 32597 30617 32631 30651
rect 3249 30549 3283 30583
rect 4905 30549 4939 30583
rect 5549 30549 5583 30583
rect 22293 30549 22327 30583
rect 26617 30549 26651 30583
rect 27445 30549 27479 30583
rect 4997 30345 5031 30379
rect 12909 30345 12943 30379
rect 16037 30345 16071 30379
rect 22753 30345 22787 30379
rect 32413 30345 32447 30379
rect 32781 30345 32815 30379
rect 3617 30277 3651 30311
rect 5165 30277 5199 30311
rect 5365 30277 5399 30311
rect 6377 30277 6411 30311
rect 6745 30277 6779 30311
rect 8033 30277 8067 30311
rect 11529 30277 11563 30311
rect 11729 30277 11763 30311
rect 13001 30277 13035 30311
rect 14381 30277 14415 30311
rect 15485 30277 15519 30311
rect 19149 30277 19183 30311
rect 19349 30277 19383 30311
rect 20085 30277 20119 30311
rect 32229 30277 32263 30311
rect 1869 30209 1903 30243
rect 3801 30209 3835 30243
rect 6561 30209 6595 30243
rect 6653 30209 6687 30243
rect 6929 30209 6963 30243
rect 7849 30209 7883 30243
rect 12817 30209 12851 30243
rect 14565 30209 14599 30243
rect 14841 30209 14875 30243
rect 15393 30209 15427 30243
rect 15589 30209 15623 30243
rect 17233 30209 17267 30243
rect 18245 30209 18279 30243
rect 18337 30209 18371 30243
rect 18521 30209 18555 30243
rect 19993 30209 20027 30243
rect 20177 30209 20211 30243
rect 22569 30209 22603 30243
rect 32505 30209 32539 30243
rect 4077 30141 4111 30175
rect 14749 30141 14783 30175
rect 17509 30141 17543 30175
rect 19809 30141 19843 30175
rect 22293 30141 22327 30175
rect 32137 30141 32171 30175
rect 32597 30141 32631 30175
rect 2145 30073 2179 30107
rect 11897 30073 11931 30107
rect 12633 30073 12667 30107
rect 18981 30073 19015 30107
rect 22385 30073 22419 30107
rect 3985 30005 4019 30039
rect 5181 30005 5215 30039
rect 11713 30005 11747 30039
rect 13185 30005 13219 30039
rect 18521 30005 18555 30039
rect 19165 30005 19199 30039
rect 20361 30005 20395 30039
rect 31493 30005 31527 30039
rect 1593 29801 1627 29835
rect 32689 29801 32723 29835
rect 37933 29801 37967 29835
rect 9873 29733 9907 29767
rect 11345 29733 11379 29767
rect 32321 29665 32355 29699
rect 32413 29665 32447 29699
rect 11069 29597 11103 29631
rect 11161 29597 11195 29631
rect 25421 29597 25455 29631
rect 32229 29597 32263 29631
rect 32505 29597 32539 29631
rect 37473 29597 37507 29631
rect 38117 29597 38151 29631
rect 10057 29529 10091 29563
rect 11345 29529 11379 29563
rect 25237 29529 25271 29563
rect 10517 29257 10551 29291
rect 11529 29257 11563 29291
rect 22937 29257 22971 29291
rect 23489 29189 23523 29223
rect 8677 29121 8711 29155
rect 8944 29121 8978 29155
rect 11529 29121 11563 29155
rect 11621 29121 11655 29155
rect 22845 29121 22879 29155
rect 23029 29121 23063 29155
rect 31125 29121 31159 29155
rect 11805 29053 11839 29087
rect 12265 29053 12299 29087
rect 10057 28985 10091 29019
rect 31309 28985 31343 29019
rect 6193 28713 6227 28747
rect 6929 28713 6963 28747
rect 18337 28645 18371 28679
rect 6745 28509 6779 28543
rect 18429 28509 18463 28543
rect 18153 28441 18187 28475
rect 30665 28441 30699 28475
rect 17601 28373 17635 28407
rect 18429 28373 18463 28407
rect 26525 28373 26559 28407
rect 30757 28373 30791 28407
rect 28549 28169 28583 28203
rect 32229 28169 32263 28203
rect 29009 28101 29043 28135
rect 26157 28033 26191 28067
rect 26249 28033 26283 28067
rect 26433 28033 26467 28067
rect 27169 28033 27203 28067
rect 27436 28033 27470 28067
rect 32137 28033 32171 28067
rect 32413 28033 32447 28067
rect 37473 28033 37507 28067
rect 38117 28033 38151 28067
rect 26433 27829 26467 27863
rect 32413 27829 32447 27863
rect 37933 27829 37967 27863
rect 27353 27625 27387 27659
rect 4813 27557 4847 27591
rect 6009 27557 6043 27591
rect 18705 27557 18739 27591
rect 35633 27557 35667 27591
rect 37565 27557 37599 27591
rect 26985 27489 27019 27523
rect 31677 27489 31711 27523
rect 31769 27489 31803 27523
rect 31953 27489 31987 27523
rect 36185 27489 36219 27523
rect 4537 27421 4571 27455
rect 4629 27421 4663 27455
rect 5273 27421 5307 27455
rect 5457 27421 5491 27455
rect 17325 27421 17359 27455
rect 17592 27421 17626 27455
rect 26893 27421 26927 27455
rect 27169 27421 27203 27455
rect 31493 27421 31527 27455
rect 31585 27421 31619 27455
rect 32413 27421 32447 27455
rect 32597 27421 32631 27455
rect 36430 27353 36464 27387
rect 5365 27285 5399 27319
rect 16773 27285 16807 27319
rect 30849 27285 30883 27319
rect 32505 27285 32539 27319
rect 33885 27081 33919 27115
rect 35458 27013 35492 27047
rect 15025 26945 15059 26979
rect 35725 26945 35759 26979
rect 34345 26809 34379 26843
rect 15209 26741 15243 26775
rect 15853 26741 15887 26775
rect 4169 26537 4203 26571
rect 3985 26333 4019 26367
rect 4261 26333 4295 26367
rect 3801 26197 3835 26231
rect 3709 25993 3743 26027
rect 4261 25993 4295 26027
rect 27077 25993 27111 26027
rect 30849 25993 30883 26027
rect 23765 25925 23799 25959
rect 30205 25925 30239 25959
rect 30757 25925 30791 25959
rect 2329 25857 2363 25891
rect 2596 25857 2630 25891
rect 21833 25857 21867 25891
rect 22100 25857 22134 25891
rect 26433 25857 26467 25891
rect 27261 25857 27295 25891
rect 8493 25721 8527 25755
rect 13921 25721 13955 25755
rect 38117 25721 38151 25755
rect 23213 25653 23247 25687
rect 13093 25449 13127 25483
rect 22017 25449 22051 25483
rect 22385 25449 22419 25483
rect 31033 25449 31067 25483
rect 22937 25381 22971 25415
rect 15485 25313 15519 25347
rect 31585 25313 31619 25347
rect 6929 25245 6963 25279
rect 9229 25245 9263 25279
rect 9873 25245 9907 25279
rect 10149 25245 10183 25279
rect 10333 25245 10367 25279
rect 22201 25245 22235 25279
rect 22477 25245 22511 25279
rect 23121 25245 23155 25279
rect 23213 25245 23247 25279
rect 31493 25245 31527 25279
rect 7196 25177 7230 25211
rect 15218 25177 15252 25211
rect 22937 25177 22971 25211
rect 28825 25177 28859 25211
rect 29009 25177 29043 25211
rect 31401 25177 31435 25211
rect 32229 25177 32263 25211
rect 8309 25109 8343 25143
rect 9689 25109 9723 25143
rect 14105 25109 14139 25143
rect 23673 25109 23707 25143
rect 28181 25109 28215 25143
rect 7941 24905 7975 24939
rect 13001 24905 13035 24939
rect 8125 24769 8159 24803
rect 9321 24769 9355 24803
rect 9505 24769 9539 24803
rect 10333 24769 10367 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 12541 24769 12575 24803
rect 12633 24769 12667 24803
rect 12725 24769 12759 24803
rect 12909 24769 12943 24803
rect 13001 24769 13035 24803
rect 13645 24769 13679 24803
rect 9689 24701 9723 24735
rect 10885 24701 10919 24735
rect 13553 24701 13587 24735
rect 10149 24633 10183 24667
rect 11621 24565 11655 24599
rect 20913 24361 20947 24395
rect 25697 24361 25731 24395
rect 30389 24293 30423 24327
rect 29561 24225 29595 24259
rect 12633 24157 12667 24191
rect 12817 24157 12851 24191
rect 25053 24157 25087 24191
rect 25237 24157 25271 24191
rect 29745 24157 29779 24191
rect 30573 24157 30607 24191
rect 19625 24089 19659 24123
rect 29929 24089 29963 24123
rect 30757 24089 30791 24123
rect 31217 24089 31251 24123
rect 37381 24089 37415 24123
rect 38025 24089 38059 24123
rect 12449 24021 12483 24055
rect 25145 24021 25179 24055
rect 37933 24021 37967 24055
rect 37289 23817 37323 23851
rect 37749 23817 37783 23851
rect 31217 23749 31251 23783
rect 31401 23749 31435 23783
rect 17592 23681 17626 23715
rect 31585 23681 31619 23715
rect 37657 23681 37691 23715
rect 17325 23613 17359 23647
rect 37841 23613 37875 23647
rect 18705 23545 18739 23579
rect 16773 23477 16807 23511
rect 19441 23477 19475 23511
rect 30113 23477 30147 23511
rect 32229 23477 32263 23511
rect 17325 23273 17359 23307
rect 18061 23273 18095 23307
rect 21005 23205 21039 23239
rect 17785 23137 17819 23171
rect 32505 23137 32539 23171
rect 17969 23069 18003 23103
rect 18061 23069 18095 23103
rect 21281 23069 21315 23103
rect 25789 23069 25823 23103
rect 27629 23069 27663 23103
rect 32229 23069 32263 23103
rect 21005 23001 21039 23035
rect 21189 23001 21223 23035
rect 26056 23001 26090 23035
rect 27169 22933 27203 22967
rect 37565 22933 37599 22967
rect 38025 22933 38059 22967
rect 25973 22729 26007 22763
rect 33241 22729 33275 22763
rect 35633 22661 35667 22695
rect 37841 22661 37875 22695
rect 22017 22593 22051 22627
rect 22109 22593 22143 22627
rect 26157 22593 26191 22627
rect 33609 22593 33643 22627
rect 33701 22593 33735 22627
rect 37657 22593 37691 22627
rect 26433 22525 26467 22559
rect 33885 22525 33919 22559
rect 35081 22457 35115 22491
rect 35909 22457 35943 22491
rect 21833 22389 21867 22423
rect 26341 22389 26375 22423
rect 32689 22389 32723 22423
rect 36093 22389 36127 22423
rect 6009 22117 6043 22151
rect 20821 22049 20855 22083
rect 21189 22049 21223 22083
rect 31217 22049 31251 22083
rect 4629 21981 4663 22015
rect 21005 21981 21039 22015
rect 37473 21981 37507 22015
rect 38117 21981 38151 22015
rect 4896 21913 4930 21947
rect 30941 21913 30975 21947
rect 6561 21845 6595 21879
rect 30113 21845 30147 21879
rect 30573 21845 30607 21879
rect 31033 21845 31067 21879
rect 37933 21845 37967 21879
rect 3433 21641 3467 21675
rect 23397 21573 23431 21607
rect 2053 21505 2087 21539
rect 2320 21505 2354 21539
rect 23581 21505 23615 21539
rect 3985 21301 4019 21335
rect 6377 21097 6411 21131
rect 6561 20961 6595 20995
rect 6653 20961 6687 20995
rect 7297 20961 7331 20995
rect 37013 20961 37047 20995
rect 6745 20893 6779 20927
rect 10977 20893 11011 20927
rect 37289 20893 37323 20927
rect 11222 20825 11256 20859
rect 10425 20757 10459 20791
rect 12357 20757 12391 20791
rect 6561 20553 6595 20587
rect 6745 20553 6779 20587
rect 10149 20553 10183 20587
rect 37933 20553 37967 20587
rect 6929 20485 6963 20519
rect 28457 20485 28491 20519
rect 6837 20417 6871 20451
rect 10425 20417 10459 20451
rect 11529 20417 11563 20451
rect 15209 20417 15243 20451
rect 15945 20417 15979 20451
rect 37473 20417 37507 20451
rect 38117 20417 38151 20451
rect 7113 20349 7147 20383
rect 10333 20349 10367 20383
rect 10517 20349 10551 20383
rect 15393 20281 15427 20315
rect 28273 20281 28307 20315
rect 6837 20009 6871 20043
rect 18153 20009 18187 20043
rect 26709 20009 26743 20043
rect 12541 19941 12575 19975
rect 13093 19941 13127 19975
rect 17325 19941 17359 19975
rect 23029 19941 23063 19975
rect 27261 19941 27295 19975
rect 4169 19873 4203 19907
rect 7205 19873 7239 19907
rect 7297 19873 7331 19907
rect 18245 19873 18279 19907
rect 4353 19805 4387 19839
rect 7021 19805 7055 19839
rect 7113 19805 7147 19839
rect 10149 19805 10183 19839
rect 12725 19805 12759 19839
rect 15485 19805 15519 19839
rect 15945 19805 15979 19839
rect 17969 19805 18003 19839
rect 23305 19805 23339 19839
rect 30113 19805 30147 19839
rect 30389 19805 30423 19839
rect 30849 19805 30883 19839
rect 31033 19805 31067 19839
rect 31493 19805 31527 19839
rect 16212 19737 16246 19771
rect 17785 19737 17819 19771
rect 22569 19737 22603 19771
rect 23029 19737 23063 19771
rect 26893 19737 26927 19771
rect 10057 19669 10091 19703
rect 12817 19669 12851 19703
rect 12909 19669 12943 19703
rect 23213 19669 23247 19703
rect 26985 19669 27019 19703
rect 27077 19669 27111 19703
rect 30941 19669 30975 19703
rect 12265 19465 12299 19499
rect 19993 19465 20027 19499
rect 26985 19465 27019 19499
rect 30205 19465 30239 19499
rect 33425 19465 33459 19499
rect 34345 19465 34379 19499
rect 36277 19465 36311 19499
rect 19901 19397 19935 19431
rect 27137 19397 27171 19431
rect 27353 19397 27387 19431
rect 37473 19397 37507 19431
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 19625 19329 19659 19363
rect 19809 19329 19843 19363
rect 26157 19329 26191 19363
rect 26249 19329 26283 19363
rect 26433 19329 26467 19363
rect 31318 19329 31352 19363
rect 31585 19329 31619 19363
rect 34161 19329 34195 19363
rect 34437 19329 34471 19363
rect 34897 19329 34931 19363
rect 35153 19329 35187 19363
rect 37657 19329 37691 19363
rect 12541 19261 12575 19295
rect 12633 19261 12667 19295
rect 33977 19261 34011 19295
rect 37289 19261 37323 19295
rect 20177 19193 20211 19227
rect 26433 19125 26467 19159
rect 27169 19125 27203 19159
rect 29653 19125 29687 19159
rect 19809 18921 19843 18955
rect 23121 18921 23155 18955
rect 25697 18921 25731 18955
rect 34713 18921 34747 18955
rect 26341 18853 26375 18887
rect 26525 18785 26559 18819
rect 23029 18717 23063 18751
rect 23305 18717 23339 18751
rect 26249 18717 26283 18751
rect 37473 18717 37507 18751
rect 38117 18717 38151 18751
rect 19793 18649 19827 18683
rect 19993 18649 20027 18683
rect 19625 18581 19659 18615
rect 23489 18581 23523 18615
rect 26249 18581 26283 18615
rect 37933 18581 37967 18615
rect 2973 18377 3007 18411
rect 17785 18377 17819 18411
rect 3157 18241 3191 18275
rect 17693 18241 17727 18275
rect 17877 18241 17911 18275
rect 3433 18173 3467 18207
rect 3341 18037 3375 18071
rect 3249 17833 3283 17867
rect 8309 17833 8343 17867
rect 9781 17833 9815 17867
rect 22385 17833 22419 17867
rect 4169 17697 4203 17731
rect 3065 17629 3099 17663
rect 3249 17629 3283 17663
rect 3985 17629 4019 17663
rect 8217 17629 8251 17663
rect 8953 17629 8987 17663
rect 23498 17629 23532 17663
rect 23765 17629 23799 17663
rect 38117 17629 38151 17663
rect 3801 17493 3835 17527
rect 9137 17493 9171 17527
rect 24501 17493 24535 17527
rect 8493 17289 8527 17323
rect 7665 17153 7699 17187
rect 7849 17153 7883 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 13185 17153 13219 17187
rect 33885 17153 33919 17187
rect 7573 17085 7607 17119
rect 7757 17085 7791 17119
rect 13001 17085 13035 17119
rect 13369 17085 13403 17119
rect 34161 17085 34195 17119
rect 7389 16949 7423 16983
rect 12265 16949 12299 16983
rect 7021 16745 7055 16779
rect 12449 16745 12483 16779
rect 17877 16677 17911 16711
rect 31677 16609 31711 16643
rect 12265 16541 12299 16575
rect 12541 16541 12575 16575
rect 17693 16541 17727 16575
rect 17877 16541 17911 16575
rect 31401 16541 31435 16575
rect 7205 16473 7239 16507
rect 6837 16405 6871 16439
rect 7005 16405 7039 16439
rect 12081 16405 12115 16439
rect 37565 16405 37599 16439
rect 30665 16201 30699 16235
rect 33977 16201 34011 16235
rect 34437 16201 34471 16235
rect 37841 16201 37875 16235
rect 30021 16133 30055 16167
rect 4261 16065 4295 16099
rect 4445 16065 4479 16099
rect 18705 16065 18739 16099
rect 18889 16065 18923 16099
rect 18981 16065 19015 16099
rect 29837 16065 29871 16099
rect 30573 16065 30607 16099
rect 34345 16065 34379 16099
rect 37749 16065 37783 16099
rect 34621 15997 34655 16031
rect 4445 15861 4479 15895
rect 18521 15861 18555 15895
rect 33425 15861 33459 15895
rect 4169 15657 4203 15691
rect 12449 15657 12483 15691
rect 20637 15657 20671 15691
rect 27169 15657 27203 15691
rect 30665 15657 30699 15691
rect 32413 15657 32447 15691
rect 34805 15657 34839 15691
rect 37933 15657 37967 15691
rect 31677 15589 31711 15623
rect 31953 15521 31987 15555
rect 3985 15453 4019 15487
rect 4261 15453 4295 15487
rect 11069 15453 11103 15487
rect 18613 15453 18647 15487
rect 19257 15453 19291 15487
rect 19513 15453 19547 15487
rect 25789 15453 25823 15487
rect 27629 15453 27663 15487
rect 30481 15453 30515 15487
rect 34897 15453 34931 15487
rect 35357 15453 35391 15487
rect 38025 15453 38059 15487
rect 11336 15385 11370 15419
rect 26056 15385 26090 15419
rect 29745 15385 29779 15419
rect 30297 15385 30331 15419
rect 36461 15385 36495 15419
rect 37197 15385 37231 15419
rect 3801 15317 3835 15351
rect 10517 15317 10551 15351
rect 31493 15317 31527 15351
rect 37105 15317 37139 15351
rect 7297 15113 7331 15147
rect 17141 15113 17175 15147
rect 23213 15113 23247 15147
rect 28273 15113 28307 15147
rect 29653 15113 29687 15147
rect 36645 15113 36679 15147
rect 38025 15113 38059 15147
rect 22385 15045 22419 15079
rect 28733 15045 28767 15079
rect 29193 15045 29227 15079
rect 7481 14977 7515 15011
rect 17233 14977 17267 15011
rect 22569 14977 22603 15011
rect 36553 14977 36587 15011
rect 37289 14977 37323 15011
rect 7665 14909 7699 14943
rect 23765 14841 23799 14875
rect 27813 14841 27847 14875
rect 28457 14841 28491 14875
rect 29469 14841 29503 14875
rect 37473 14841 37507 14875
rect 14657 14773 14691 14807
rect 36001 14773 36035 14807
rect 14289 14569 14323 14603
rect 15117 14569 15151 14603
rect 15761 14569 15795 14603
rect 23857 14501 23891 14535
rect 23121 14433 23155 14467
rect 37565 14433 37599 14467
rect 7297 14365 7331 14399
rect 7573 14365 7607 14399
rect 7757 14365 7791 14399
rect 15025 14365 15059 14399
rect 22845 14365 22879 14399
rect 23673 14365 23707 14399
rect 29561 14365 29595 14399
rect 36829 14365 36863 14399
rect 37289 14365 37323 14399
rect 14841 14297 14875 14331
rect 7113 14229 7147 14263
rect 24409 14229 24443 14263
rect 4077 14025 4111 14059
rect 15117 14025 15151 14059
rect 25605 14025 25639 14059
rect 26341 14025 26375 14059
rect 31401 14025 31435 14059
rect 4537 13957 4571 13991
rect 14197 13957 14231 13991
rect 17049 13957 17083 13991
rect 24317 13957 24351 13991
rect 24501 13957 24535 13991
rect 25697 13957 25731 13991
rect 31493 13957 31527 13991
rect 37933 13957 37967 13991
rect 2697 13889 2731 13923
rect 2964 13889 2998 13923
rect 14013 13889 14047 13923
rect 17233 13889 17267 13923
rect 23765 13889 23799 13923
rect 37749 13889 37783 13923
rect 14657 13821 14691 13855
rect 23489 13821 23523 13855
rect 14933 13753 14967 13787
rect 22845 13481 22879 13515
rect 24409 13481 24443 13515
rect 23305 13345 23339 13379
rect 23489 13345 23523 13379
rect 22293 13209 22327 13243
rect 23213 13209 23247 13243
rect 14473 13141 14507 13175
rect 37565 13141 37599 13175
rect 8309 12937 8343 12971
rect 23673 12937 23707 12971
rect 8769 12869 8803 12903
rect 13277 12869 13311 12903
rect 34069 12869 34103 12903
rect 6929 12801 6963 12835
rect 7196 12801 7230 12835
rect 13093 12801 13127 12835
rect 25973 12801 26007 12835
rect 32137 12801 32171 12835
rect 33425 12801 33459 12835
rect 32413 12733 32447 12767
rect 25789 12665 25823 12699
rect 19809 12597 19843 12631
rect 33609 12597 33643 12631
rect 38117 12597 38151 12631
rect 19533 12393 19567 12427
rect 4445 12325 4479 12359
rect 9689 12325 9723 12359
rect 20637 12325 20671 12359
rect 21925 12325 21959 12359
rect 9505 12189 9539 12223
rect 31033 12189 31067 12223
rect 4261 12121 4295 12155
rect 19257 12121 19291 12155
rect 19441 12121 19475 12155
rect 20913 12121 20947 12155
rect 21465 12121 21499 12155
rect 31401 12121 31435 12155
rect 10241 12053 10275 12087
rect 18613 12053 18647 12087
rect 20453 12053 20487 12087
rect 27905 12053 27939 12087
rect 17693 11849 17727 11883
rect 19073 11849 19107 11883
rect 22385 11849 22419 11883
rect 30205 11849 30239 11883
rect 31125 11849 31159 11883
rect 2973 11781 3007 11815
rect 3709 11781 3743 11815
rect 27629 11781 27663 11815
rect 28089 11781 28123 11815
rect 30665 11781 30699 11815
rect 31585 11781 31619 11815
rect 2789 11713 2823 11747
rect 3525 11713 3559 11747
rect 10149 11713 10183 11747
rect 22293 11713 22327 11747
rect 12081 11645 12115 11679
rect 18153 11645 18187 11679
rect 18613 11645 18647 11679
rect 19533 11645 19567 11679
rect 12449 11577 12483 11611
rect 17785 11577 17819 11611
rect 18889 11577 18923 11611
rect 27261 11577 27295 11611
rect 28365 11577 28399 11611
rect 30389 11577 30423 11611
rect 31217 11577 31251 11611
rect 10333 11509 10367 11543
rect 12541 11509 12575 11543
rect 13093 11509 13127 11543
rect 27169 11509 27203 11543
rect 28549 11509 28583 11543
rect 2053 11305 2087 11339
rect 12725 11305 12759 11339
rect 27077 11305 27111 11339
rect 33241 11305 33275 11339
rect 37933 11305 37967 11339
rect 18337 11237 18371 11271
rect 28273 11237 28307 11271
rect 2881 11169 2915 11203
rect 27997 11169 28031 11203
rect 28457 11169 28491 11203
rect 2697 11101 2731 11135
rect 12817 11101 12851 11135
rect 37381 11101 37415 11135
rect 38117 11101 38151 11135
rect 13001 11033 13035 11067
rect 22109 11033 22143 11067
rect 33149 11033 33183 11067
rect 27813 10761 27847 10795
rect 5089 10693 5123 10727
rect 4905 10625 4939 10659
rect 12173 10625 12207 10659
rect 36001 10625 36035 10659
rect 36553 10625 36587 10659
rect 37289 10625 37323 10659
rect 37473 10489 37507 10523
rect 12357 10421 12391 10455
rect 17509 10421 17543 10455
rect 36737 10421 36771 10455
rect 2881 10217 2915 10251
rect 17693 10217 17727 10251
rect 6193 10149 6227 10183
rect 14841 10149 14875 10183
rect 17049 10149 17083 10183
rect 17141 10081 17175 10115
rect 15485 10013 15519 10047
rect 28457 10013 28491 10047
rect 2789 9945 2823 9979
rect 6009 9945 6043 9979
rect 14473 9945 14507 9979
rect 16681 9945 16715 9979
rect 17785 9945 17819 9979
rect 17969 9945 18003 9979
rect 14933 9877 14967 9911
rect 16221 9877 16255 9911
rect 18521 9877 18555 9911
rect 28641 9877 28675 9911
rect 17325 9673 17359 9707
rect 13461 9537 13495 9571
rect 14289 9537 14323 9571
rect 14473 9537 14507 9571
rect 24317 9537 24351 9571
rect 24777 9537 24811 9571
rect 29009 9537 29043 9571
rect 30021 9537 30055 9571
rect 37749 9537 37783 9571
rect 9873 9469 9907 9503
rect 24409 9469 24443 9503
rect 25329 9469 25363 9503
rect 38025 9469 38059 9503
rect 29193 9401 29227 9435
rect 13645 9333 13679 9367
rect 14197 9333 14231 9367
rect 30205 9333 30239 9367
rect 3801 9129 3835 9163
rect 4997 9129 5031 9163
rect 25789 9129 25823 9163
rect 34805 9129 34839 9163
rect 2881 9061 2915 9095
rect 5733 9061 5767 9095
rect 9597 9061 9631 9095
rect 10517 9061 10551 9095
rect 21005 9061 21039 9095
rect 35357 8993 35391 9027
rect 10333 8925 10367 8959
rect 20177 8925 20211 8959
rect 20637 8925 20671 8959
rect 24501 8925 24535 8959
rect 24961 8925 24995 8959
rect 25881 8925 25915 8959
rect 35909 8925 35943 8959
rect 36553 8925 36587 8959
rect 37473 8925 37507 8959
rect 38117 8925 38151 8959
rect 2513 8857 2547 8891
rect 5457 8857 5491 8891
rect 9229 8857 9263 8891
rect 10149 8857 10183 8891
rect 21649 8857 21683 8891
rect 26065 8857 26099 8891
rect 35081 8857 35115 8891
rect 2973 8789 3007 8823
rect 5917 8789 5951 8823
rect 9689 8789 9723 8823
rect 21097 8789 21131 8823
rect 24685 8789 24719 8823
rect 26525 8789 26559 8823
rect 35265 8789 35299 8823
rect 36093 8789 36127 8823
rect 37933 8789 37967 8823
rect 2697 8585 2731 8619
rect 4169 8585 4203 8619
rect 23949 8585 23983 8619
rect 38117 8585 38151 8619
rect 4077 8517 4111 8551
rect 6377 8517 6411 8551
rect 7297 8517 7331 8551
rect 20729 8517 20763 8551
rect 20913 8517 20947 8551
rect 32321 8517 32355 8551
rect 33241 8517 33275 8551
rect 33425 8517 33459 8551
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 9781 8449 9815 8483
rect 12541 8449 12575 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 32689 8449 32723 8483
rect 33609 8449 33643 8483
rect 11529 8381 11563 8415
rect 24409 8381 24443 8415
rect 32229 8381 32263 8415
rect 35725 8381 35759 8415
rect 9965 8313 9999 8347
rect 11897 8313 11931 8347
rect 20085 8313 20119 8347
rect 23489 8313 23523 8347
rect 24041 8313 24075 8347
rect 24961 8313 24995 8347
rect 25513 8313 25547 8347
rect 36277 8313 36311 8347
rect 37473 8313 37507 8347
rect 11989 8245 12023 8279
rect 37197 8041 37231 8075
rect 11805 7973 11839 8007
rect 30205 7973 30239 8007
rect 32045 7905 32079 7939
rect 11621 7837 11655 7871
rect 24869 7837 24903 7871
rect 32413 7837 32447 7871
rect 38117 7837 38151 7871
rect 11437 7769 11471 7803
rect 30021 7769 30055 7803
rect 31953 7769 31987 7803
rect 35081 7769 35115 7803
rect 37105 7769 37139 7803
rect 3249 7701 3283 7735
rect 20361 7701 20395 7735
rect 25053 7701 25087 7735
rect 35541 7701 35575 7735
rect 36553 7701 36587 7735
rect 7021 7497 7055 7531
rect 28641 7497 28675 7531
rect 7481 7429 7515 7463
rect 15209 7429 15243 7463
rect 28089 7429 28123 7463
rect 37841 7429 37875 7463
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 11529 7361 11563 7395
rect 15393 7361 15427 7395
rect 15577 7361 15611 7395
rect 26433 7361 26467 7395
rect 26985 7361 27019 7395
rect 6561 7293 6595 7327
rect 14289 7293 14323 7327
rect 20361 7293 20395 7327
rect 34069 7293 34103 7327
rect 6837 7225 6871 7259
rect 8401 7225 8435 7259
rect 14657 7225 14691 7259
rect 20637 7225 20671 7259
rect 27905 7225 27939 7259
rect 37657 7225 37691 7259
rect 11713 7157 11747 7191
rect 14749 7157 14783 7191
rect 16129 7157 16163 7191
rect 20821 7157 20855 7191
rect 27169 7157 27203 7191
rect 34621 7157 34655 7191
rect 35633 7157 35667 7191
rect 36185 7157 36219 7191
rect 36737 7157 36771 7191
rect 14933 6953 14967 6987
rect 16865 6885 16899 6919
rect 20913 6885 20947 6919
rect 31769 6885 31803 6919
rect 7113 6817 7147 6851
rect 16037 6817 16071 6851
rect 17049 6817 17083 6851
rect 25053 6817 25087 6851
rect 31125 6817 31159 6851
rect 32137 6817 32171 6851
rect 19533 6749 19567 6783
rect 27629 6749 27663 6783
rect 28273 6749 28307 6783
rect 35265 6749 35299 6783
rect 37197 6749 37231 6783
rect 37841 6749 37875 6783
rect 16589 6681 16623 6715
rect 19993 6681 20027 6715
rect 20177 6681 20211 6715
rect 20361 6681 20395 6715
rect 24869 6681 24903 6715
rect 33241 6681 33275 6715
rect 34805 6681 34839 6715
rect 36737 6681 36771 6715
rect 5273 6613 5307 6647
rect 19349 6613 19383 6647
rect 27813 6613 27847 6647
rect 29929 6613 29963 6647
rect 30573 6613 30607 6647
rect 31677 6613 31711 6647
rect 32597 6613 32631 6647
rect 33793 6613 33827 6647
rect 36093 6613 36127 6647
rect 37381 6613 37415 6647
rect 38025 6613 38059 6647
rect 4353 6409 4387 6443
rect 15577 6409 15611 6443
rect 35449 6409 35483 6443
rect 36737 6409 36771 6443
rect 16681 6341 16715 6375
rect 34805 6341 34839 6375
rect 37841 6341 37875 6375
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 35265 6273 35299 6307
rect 36093 6273 36127 6307
rect 36553 6273 36587 6307
rect 3341 6205 3375 6239
rect 3801 6205 3835 6239
rect 3709 6137 3743 6171
rect 31493 6137 31527 6171
rect 33701 6137 33735 6171
rect 35909 6137 35943 6171
rect 1501 6069 1535 6103
rect 2513 6069 2547 6103
rect 4813 6069 4847 6103
rect 5457 6069 5491 6103
rect 15117 6069 15151 6103
rect 17601 6069 17635 6103
rect 29653 6069 29687 6103
rect 30481 6069 30515 6103
rect 30941 6069 30975 6103
rect 32137 6069 32171 6103
rect 32965 6069 32999 6103
rect 34161 6069 34195 6103
rect 37749 6069 37783 6103
rect 3801 5865 3835 5899
rect 16129 5865 16163 5899
rect 18521 5865 18555 5899
rect 30665 5865 30699 5899
rect 31217 5865 31251 5899
rect 33333 5865 33367 5899
rect 33977 5865 34011 5899
rect 34897 5865 34931 5899
rect 36461 5865 36495 5899
rect 12541 5729 12575 5763
rect 29929 5729 29963 5763
rect 37841 5729 37875 5763
rect 12633 5661 12667 5695
rect 25697 5661 25731 5695
rect 26341 5661 26375 5695
rect 30113 5661 30147 5695
rect 33517 5661 33551 5695
rect 34713 5661 34747 5695
rect 35449 5661 35483 5695
rect 36645 5661 36679 5695
rect 37105 5661 37139 5695
rect 2513 5593 2547 5627
rect 3985 5593 4019 5627
rect 4169 5593 4203 5627
rect 4721 5593 4755 5627
rect 38025 5593 38059 5627
rect 1409 5525 1443 5559
rect 1961 5525 1995 5559
rect 3157 5525 3191 5559
rect 5181 5525 5215 5559
rect 5733 5525 5767 5559
rect 6377 5525 6411 5559
rect 6929 5525 6963 5559
rect 8033 5525 8067 5559
rect 9413 5525 9447 5559
rect 11069 5525 11103 5559
rect 12725 5525 12759 5559
rect 13093 5525 13127 5559
rect 14197 5525 14231 5559
rect 14657 5525 14691 5559
rect 15669 5525 15703 5559
rect 20361 5525 20395 5559
rect 21189 5525 21223 5559
rect 22109 5525 22143 5559
rect 24501 5525 24535 5559
rect 25237 5525 25271 5559
rect 25881 5525 25915 5559
rect 26893 5525 26927 5559
rect 29009 5525 29043 5559
rect 31953 5525 31987 5559
rect 32873 5525 32907 5559
rect 35633 5525 35667 5559
rect 37289 5525 37323 5559
rect 26341 5321 26375 5355
rect 29285 5321 29319 5355
rect 32137 5321 32171 5355
rect 33057 5321 33091 5355
rect 33885 5321 33919 5355
rect 34897 5321 34931 5355
rect 35541 5321 35575 5355
rect 37381 5321 37415 5355
rect 35633 5253 35667 5287
rect 29837 5185 29871 5219
rect 30573 5185 30607 5219
rect 31401 5185 31435 5219
rect 32321 5185 32355 5219
rect 33241 5185 33275 5219
rect 34069 5185 34103 5219
rect 34805 5185 34839 5219
rect 36461 5185 36495 5219
rect 38117 5185 38151 5219
rect 12265 5117 12299 5151
rect 4537 5049 4571 5083
rect 30021 5049 30055 5083
rect 37933 5049 37967 5083
rect 1501 4981 1535 5015
rect 1961 4981 1995 5015
rect 2605 4981 2639 5015
rect 3065 4981 3099 5015
rect 3709 4981 3743 5015
rect 4997 4981 5031 5015
rect 5825 4981 5859 5015
rect 6469 4981 6503 5015
rect 7205 4981 7239 5015
rect 7941 4981 7975 5015
rect 8493 4981 8527 5015
rect 9045 4981 9079 5015
rect 9597 4981 9631 5015
rect 10149 4981 10183 5015
rect 10701 4981 10735 5015
rect 11713 4981 11747 5015
rect 12817 4981 12851 5015
rect 13369 4981 13403 5015
rect 14013 4981 14047 5015
rect 14841 4981 14875 5015
rect 15761 4981 15795 5015
rect 16681 4981 16715 5015
rect 17233 4981 17267 5015
rect 18337 4981 18371 5015
rect 18981 4981 19015 5015
rect 19441 4981 19475 5015
rect 20361 4981 20395 5015
rect 21097 4981 21131 5015
rect 21833 4981 21867 5015
rect 22385 4981 22419 5015
rect 22937 4981 22971 5015
rect 23765 4981 23799 5015
rect 24317 4981 24351 5015
rect 25053 4981 25087 5015
rect 25789 4981 25823 5015
rect 27537 4981 27571 5015
rect 27997 4981 28031 5015
rect 28641 4981 28675 5015
rect 31585 4981 31619 5015
rect 36645 4981 36679 5015
rect 2237 4777 2271 4811
rect 9597 4777 9631 4811
rect 14105 4777 14139 4811
rect 25145 4777 25179 4811
rect 30573 4777 30607 4811
rect 33425 4777 33459 4811
rect 1593 4709 1627 4743
rect 5549 4709 5583 4743
rect 12265 4709 12299 4743
rect 21097 4709 21131 4743
rect 27997 4709 28031 4743
rect 32321 4709 32355 4743
rect 35357 4709 35391 4743
rect 8401 4641 8435 4675
rect 25973 4641 26007 4675
rect 1409 4573 1443 4607
rect 2053 4573 2087 4607
rect 2697 4573 2731 4607
rect 5365 4573 5399 4607
rect 7113 4573 7147 4607
rect 11345 4573 11379 4607
rect 13001 4573 13035 4607
rect 14289 4573 14323 4607
rect 15761 4573 15795 4607
rect 16589 4573 16623 4607
rect 20085 4573 20119 4607
rect 20913 4573 20947 4607
rect 21557 4573 21591 4607
rect 22201 4573 22235 4607
rect 25329 4573 25363 4607
rect 26433 4573 26467 4607
rect 26617 4573 26651 4607
rect 26709 4573 26743 4607
rect 30389 4573 30423 4607
rect 31033 4573 31067 4607
rect 32137 4573 32171 4607
rect 33241 4573 33275 4607
rect 33977 4573 34011 4607
rect 36093 4573 36127 4607
rect 38117 4573 38151 4607
rect 8217 4505 8251 4539
rect 9045 4505 9079 4539
rect 9137 4505 9171 4539
rect 9321 4505 9355 4539
rect 17141 4505 17175 4539
rect 28549 4505 28583 4539
rect 35173 4505 35207 4539
rect 37197 4505 37231 4539
rect 37381 4505 37415 4539
rect 2881 4437 2915 4471
rect 3893 4437 3927 4471
rect 4353 4437 4387 4471
rect 6101 4437 6135 4471
rect 6561 4437 6595 4471
rect 7297 4437 7331 4471
rect 10149 4437 10183 4471
rect 11161 4437 11195 4471
rect 12817 4437 12851 4471
rect 13553 4437 13587 4471
rect 14933 4437 14967 4471
rect 15577 4437 15611 4471
rect 16405 4437 16439 4471
rect 17601 4437 17635 4471
rect 18153 4437 18187 4471
rect 19625 4437 19659 4471
rect 20269 4437 20303 4471
rect 21741 4437 21775 4471
rect 22385 4437 22419 4471
rect 22937 4437 22971 4471
rect 23765 4437 23799 4471
rect 24593 4437 24627 4471
rect 27445 4437 27479 4471
rect 29653 4437 29687 4471
rect 31217 4437 31251 4471
rect 34161 4437 34195 4471
rect 36277 4437 36311 4471
rect 2789 4233 2823 4267
rect 10149 4233 10183 4267
rect 12357 4233 12391 4267
rect 19257 4233 19291 4267
rect 20545 4233 20579 4267
rect 20913 4233 20947 4267
rect 24501 4233 24535 4267
rect 27629 4233 27663 4267
rect 7481 4165 7515 4199
rect 36553 4165 36587 4199
rect 1409 4097 1443 4131
rect 2881 4097 2915 4131
rect 3617 4097 3651 4131
rect 4261 4097 4295 4131
rect 4905 4097 4939 4131
rect 5549 4097 5583 4131
rect 6469 4097 6503 4131
rect 8953 4097 8987 4131
rect 11897 4097 11931 4131
rect 12541 4097 12575 4131
rect 13001 4097 13035 4131
rect 13737 4097 13771 4131
rect 14749 4097 14783 4131
rect 15485 4097 15519 4131
rect 17417 4097 17451 4131
rect 19349 4097 19383 4131
rect 22385 4097 22419 4131
rect 23213 4097 23247 4131
rect 24041 4097 24075 4131
rect 25237 4097 25271 4131
rect 27169 4097 27203 4131
rect 27813 4097 27847 4131
rect 28641 4097 28675 4131
rect 30481 4097 30515 4131
rect 31033 4097 31067 4131
rect 32137 4097 32171 4131
rect 32873 4097 32907 4131
rect 33977 4097 34011 4131
rect 35265 4097 35299 4131
rect 37289 4097 37323 4131
rect 38117 4097 38151 4131
rect 3065 4029 3099 4063
rect 7665 4029 7699 4063
rect 8677 4029 8711 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 19073 4029 19107 4063
rect 20269 4029 20303 4063
rect 20453 4029 20487 4063
rect 25697 4029 25731 4063
rect 26157 4029 26191 4063
rect 29837 4029 29871 4063
rect 2421 3961 2455 3995
rect 4445 3961 4479 3995
rect 5733 3961 5767 3995
rect 10609 3961 10643 3995
rect 11713 3961 11747 3995
rect 13921 3961 13955 3995
rect 17969 3961 18003 3995
rect 19717 3961 19751 3995
rect 25053 3961 25087 3995
rect 26065 3961 26099 3995
rect 26985 3961 27019 3995
rect 29469 3961 29503 3995
rect 30297 3961 30331 3995
rect 31217 3961 31251 3995
rect 34713 3961 34747 3995
rect 37473 3961 37507 3995
rect 1593 3893 1627 3927
rect 3801 3893 3835 3927
rect 5089 3893 5123 3927
rect 6653 3893 6687 3927
rect 8125 3893 8159 3927
rect 13185 3893 13219 3927
rect 14565 3893 14599 3927
rect 15301 3893 15335 3927
rect 16129 3893 16163 3927
rect 17233 3893 17267 3927
rect 18429 3893 18463 3927
rect 22201 3893 22235 3927
rect 23029 3893 23063 3927
rect 23857 3893 23891 3927
rect 28825 3893 28859 3927
rect 29377 3893 29411 3927
rect 32321 3893 32355 3927
rect 33057 3893 33091 3927
rect 34161 3893 34195 3927
rect 35449 3893 35483 3927
rect 36461 3893 36495 3927
rect 4997 3689 5031 3723
rect 6193 3689 6227 3723
rect 11529 3689 11563 3723
rect 13185 3689 13219 3723
rect 14105 3689 14139 3723
rect 16957 3689 16991 3723
rect 19349 3689 19383 3723
rect 19993 3689 20027 3723
rect 20729 3689 20763 3723
rect 22569 3689 22603 3723
rect 23765 3689 23799 3723
rect 3985 3621 4019 3655
rect 7757 3621 7791 3655
rect 16497 3621 16531 3655
rect 31585 3621 31619 3655
rect 36185 3621 36219 3655
rect 5457 3553 5491 3587
rect 5549 3553 5583 3587
rect 6653 3553 6687 3587
rect 6745 3553 6779 3587
rect 9781 3553 9815 3587
rect 12541 3553 12575 3587
rect 14657 3553 14691 3587
rect 15853 3553 15887 3587
rect 16037 3553 16071 3587
rect 17509 3553 17543 3587
rect 21925 3553 21959 3587
rect 22109 3553 22143 3587
rect 23121 3553 23155 3587
rect 30297 3553 30331 3587
rect 37841 3553 37875 3587
rect 38117 3553 38151 3587
rect 1777 3485 1811 3519
rect 2053 3485 2087 3519
rect 3249 3485 3283 3519
rect 3801 3485 3835 3519
rect 8217 3485 8251 3519
rect 9505 3485 9539 3519
rect 11253 3485 11287 3519
rect 14565 3485 14599 3519
rect 16129 3485 16163 3519
rect 17325 3485 17359 3519
rect 18429 3485 18463 3519
rect 19533 3485 19567 3519
rect 20545 3485 20579 3519
rect 21189 3485 21223 3519
rect 22201 3485 22235 3519
rect 23397 3485 23431 3519
rect 25237 3485 25271 3519
rect 25421 3485 25455 3519
rect 26525 3485 26559 3519
rect 26985 3485 27019 3519
rect 27813 3485 27847 3519
rect 28825 3485 28859 3519
rect 30021 3485 30055 3519
rect 31401 3485 31435 3519
rect 32045 3485 32079 3519
rect 32781 3485 32815 3519
rect 33885 3485 33919 3519
rect 35265 3485 35299 3519
rect 36369 3485 36403 3519
rect 4537 3417 4571 3451
rect 5365 3417 5399 3451
rect 6561 3417 6595 3451
rect 7573 3417 7607 3451
rect 8953 3417 8987 3451
rect 10977 3417 11011 3451
rect 14473 3417 14507 3451
rect 17417 3417 17451 3451
rect 24593 3417 24627 3451
rect 24777 3417 24811 3451
rect 28641 3417 28675 3451
rect 29009 3417 29043 3451
rect 35081 3417 35115 3451
rect 3065 3349 3099 3383
rect 8401 3349 8435 3383
rect 11069 3349 11103 3383
rect 12725 3349 12759 3383
rect 12817 3349 12851 3383
rect 18245 3349 18279 3383
rect 21373 3349 21407 3383
rect 23305 3349 23339 3383
rect 25605 3349 25639 3383
rect 26341 3349 26375 3383
rect 27169 3349 27203 3383
rect 27997 3349 28031 3383
rect 32229 3349 32263 3383
rect 32965 3349 32999 3383
rect 34069 3349 34103 3383
rect 2973 3145 3007 3179
rect 3433 3145 3467 3179
rect 5825 3145 5859 3179
rect 9597 3145 9631 3179
rect 13737 3145 13771 3179
rect 14565 3145 14599 3179
rect 15393 3145 15427 3179
rect 15945 3145 15979 3179
rect 16865 3145 16899 3179
rect 18613 3145 18647 3179
rect 20085 3145 20119 3179
rect 24869 3145 24903 3179
rect 36645 3145 36679 3179
rect 3065 3077 3099 3111
rect 4169 3077 4203 3111
rect 4905 3077 4939 3111
rect 17969 3077 18003 3111
rect 28365 3077 28399 3111
rect 28825 3077 28859 3111
rect 29561 3077 29595 3111
rect 34897 3077 34931 3111
rect 35725 3077 35759 3111
rect 1409 3009 1443 3043
rect 3985 3009 4019 3043
rect 4721 3009 4755 3043
rect 5641 3009 5675 3043
rect 6801 3009 6835 3043
rect 8125 3009 8159 3043
rect 9413 3009 9447 3043
rect 11529 3009 11563 3043
rect 12265 3009 12299 3043
rect 13001 3009 13035 3043
rect 13921 3009 13955 3043
rect 14381 3009 14415 3043
rect 15209 3009 15243 3043
rect 16129 3009 16163 3043
rect 16681 3009 16715 3043
rect 17785 3009 17819 3043
rect 18429 3009 18463 3043
rect 19441 3009 19475 3043
rect 19901 3009 19935 3043
rect 21005 3009 21039 3043
rect 22109 3009 22143 3043
rect 22937 3009 22971 3043
rect 24041 3009 24075 3043
rect 24777 3009 24811 3043
rect 25421 3009 25455 3043
rect 26157 3009 26191 3043
rect 27721 3009 27755 3043
rect 29009 3009 29043 3043
rect 29745 3009 29779 3043
rect 30573 3009 30607 3043
rect 30849 3009 30883 3043
rect 32505 3009 32539 3043
rect 33793 3009 33827 3043
rect 35081 3009 35115 3043
rect 36461 3009 36495 3043
rect 37289 3009 37323 3043
rect 1685 2941 1719 2975
rect 2789 2941 2823 2975
rect 7021 2941 7055 2975
rect 8401 2941 8435 2975
rect 10057 2941 10091 2975
rect 10333 2941 10367 2975
rect 22661 2941 22695 2975
rect 24225 2941 24259 2975
rect 32781 2941 32815 2975
rect 37565 2941 37599 2975
rect 13185 2873 13219 2907
rect 25605 2873 25639 2907
rect 26341 2873 26375 2907
rect 27537 2873 27571 2907
rect 35541 2873 35575 2907
rect 7573 2805 7607 2839
rect 11713 2805 11747 2839
rect 12449 2805 12483 2839
rect 19257 2805 19291 2839
rect 20821 2805 20855 2839
rect 21925 2805 21959 2839
rect 26985 2805 27019 2839
rect 33977 2805 34011 2839
rect 6607 2601 6641 2635
rect 12817 2601 12851 2635
rect 15945 2601 15979 2635
rect 21925 2601 21959 2635
rect 23857 2601 23891 2635
rect 34897 2601 34931 2635
rect 18521 2533 18555 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 4537 2465 4571 2499
rect 4813 2465 4847 2499
rect 9229 2465 9263 2499
rect 24685 2465 24719 2499
rect 30021 2465 30055 2499
rect 32229 2465 32263 2499
rect 32505 2465 32539 2499
rect 35909 2465 35943 2499
rect 37565 2465 37599 2499
rect 2789 2397 2823 2431
rect 3893 2397 3927 2431
rect 6377 2397 6411 2431
rect 7757 2397 7791 2431
rect 9505 2397 9539 2431
rect 10609 2397 10643 2431
rect 10793 2397 10827 2431
rect 12633 2397 12667 2431
rect 14105 2397 14139 2431
rect 14933 2397 14967 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 20361 2397 20395 2431
rect 22385 2397 22419 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 27537 2397 27571 2431
rect 28089 2397 28123 2431
rect 29009 2397 29043 2431
rect 29745 2397 29779 2431
rect 34069 2397 34103 2431
rect 34713 2397 34747 2431
rect 36185 2397 36219 2431
rect 37289 2397 37323 2431
rect 11989 2329 12023 2363
rect 12173 2329 12207 2363
rect 18337 2329 18371 2363
rect 19717 2329 19751 2363
rect 19901 2329 19935 2363
rect 21281 2329 21315 2363
rect 26157 2329 26191 2363
rect 26341 2329 26375 2363
rect 27353 2329 27387 2363
rect 28273 2329 28307 2363
rect 31217 2329 31251 2363
rect 33885 2329 33919 2363
rect 2881 2261 2915 2295
rect 3985 2261 4019 2295
rect 7849 2261 7883 2295
rect 13461 2261 13495 2295
rect 14289 2261 14323 2295
rect 15117 2261 15151 2295
rect 16865 2261 16899 2295
rect 17601 2261 17635 2295
rect 20545 2261 20579 2295
rect 22615 2261 22649 2295
rect 28825 2261 28859 2295
rect 31125 2261 31159 2295
<< metal1 >>
rect 9674 37612 9680 37664
rect 9732 37652 9738 37664
rect 16022 37652 16028 37664
rect 9732 37624 16028 37652
rect 9732 37612 9738 37624
rect 16022 37612 16028 37624
rect 16080 37612 16086 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 4249 37451 4307 37457
rect 4249 37417 4261 37451
rect 4295 37448 4307 37451
rect 4890 37448 4896 37460
rect 4295 37420 4896 37448
rect 4295 37417 4307 37420
rect 4249 37411 4307 37417
rect 4890 37408 4896 37420
rect 4948 37408 4954 37460
rect 9674 37448 9680 37460
rect 9635 37420 9680 37448
rect 9674 37408 9680 37420
rect 9732 37408 9738 37460
rect 14550 37408 14556 37460
rect 14608 37448 14614 37460
rect 15933 37451 15991 37457
rect 15933 37448 15945 37451
rect 14608 37420 15945 37448
rect 14608 37408 14614 37420
rect 15933 37417 15945 37420
rect 15979 37417 15991 37451
rect 15933 37411 15991 37417
rect 16022 37408 16028 37460
rect 16080 37448 16086 37460
rect 29086 37448 29092 37460
rect 16080 37420 29092 37448
rect 16080 37408 16086 37420
rect 29086 37408 29092 37420
rect 29144 37408 29150 37460
rect 7101 37383 7159 37389
rect 7101 37349 7113 37383
rect 7147 37380 7159 37383
rect 7650 37380 7656 37392
rect 7147 37352 7656 37380
rect 7147 37349 7159 37352
rect 7101 37343 7159 37349
rect 7650 37340 7656 37352
rect 7708 37340 7714 37392
rect 13173 37383 13231 37389
rect 13173 37349 13185 37383
rect 13219 37380 13231 37383
rect 28442 37380 28448 37392
rect 13219 37352 28448 37380
rect 13219 37349 13231 37352
rect 13173 37343 13231 37349
rect 28442 37340 28448 37352
rect 28500 37340 28506 37392
rect 2961 37315 3019 37321
rect 2961 37281 2973 37315
rect 3007 37312 3019 37315
rect 3510 37312 3516 37324
rect 3007 37284 3516 37312
rect 3007 37281 3019 37284
rect 2961 37275 3019 37281
rect 3510 37272 3516 37284
rect 3568 37272 3574 37324
rect 4893 37315 4951 37321
rect 4893 37281 4905 37315
rect 4939 37312 4951 37315
rect 5074 37312 5080 37324
rect 4939 37284 5080 37312
rect 4939 37281 4951 37284
rect 4893 37275 4951 37281
rect 5074 37272 5080 37284
rect 5132 37272 5138 37324
rect 14737 37315 14795 37321
rect 14737 37281 14749 37315
rect 14783 37312 14795 37315
rect 14918 37312 14924 37324
rect 14783 37284 14924 37312
rect 14783 37281 14795 37284
rect 14737 37275 14795 37281
rect 14918 37272 14924 37284
rect 14976 37272 14982 37324
rect 15473 37315 15531 37321
rect 15473 37281 15485 37315
rect 15519 37312 15531 37315
rect 16022 37312 16028 37324
rect 15519 37284 16028 37312
rect 15519 37281 15531 37284
rect 15473 37275 15531 37281
rect 16022 37272 16028 37284
rect 16080 37272 16086 37324
rect 17037 37315 17095 37321
rect 17037 37281 17049 37315
rect 17083 37312 17095 37315
rect 17402 37312 17408 37324
rect 17083 37284 17408 37312
rect 17083 37281 17095 37284
rect 17037 37275 17095 37281
rect 17402 37272 17408 37284
rect 17460 37272 17466 37324
rect 18417 37315 18475 37321
rect 18417 37281 18429 37315
rect 18463 37312 18475 37315
rect 18874 37312 18880 37324
rect 18463 37284 18880 37312
rect 18463 37281 18475 37284
rect 18417 37275 18475 37281
rect 18874 37272 18880 37284
rect 18932 37272 18938 37324
rect 22189 37315 22247 37321
rect 22189 37281 22201 37315
rect 22235 37312 22247 37315
rect 22646 37312 22652 37324
rect 22235 37284 22652 37312
rect 22235 37281 22247 37284
rect 22189 37275 22247 37281
rect 22646 37272 22652 37284
rect 22704 37272 22710 37324
rect 23661 37315 23719 37321
rect 23661 37312 23673 37315
rect 22756 37284 23673 37312
rect 1118 37204 1124 37256
rect 1176 37244 1182 37256
rect 1762 37244 1768 37256
rect 1176 37216 1768 37244
rect 1176 37204 1182 37216
rect 1762 37204 1768 37216
rect 1820 37244 1826 37256
rect 1857 37247 1915 37253
rect 1857 37244 1869 37247
rect 1820 37216 1869 37244
rect 1820 37204 1826 37216
rect 1857 37213 1869 37216
rect 1903 37213 1915 37247
rect 1857 37207 1915 37213
rect 2130 37204 2136 37256
rect 2188 37244 2194 37256
rect 2590 37244 2596 37256
rect 2188 37216 2596 37244
rect 2188 37204 2194 37216
rect 2590 37204 2596 37216
rect 2648 37244 2654 37256
rect 2777 37247 2835 37253
rect 2777 37244 2789 37247
rect 2648 37216 2789 37244
rect 2648 37204 2654 37216
rect 2777 37213 2789 37216
rect 2823 37213 2835 37247
rect 2777 37207 2835 37213
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4062 37244 4068 37256
rect 3292 37216 4068 37244
rect 3292 37204 3298 37216
rect 4062 37204 4068 37216
rect 4120 37244 4126 37256
rect 4341 37247 4399 37253
rect 4341 37244 4353 37247
rect 4120 37216 4353 37244
rect 4120 37204 4126 37216
rect 4341 37213 4353 37216
rect 4387 37213 4399 37247
rect 4341 37207 4399 37213
rect 5718 37204 5724 37256
rect 5776 37244 5782 37256
rect 5813 37247 5871 37253
rect 5813 37244 5825 37247
rect 5776 37216 5825 37244
rect 5776 37204 5782 37216
rect 5813 37213 5825 37216
rect 5859 37213 5871 37247
rect 5813 37207 5871 37213
rect 6362 37204 6368 37256
rect 6420 37244 6426 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6420 37216 6837 37244
rect 6420 37204 6426 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 6825 37207 6883 37213
rect 7466 37204 7472 37256
rect 7524 37244 7530 37256
rect 7653 37247 7711 37253
rect 7653 37244 7665 37247
rect 7524 37216 7665 37244
rect 7524 37204 7530 37216
rect 7653 37213 7665 37216
rect 7699 37213 7711 37247
rect 7653 37207 7711 37213
rect 8478 37204 8484 37256
rect 8536 37244 8542 37256
rect 9398 37244 9404 37256
rect 8536 37216 9404 37244
rect 8536 37204 8542 37216
rect 9398 37204 9404 37216
rect 9456 37204 9462 37256
rect 10134 37204 10140 37256
rect 10192 37244 10198 37256
rect 10229 37247 10287 37253
rect 10229 37244 10241 37247
rect 10192 37216 10241 37244
rect 10192 37204 10198 37216
rect 10229 37213 10241 37216
rect 10275 37213 10287 37247
rect 10229 37207 10287 37213
rect 10594 37204 10600 37256
rect 10652 37244 10658 37256
rect 11977 37247 12035 37253
rect 11977 37244 11989 37247
rect 10652 37216 11989 37244
rect 10652 37204 10658 37216
rect 11977 37213 11989 37216
rect 12023 37244 12035 37247
rect 12158 37244 12164 37256
rect 12023 37216 12164 37244
rect 12023 37213 12035 37216
rect 11977 37207 12035 37213
rect 12158 37204 12164 37216
rect 12216 37204 12222 37256
rect 13814 37204 13820 37256
rect 13872 37244 13878 37256
rect 14550 37244 14556 37256
rect 13872 37216 14556 37244
rect 13872 37204 13878 37216
rect 14550 37204 14556 37216
rect 14608 37204 14614 37256
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15286 37244 15292 37256
rect 14884 37216 15292 37244
rect 14884 37204 14890 37216
rect 15286 37204 15292 37216
rect 15344 37204 15350 37256
rect 17954 37204 17960 37256
rect 18012 37244 18018 37256
rect 18141 37247 18199 37253
rect 18141 37244 18153 37247
rect 18012 37216 18153 37244
rect 18012 37204 18018 37216
rect 18141 37213 18153 37216
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 19058 37204 19064 37256
rect 19116 37244 19122 37256
rect 19242 37244 19248 37256
rect 19116 37216 19248 37244
rect 19116 37204 19122 37216
rect 19242 37204 19248 37216
rect 19300 37204 19306 37256
rect 20070 37204 20076 37256
rect 20128 37244 20134 37256
rect 20165 37247 20223 37253
rect 20165 37244 20177 37247
rect 20128 37216 20177 37244
rect 20128 37204 20134 37216
rect 20165 37213 20177 37216
rect 20211 37213 20223 37247
rect 20898 37244 20904 37256
rect 20859 37216 20904 37244
rect 20165 37207 20223 37213
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 21082 37204 21088 37256
rect 21140 37244 21146 37256
rect 22373 37247 22431 37253
rect 22373 37244 22385 37247
rect 21140 37216 22385 37244
rect 21140 37204 21146 37216
rect 22373 37213 22385 37216
rect 22419 37244 22431 37247
rect 22756 37244 22784 37284
rect 23661 37281 23673 37284
rect 23707 37281 23719 37315
rect 30650 37312 30656 37324
rect 30611 37284 30656 37312
rect 23661 37275 23719 37281
rect 30650 37272 30656 37284
rect 30708 37272 30714 37324
rect 32306 37272 32312 37324
rect 32364 37312 32370 37324
rect 32493 37315 32551 37321
rect 32493 37312 32505 37315
rect 32364 37284 32505 37312
rect 32364 37272 32370 37284
rect 32493 37281 32505 37284
rect 32539 37281 32551 37315
rect 33965 37315 34023 37321
rect 33965 37312 33977 37315
rect 32493 37275 32551 37281
rect 32692 37284 33977 37312
rect 22419 37216 22784 37244
rect 22925 37247 22983 37253
rect 22419 37213 22431 37216
rect 22373 37207 22431 37213
rect 22925 37213 22937 37247
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 4154 37136 4160 37188
rect 4212 37176 4218 37188
rect 5077 37179 5135 37185
rect 5077 37176 5089 37179
rect 4212 37148 5089 37176
rect 4212 37136 4218 37148
rect 5077 37145 5089 37148
rect 5123 37176 5135 37179
rect 5258 37176 5264 37188
rect 5123 37148 5264 37176
rect 5123 37145 5135 37148
rect 5077 37139 5135 37145
rect 5258 37136 5264 37148
rect 5316 37136 5322 37188
rect 11606 37136 11612 37188
rect 11664 37176 11670 37188
rect 12897 37179 12955 37185
rect 12897 37176 12909 37179
rect 11664 37148 12909 37176
rect 11664 37136 11670 37148
rect 12897 37145 12909 37148
rect 12943 37176 12955 37179
rect 13722 37176 13728 37188
rect 12943 37148 13728 37176
rect 12943 37145 12955 37148
rect 12897 37139 12955 37145
rect 13722 37136 13728 37148
rect 13780 37136 13786 37188
rect 15838 37136 15844 37188
rect 15896 37176 15902 37188
rect 17221 37179 17279 37185
rect 17221 37176 17233 37179
rect 15896 37148 17233 37176
rect 15896 37136 15902 37148
rect 17221 37145 17233 37148
rect 17267 37176 17279 37179
rect 17494 37176 17500 37188
rect 17267 37148 17500 37176
rect 17267 37145 17279 37148
rect 17221 37139 17279 37145
rect 17494 37136 17500 37148
rect 17552 37136 17558 37188
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 22940 37176 22968 37207
rect 24302 37204 24308 37256
rect 24360 37244 24366 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 24360 37216 24409 37244
rect 24360 37204 24366 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 25314 37204 25320 37256
rect 25372 37244 25378 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25372 37216 25421 37244
rect 25372 37204 25378 37216
rect 25409 37213 25421 37216
rect 25455 37213 25467 37247
rect 25409 37207 25467 37213
rect 25498 37204 25504 37256
rect 25556 37244 25562 37256
rect 26145 37247 26203 37253
rect 26145 37244 26157 37247
rect 25556 37216 26157 37244
rect 25556 37204 25562 37216
rect 26145 37213 26157 37216
rect 26191 37213 26203 37247
rect 26970 37244 26976 37256
rect 26931 37216 26976 37244
rect 26145 37207 26203 37213
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27893 37247 27951 37253
rect 27893 37244 27905 37247
rect 27120 37216 27905 37244
rect 27120 37204 27126 37216
rect 27893 37213 27905 37216
rect 27939 37213 27951 37247
rect 27893 37207 27951 37213
rect 28534 37204 28540 37256
rect 28592 37244 28598 37256
rect 28813 37247 28871 37253
rect 28813 37244 28825 37247
rect 28592 37216 28825 37244
rect 28592 37204 28598 37216
rect 28813 37213 28825 37216
rect 28859 37244 28871 37247
rect 28902 37244 28908 37256
rect 28859 37216 28908 37244
rect 28859 37213 28871 37216
rect 28813 37207 28871 37213
rect 28902 37204 28908 37216
rect 28960 37204 28966 37256
rect 29454 37204 29460 37256
rect 29512 37244 29518 37256
rect 29549 37247 29607 37253
rect 29549 37244 29561 37247
rect 29512 37216 29561 37244
rect 29512 37204 29518 37216
rect 29549 37213 29561 37216
rect 29595 37213 29607 37247
rect 29549 37207 29607 37213
rect 30558 37204 30564 37256
rect 30616 37244 30622 37256
rect 30837 37247 30895 37253
rect 30837 37244 30849 37247
rect 30616 37216 30849 37244
rect 30616 37204 30622 37216
rect 30837 37213 30849 37216
rect 30883 37213 30895 37247
rect 30837 37207 30895 37213
rect 31573 37247 31631 37253
rect 31573 37213 31585 37247
rect 31619 37213 31631 37247
rect 31573 37207 31631 37213
rect 22244 37148 22968 37176
rect 22244 37136 22250 37148
rect 29638 37136 29644 37188
rect 29696 37176 29702 37188
rect 31202 37176 31208 37188
rect 29696 37148 31208 37176
rect 29696 37136 29702 37148
rect 31202 37136 31208 37148
rect 31260 37176 31266 37188
rect 31588 37176 31616 37207
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32692 37253 32720 37284
rect 33965 37281 33977 37284
rect 34011 37281 34023 37315
rect 38013 37315 38071 37321
rect 38013 37312 38025 37315
rect 33965 37275 34023 37281
rect 34716 37284 34928 37312
rect 32677 37247 32735 37253
rect 32677 37244 32689 37247
rect 31812 37216 32689 37244
rect 31812 37204 31818 37216
rect 32677 37213 32689 37216
rect 32723 37213 32735 37247
rect 32677 37207 32735 37213
rect 32766 37204 32772 37256
rect 32824 37244 32830 37256
rect 33502 37244 33508 37256
rect 32824 37216 33508 37244
rect 32824 37204 32830 37216
rect 33502 37204 33508 37216
rect 33560 37204 33566 37256
rect 33778 37204 33784 37256
rect 33836 37244 33842 37256
rect 34716 37244 34744 37284
rect 33836 37216 34744 37244
rect 34900 37244 34928 37284
rect 36464 37284 38025 37312
rect 34977 37247 35035 37253
rect 34977 37244 34989 37247
rect 34900 37216 34989 37244
rect 33836 37204 33842 37216
rect 34977 37213 34989 37216
rect 35023 37244 35035 37247
rect 35434 37244 35440 37256
rect 35023 37216 35440 37244
rect 35023 37213 35035 37216
rect 34977 37207 35035 37213
rect 35434 37204 35440 37216
rect 35492 37204 35498 37256
rect 35710 37244 35716 37256
rect 35671 37216 35716 37244
rect 35710 37204 35716 37216
rect 35768 37204 35774 37256
rect 35894 37204 35900 37256
rect 35952 37244 35958 37256
rect 36464 37253 36492 37284
rect 38013 37281 38025 37284
rect 38059 37281 38071 37315
rect 38013 37275 38071 37281
rect 36449 37247 36507 37253
rect 36449 37244 36461 37247
rect 35952 37216 36461 37244
rect 35952 37204 35958 37216
rect 36449 37213 36461 37216
rect 36495 37213 36507 37247
rect 37274 37244 37280 37256
rect 37235 37216 37280 37244
rect 36449 37207 36507 37213
rect 37274 37204 37280 37216
rect 37332 37204 37338 37256
rect 38378 37176 38384 37188
rect 31260 37148 31616 37176
rect 37476 37148 38384 37176
rect 31260 37136 31266 37148
rect 1946 37108 1952 37120
rect 1907 37080 1952 37108
rect 1946 37068 1952 37080
rect 2004 37068 2010 37120
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 5629 37111 5687 37117
rect 5629 37108 5641 37111
rect 2832 37080 5641 37108
rect 2832 37068 2838 37080
rect 5629 37077 5641 37080
rect 5675 37077 5687 37111
rect 7834 37108 7840 37120
rect 7795 37080 7840 37108
rect 5629 37071 5687 37077
rect 7834 37068 7840 37080
rect 7892 37068 7898 37120
rect 10413 37111 10471 37117
rect 10413 37077 10425 37111
rect 10459 37108 10471 37111
rect 10594 37108 10600 37120
rect 10459 37080 10600 37108
rect 10459 37077 10471 37080
rect 10413 37071 10471 37077
rect 10594 37068 10600 37080
rect 10652 37068 10658 37120
rect 12066 37108 12072 37120
rect 12027 37080 12072 37108
rect 12066 37068 12072 37080
rect 12124 37068 12130 37120
rect 19429 37111 19487 37117
rect 19429 37077 19441 37111
rect 19475 37108 19487 37111
rect 20162 37108 20168 37120
rect 19475 37080 20168 37108
rect 19475 37077 19487 37080
rect 19429 37071 19487 37077
rect 20162 37068 20168 37080
rect 20220 37068 20226 37120
rect 20346 37108 20352 37120
rect 20307 37080 20352 37108
rect 20346 37068 20352 37080
rect 20404 37068 20410 37120
rect 20438 37068 20444 37120
rect 20496 37108 20502 37120
rect 21085 37111 21143 37117
rect 21085 37108 21097 37111
rect 20496 37080 21097 37108
rect 20496 37068 20502 37080
rect 21085 37077 21097 37080
rect 21131 37077 21143 37111
rect 21085 37071 21143 37077
rect 23014 37068 23020 37120
rect 23072 37108 23078 37120
rect 23109 37111 23167 37117
rect 23109 37108 23121 37111
rect 23072 37080 23121 37108
rect 23072 37068 23078 37080
rect 23109 37077 23121 37080
rect 23155 37077 23167 37111
rect 24578 37108 24584 37120
rect 24539 37080 24584 37108
rect 23109 37071 23167 37077
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 25590 37108 25596 37120
rect 25551 37080 25596 37108
rect 25590 37068 25596 37080
rect 25648 37068 25654 37120
rect 25682 37068 25688 37120
rect 25740 37108 25746 37120
rect 26329 37111 26387 37117
rect 26329 37108 26341 37111
rect 25740 37080 26341 37108
rect 25740 37068 25746 37080
rect 26329 37077 26341 37080
rect 26375 37077 26387 37111
rect 26329 37071 26387 37077
rect 26786 37068 26792 37120
rect 26844 37108 26850 37120
rect 27157 37111 27215 37117
rect 27157 37108 27169 37111
rect 26844 37080 27169 37108
rect 26844 37068 26850 37080
rect 27157 37077 27169 37080
rect 27203 37077 27215 37111
rect 27157 37071 27215 37077
rect 27798 37068 27804 37120
rect 27856 37108 27862 37120
rect 28077 37111 28135 37117
rect 28077 37108 28089 37111
rect 27856 37080 28089 37108
rect 27856 37068 27862 37080
rect 28077 37077 28089 37080
rect 28123 37077 28135 37111
rect 28718 37108 28724 37120
rect 28679 37080 28724 37108
rect 28077 37071 28135 37077
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 29730 37108 29736 37120
rect 29691 37080 29736 37108
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 31386 37108 31392 37120
rect 31347 37080 31392 37108
rect 31386 37068 31392 37080
rect 31444 37068 31450 37120
rect 33321 37111 33379 37117
rect 33321 37077 33333 37111
rect 33367 37108 33379 37111
rect 33686 37108 33692 37120
rect 33367 37080 33692 37108
rect 33367 37077 33379 37080
rect 33321 37071 33379 37077
rect 33686 37068 33692 37080
rect 33744 37068 33750 37120
rect 34606 37068 34612 37120
rect 34664 37108 34670 37120
rect 34793 37111 34851 37117
rect 34793 37108 34805 37111
rect 34664 37080 34805 37108
rect 34664 37068 34670 37080
rect 34793 37077 34805 37080
rect 34839 37077 34851 37111
rect 34793 37071 34851 37077
rect 34882 37068 34888 37120
rect 34940 37108 34946 37120
rect 35529 37111 35587 37117
rect 35529 37108 35541 37111
rect 34940 37080 35541 37108
rect 34940 37068 34946 37080
rect 35529 37077 35541 37080
rect 35575 37077 35587 37111
rect 36262 37108 36268 37120
rect 36223 37080 36268 37108
rect 35529 37071 35587 37077
rect 36262 37068 36268 37080
rect 36320 37068 36326 37120
rect 37476 37117 37504 37148
rect 38378 37136 38384 37148
rect 38436 37136 38442 37188
rect 37461 37111 37519 37117
rect 37461 37077 37473 37111
rect 37507 37077 37519 37111
rect 37461 37071 37519 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 2498 36864 2504 36916
rect 2556 36904 2562 36916
rect 3421 36907 3479 36913
rect 3421 36904 3433 36907
rect 2556 36876 3433 36904
rect 2556 36864 2562 36876
rect 3421 36873 3433 36876
rect 3467 36873 3479 36907
rect 3421 36867 3479 36873
rect 3602 36864 3608 36916
rect 3660 36904 3666 36916
rect 4065 36907 4123 36913
rect 4065 36904 4077 36907
rect 3660 36876 4077 36904
rect 3660 36864 3666 36876
rect 4065 36873 4077 36876
rect 4111 36873 4123 36907
rect 4065 36867 4123 36873
rect 4614 36864 4620 36916
rect 4672 36904 4678 36916
rect 4801 36907 4859 36913
rect 4801 36904 4813 36907
rect 4672 36876 4813 36904
rect 4672 36864 4678 36876
rect 4801 36873 4813 36876
rect 4847 36873 4859 36907
rect 4801 36867 4859 36873
rect 4982 36864 4988 36916
rect 5040 36904 5046 36916
rect 5629 36907 5687 36913
rect 5629 36904 5641 36907
rect 5040 36876 5641 36904
rect 5040 36864 5046 36876
rect 5629 36873 5641 36876
rect 5675 36873 5687 36907
rect 5629 36867 5687 36873
rect 5810 36864 5816 36916
rect 5868 36904 5874 36916
rect 7285 36907 7343 36913
rect 7285 36904 7297 36907
rect 5868 36876 7297 36904
rect 5868 36864 5874 36876
rect 7285 36873 7297 36876
rect 7331 36873 7343 36907
rect 7285 36867 7343 36873
rect 7742 36864 7748 36916
rect 7800 36904 7806 36916
rect 8757 36907 8815 36913
rect 8757 36904 8769 36907
rect 7800 36876 8769 36904
rect 7800 36864 7806 36876
rect 8757 36873 8769 36876
rect 8803 36873 8815 36907
rect 8757 36867 8815 36873
rect 8846 36864 8852 36916
rect 8904 36904 8910 36916
rect 9401 36907 9459 36913
rect 9401 36904 9413 36907
rect 8904 36876 9413 36904
rect 8904 36864 8910 36876
rect 9401 36873 9413 36876
rect 9447 36873 9459 36907
rect 9401 36867 9459 36873
rect 10873 36907 10931 36913
rect 10873 36873 10885 36907
rect 10919 36904 10931 36907
rect 10962 36904 10968 36916
rect 10919 36876 10968 36904
rect 10919 36873 10931 36876
rect 10873 36867 10931 36873
rect 10962 36864 10968 36876
rect 11020 36864 11026 36916
rect 11974 36864 11980 36916
rect 12032 36904 12038 36916
rect 12161 36907 12219 36913
rect 12161 36904 12173 36907
rect 12032 36876 12173 36904
rect 12032 36864 12038 36876
rect 12161 36873 12173 36876
rect 12207 36873 12219 36907
rect 12161 36867 12219 36873
rect 13078 36864 13084 36916
rect 13136 36904 13142 36916
rect 13633 36907 13691 36913
rect 13633 36904 13645 36907
rect 13136 36876 13645 36904
rect 13136 36864 13142 36876
rect 13633 36873 13645 36876
rect 13679 36873 13691 36907
rect 13633 36867 13691 36873
rect 14090 36864 14096 36916
rect 14148 36904 14154 36916
rect 14461 36907 14519 36913
rect 14461 36904 14473 36907
rect 14148 36876 14473 36904
rect 14148 36864 14154 36876
rect 14461 36873 14473 36876
rect 14507 36873 14519 36907
rect 14461 36867 14519 36873
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 15749 36907 15807 36913
rect 15749 36904 15761 36907
rect 15252 36876 15761 36904
rect 15252 36864 15258 36876
rect 15749 36873 15761 36876
rect 15795 36873 15807 36907
rect 15749 36867 15807 36873
rect 17218 36864 17224 36916
rect 17276 36904 17282 36916
rect 17865 36907 17923 36913
rect 17865 36904 17877 36907
rect 17276 36876 17877 36904
rect 17276 36864 17282 36876
rect 17865 36873 17877 36876
rect 17911 36873 17923 36907
rect 17865 36867 17923 36873
rect 18322 36864 18328 36916
rect 18380 36904 18386 36916
rect 18601 36907 18659 36913
rect 18601 36904 18613 36907
rect 18380 36876 18613 36904
rect 18380 36864 18386 36876
rect 18601 36873 18613 36876
rect 18647 36873 18659 36907
rect 18601 36867 18659 36873
rect 19334 36864 19340 36916
rect 19392 36904 19398 36916
rect 19521 36907 19579 36913
rect 19521 36904 19533 36907
rect 19392 36876 19533 36904
rect 19392 36864 19398 36876
rect 19521 36873 19533 36876
rect 19567 36873 19579 36907
rect 19521 36867 19579 36873
rect 19978 36864 19984 36916
rect 20036 36904 20042 36916
rect 20257 36907 20315 36913
rect 20257 36904 20269 36907
rect 20036 36876 20269 36904
rect 20036 36864 20042 36876
rect 20257 36873 20269 36876
rect 20303 36873 20315 36907
rect 20257 36867 20315 36873
rect 20806 36864 20812 36916
rect 20864 36904 20870 36916
rect 21085 36907 21143 36913
rect 21085 36904 21097 36907
rect 20864 36876 21097 36904
rect 20864 36864 20870 36876
rect 21085 36873 21097 36876
rect 21131 36873 21143 36907
rect 21085 36867 21143 36873
rect 21450 36864 21456 36916
rect 21508 36904 21514 36916
rect 22005 36907 22063 36913
rect 22005 36904 22017 36907
rect 21508 36876 22017 36904
rect 21508 36864 21514 36876
rect 22005 36873 22017 36876
rect 22051 36873 22063 36907
rect 22005 36867 22063 36873
rect 22554 36864 22560 36916
rect 22612 36904 22618 36916
rect 22741 36907 22799 36913
rect 22741 36904 22753 36907
rect 22612 36876 22753 36904
rect 22612 36864 22618 36876
rect 22741 36873 22753 36876
rect 22787 36873 22799 36907
rect 22741 36867 22799 36873
rect 23566 36864 23572 36916
rect 23624 36904 23630 36916
rect 24213 36907 24271 36913
rect 24213 36904 24225 36907
rect 23624 36876 24225 36904
rect 23624 36864 23630 36876
rect 24213 36873 24225 36876
rect 24259 36873 24271 36907
rect 24213 36867 24271 36873
rect 24854 36864 24860 36916
rect 24912 36904 24918 36916
rect 24949 36907 25007 36913
rect 24949 36904 24961 36907
rect 24912 36876 24961 36904
rect 24912 36864 24918 36876
rect 24949 36873 24961 36876
rect 24995 36873 25007 36907
rect 24949 36867 25007 36873
rect 25038 36864 25044 36916
rect 25096 36904 25102 36916
rect 25685 36907 25743 36913
rect 25685 36904 25697 36907
rect 25096 36876 25697 36904
rect 25096 36864 25102 36876
rect 25685 36873 25697 36876
rect 25731 36873 25743 36907
rect 25685 36867 25743 36873
rect 26234 36864 26240 36916
rect 26292 36904 26298 36916
rect 27157 36907 27215 36913
rect 27157 36904 27169 36907
rect 26292 36876 27169 36904
rect 26292 36864 26298 36876
rect 27157 36873 27169 36876
rect 27203 36873 27215 36907
rect 27157 36867 27215 36873
rect 27338 36864 27344 36916
rect 27396 36904 27402 36916
rect 27893 36907 27951 36913
rect 27893 36904 27905 36907
rect 27396 36876 27905 36904
rect 27396 36864 27402 36876
rect 27893 36873 27905 36876
rect 27939 36873 27951 36907
rect 27893 36867 27951 36873
rect 28166 36864 28172 36916
rect 28224 36904 28230 36916
rect 28537 36907 28595 36913
rect 28537 36904 28549 36907
rect 28224 36876 28549 36904
rect 28224 36864 28230 36876
rect 28537 36873 28549 36876
rect 28583 36873 28595 36907
rect 28537 36867 28595 36873
rect 29178 36864 29184 36916
rect 29236 36904 29242 36916
rect 29457 36907 29515 36913
rect 29457 36904 29469 36907
rect 29236 36876 29469 36904
rect 29236 36864 29242 36876
rect 29457 36873 29469 36876
rect 29503 36873 29515 36907
rect 29457 36867 29515 36873
rect 29914 36864 29920 36916
rect 29972 36904 29978 36916
rect 30193 36907 30251 36913
rect 30193 36904 30205 36907
rect 29972 36876 30205 36904
rect 29972 36864 29978 36876
rect 30193 36873 30205 36876
rect 30239 36873 30251 36907
rect 30193 36867 30251 36873
rect 30926 36864 30932 36916
rect 30984 36904 30990 36916
rect 31205 36907 31263 36913
rect 31205 36904 31217 36907
rect 30984 36876 31217 36904
rect 30984 36864 30990 36876
rect 31205 36873 31217 36876
rect 31251 36873 31263 36907
rect 31205 36867 31263 36873
rect 32030 36864 32036 36916
rect 32088 36904 32094 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 32088 36876 32321 36904
rect 32088 36864 32094 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 33134 36864 33140 36916
rect 33192 36904 33198 36916
rect 33321 36907 33379 36913
rect 33321 36904 33333 36907
rect 33192 36876 33333 36904
rect 33192 36864 33198 36876
rect 33321 36873 33333 36876
rect 33367 36873 33379 36907
rect 33321 36867 33379 36873
rect 34146 36864 34152 36916
rect 34204 36904 34210 36916
rect 34425 36907 34483 36913
rect 34425 36904 34437 36907
rect 34204 36876 34437 36904
rect 34204 36864 34210 36876
rect 34425 36873 34437 36876
rect 34471 36873 34483 36907
rect 34425 36867 34483 36873
rect 34790 36864 34796 36916
rect 34848 36904 34854 36916
rect 34848 36876 35296 36904
rect 34848 36864 34854 36876
rect 106 36796 112 36848
rect 164 36836 170 36848
rect 1578 36836 1584 36848
rect 164 36808 1584 36836
rect 164 36796 170 36808
rect 1578 36796 1584 36808
rect 1636 36836 1642 36848
rect 1857 36839 1915 36845
rect 1857 36836 1869 36839
rect 1636 36808 1869 36836
rect 1636 36796 1642 36808
rect 1857 36805 1869 36808
rect 1903 36805 1915 36839
rect 1857 36799 1915 36805
rect 7466 36796 7472 36848
rect 7524 36836 7530 36848
rect 10045 36839 10103 36845
rect 10045 36836 10057 36839
rect 7524 36808 10057 36836
rect 7524 36796 7530 36808
rect 10045 36805 10057 36808
rect 10091 36805 10103 36839
rect 10045 36799 10103 36805
rect 12710 36796 12716 36848
rect 12768 36836 12774 36848
rect 12897 36839 12955 36845
rect 12897 36836 12909 36839
rect 12768 36808 12909 36836
rect 12768 36796 12774 36808
rect 12897 36805 12909 36808
rect 12943 36805 12955 36839
rect 12897 36799 12955 36805
rect 13722 36796 13728 36848
rect 13780 36836 13786 36848
rect 15013 36839 15071 36845
rect 15013 36836 15025 36839
rect 13780 36808 15025 36836
rect 13780 36796 13786 36808
rect 15013 36805 15025 36808
rect 15059 36805 15071 36839
rect 15013 36799 15071 36805
rect 16942 36796 16948 36848
rect 17000 36836 17006 36848
rect 17129 36839 17187 36845
rect 17129 36836 17141 36839
rect 17000 36808 17141 36836
rect 17000 36796 17006 36808
rect 17129 36805 17141 36808
rect 17175 36805 17187 36839
rect 17129 36799 17187 36805
rect 22830 36796 22836 36848
rect 22888 36836 22894 36848
rect 31386 36836 31392 36848
rect 22888 36808 31392 36836
rect 22888 36796 22894 36808
rect 31386 36796 31392 36808
rect 31444 36796 31450 36848
rect 34330 36796 34336 36848
rect 34388 36836 34394 36848
rect 34882 36836 34888 36848
rect 34388 36808 34888 36836
rect 34388 36796 34394 36808
rect 34882 36796 34888 36808
rect 34940 36796 34946 36848
rect 35268 36836 35296 36876
rect 35342 36864 35348 36916
rect 35400 36904 35406 36916
rect 35437 36907 35495 36913
rect 35437 36904 35449 36907
rect 35400 36876 35449 36904
rect 35400 36864 35406 36876
rect 35437 36873 35449 36876
rect 35483 36873 35495 36907
rect 35437 36867 35495 36873
rect 36354 36864 36360 36916
rect 36412 36904 36418 36916
rect 36541 36907 36599 36913
rect 36541 36904 36553 36907
rect 36412 36876 36553 36904
rect 36412 36864 36418 36876
rect 36541 36873 36553 36876
rect 36587 36873 36599 36907
rect 36541 36867 36599 36873
rect 35710 36836 35716 36848
rect 35268 36808 35716 36836
rect 35710 36796 35716 36808
rect 35768 36836 35774 36848
rect 37277 36839 37335 36845
rect 37277 36836 37289 36839
rect 35768 36808 37289 36836
rect 35768 36796 35774 36808
rect 37277 36805 37289 36808
rect 37323 36805 37335 36839
rect 37277 36799 37335 36805
rect 37921 36839 37979 36845
rect 37921 36805 37933 36839
rect 37967 36836 37979 36839
rect 38010 36836 38016 36848
rect 37967 36808 38016 36836
rect 37967 36805 37979 36808
rect 37921 36799 37979 36805
rect 38010 36796 38016 36808
rect 38068 36796 38074 36848
rect 2774 36768 2780 36780
rect 2735 36740 2780 36768
rect 2774 36728 2780 36740
rect 2832 36728 2838 36780
rect 3234 36768 3240 36780
rect 3195 36740 3240 36768
rect 3234 36728 3240 36740
rect 3292 36728 3298 36780
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36768 4307 36771
rect 4614 36768 4620 36780
rect 4295 36740 4620 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 4985 36771 5043 36777
rect 4985 36737 4997 36771
rect 5031 36768 5043 36771
rect 5350 36768 5356 36780
rect 5031 36740 5356 36768
rect 5031 36737 5043 36740
rect 4985 36731 5043 36737
rect 5350 36728 5356 36740
rect 5408 36728 5414 36780
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 5534 36768 5540 36780
rect 5491 36740 5540 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 5534 36728 5540 36740
rect 5592 36728 5598 36780
rect 5626 36728 5632 36780
rect 5684 36768 5690 36780
rect 6178 36768 6184 36780
rect 5684 36740 6184 36768
rect 5684 36728 5690 36740
rect 6178 36728 6184 36740
rect 6236 36768 6242 36780
rect 6457 36771 6515 36777
rect 6457 36768 6469 36771
rect 6236 36740 6469 36768
rect 6236 36728 6242 36740
rect 6457 36737 6469 36740
rect 6503 36737 6515 36771
rect 7098 36768 7104 36780
rect 7059 36740 7104 36768
rect 6457 36731 6515 36737
rect 7098 36728 7104 36740
rect 7156 36728 7162 36780
rect 7926 36728 7932 36780
rect 7984 36768 7990 36780
rect 8113 36771 8171 36777
rect 8113 36768 8125 36771
rect 7984 36740 8125 36768
rect 7984 36728 7990 36740
rect 8113 36737 8125 36740
rect 8159 36737 8171 36771
rect 8570 36768 8576 36780
rect 8531 36740 8576 36768
rect 8113 36731 8171 36737
rect 8570 36728 8576 36740
rect 8628 36728 8634 36780
rect 9585 36771 9643 36777
rect 9585 36737 9597 36771
rect 9631 36768 9643 36771
rect 9766 36768 9772 36780
rect 9631 36740 9772 36768
rect 9631 36737 9643 36740
rect 9585 36731 9643 36737
rect 9766 36728 9772 36740
rect 9824 36728 9830 36780
rect 10686 36768 10692 36780
rect 10647 36740 10692 36768
rect 10686 36728 10692 36740
rect 10744 36728 10750 36780
rect 12345 36771 12403 36777
rect 12345 36737 12357 36771
rect 12391 36768 12403 36771
rect 13354 36768 13360 36780
rect 12391 36740 13360 36768
rect 12391 36737 12403 36740
rect 12345 36731 12403 36737
rect 13354 36728 13360 36740
rect 13412 36728 13418 36780
rect 13817 36771 13875 36777
rect 13817 36737 13829 36771
rect 13863 36737 13875 36771
rect 14274 36768 14280 36780
rect 14235 36740 14280 36768
rect 13817 36731 13875 36737
rect 9398 36660 9404 36712
rect 9456 36700 9462 36712
rect 11517 36703 11575 36709
rect 11517 36700 11529 36703
rect 9456 36672 11529 36700
rect 9456 36660 9462 36672
rect 11517 36669 11529 36672
rect 11563 36669 11575 36703
rect 13832 36700 13860 36731
rect 14274 36728 14280 36740
rect 14332 36728 14338 36780
rect 15933 36771 15991 36777
rect 15933 36737 15945 36771
rect 15979 36768 15991 36771
rect 16666 36768 16672 36780
rect 15979 36740 16672 36768
rect 15979 36737 15991 36740
rect 15933 36731 15991 36737
rect 16666 36728 16672 36740
rect 16724 36728 16730 36780
rect 18046 36768 18052 36780
rect 18007 36740 18052 36768
rect 18046 36728 18052 36740
rect 18104 36728 18110 36780
rect 18785 36771 18843 36777
rect 18785 36737 18797 36771
rect 18831 36768 18843 36771
rect 19426 36768 19432 36780
rect 18831 36740 19432 36768
rect 18831 36737 18843 36740
rect 18785 36731 18843 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 19705 36771 19763 36777
rect 19705 36737 19717 36771
rect 19751 36768 19763 36771
rect 20162 36768 20168 36780
rect 19751 36740 20168 36768
rect 19751 36737 19763 36740
rect 19705 36731 19763 36737
rect 20162 36728 20168 36740
rect 20220 36728 20226 36780
rect 20438 36768 20444 36780
rect 20399 36740 20444 36768
rect 20438 36728 20444 36740
rect 20496 36728 20502 36780
rect 20530 36728 20536 36780
rect 20588 36768 20594 36780
rect 20901 36771 20959 36777
rect 20901 36768 20913 36771
rect 20588 36740 20913 36768
rect 20588 36728 20594 36740
rect 20901 36737 20913 36740
rect 20947 36737 20959 36771
rect 20901 36731 20959 36737
rect 20990 36728 20996 36780
rect 21048 36768 21054 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21048 36740 21833 36768
rect 21048 36728 21054 36740
rect 21821 36737 21833 36740
rect 21867 36737 21879 36771
rect 22554 36768 22560 36780
rect 22515 36740 22560 36768
rect 21821 36731 21879 36737
rect 22554 36728 22560 36740
rect 22612 36728 22618 36780
rect 23198 36728 23204 36780
rect 23256 36768 23262 36780
rect 23474 36768 23480 36780
rect 23256 36740 23480 36768
rect 23256 36728 23262 36740
rect 23474 36728 23480 36740
rect 23532 36768 23538 36780
rect 23569 36771 23627 36777
rect 23569 36768 23581 36771
rect 23532 36740 23581 36768
rect 23532 36728 23538 36740
rect 23569 36737 23581 36740
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 23750 36728 23756 36780
rect 23808 36768 23814 36780
rect 24029 36771 24087 36777
rect 24029 36768 24041 36771
rect 23808 36740 24041 36768
rect 23808 36728 23814 36740
rect 24029 36737 24041 36740
rect 24075 36737 24087 36771
rect 24029 36731 24087 36737
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36737 24823 36771
rect 24765 36731 24823 36737
rect 14826 36700 14832 36712
rect 13832 36672 14832 36700
rect 11517 36663 11575 36669
rect 14826 36660 14832 36672
rect 14884 36660 14890 36712
rect 15378 36660 15384 36712
rect 15436 36700 15442 36712
rect 24780 36700 24808 36731
rect 25406 36728 25412 36780
rect 25464 36768 25470 36780
rect 25501 36771 25559 36777
rect 25501 36768 25513 36771
rect 25464 36740 25513 36768
rect 25464 36728 25470 36740
rect 25501 36737 25513 36740
rect 25547 36737 25559 36771
rect 26418 36768 26424 36780
rect 26379 36740 26424 36768
rect 25501 36731 25559 36737
rect 26418 36728 26424 36740
rect 26476 36728 26482 36780
rect 26878 36728 26884 36780
rect 26936 36768 26942 36780
rect 26973 36771 27031 36777
rect 26973 36768 26985 36771
rect 26936 36740 26985 36768
rect 26936 36728 26942 36740
rect 26973 36737 26985 36740
rect 27019 36737 27031 36771
rect 26973 36731 27031 36737
rect 27246 36728 27252 36780
rect 27304 36768 27310 36780
rect 27709 36771 27767 36777
rect 27709 36768 27721 36771
rect 27304 36740 27721 36768
rect 27304 36728 27310 36740
rect 27709 36737 27721 36740
rect 27755 36737 27767 36771
rect 27709 36731 27767 36737
rect 28626 36728 28632 36780
rect 28684 36768 28690 36780
rect 28721 36771 28779 36777
rect 28721 36768 28733 36771
rect 28684 36740 28733 36768
rect 28684 36728 28690 36740
rect 28721 36737 28733 36740
rect 28767 36737 28779 36771
rect 28721 36731 28779 36737
rect 29273 36771 29331 36777
rect 29273 36737 29285 36771
rect 29319 36737 29331 36771
rect 29273 36731 29331 36737
rect 15436 36672 24808 36700
rect 15436 36660 15442 36672
rect 28166 36660 28172 36712
rect 28224 36700 28230 36712
rect 29288 36700 29316 36731
rect 29362 36728 29368 36780
rect 29420 36768 29426 36780
rect 30009 36771 30067 36777
rect 30009 36768 30021 36771
rect 29420 36740 30021 36768
rect 29420 36728 29426 36740
rect 30009 36737 30021 36740
rect 30055 36737 30067 36771
rect 31018 36768 31024 36780
rect 30979 36740 31024 36768
rect 30009 36731 30067 36737
rect 31018 36728 31024 36740
rect 31076 36728 31082 36780
rect 31938 36728 31944 36780
rect 31996 36768 32002 36780
rect 32125 36771 32183 36777
rect 32125 36768 32137 36771
rect 31996 36740 32137 36768
rect 31996 36728 32002 36740
rect 32125 36737 32137 36740
rect 32171 36737 32183 36771
rect 33134 36768 33140 36780
rect 33095 36740 33140 36768
rect 32125 36731 32183 36737
rect 33134 36728 33140 36740
rect 33192 36728 33198 36780
rect 34238 36768 34244 36780
rect 34199 36740 34244 36768
rect 34238 36728 34244 36740
rect 34296 36728 34302 36780
rect 34790 36728 34796 36780
rect 34848 36768 34854 36780
rect 35253 36771 35311 36777
rect 35253 36768 35265 36771
rect 34848 36740 35265 36768
rect 34848 36728 34854 36740
rect 35253 36737 35265 36740
rect 35299 36737 35311 36771
rect 35253 36731 35311 36737
rect 36170 36728 36176 36780
rect 36228 36768 36234 36780
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 36228 36740 36369 36768
rect 36228 36728 36234 36740
rect 36357 36737 36369 36740
rect 36403 36737 36415 36771
rect 36357 36731 36415 36737
rect 28224 36672 29316 36700
rect 28224 36660 28230 36672
rect 2038 36632 2044 36644
rect 1999 36604 2044 36632
rect 2038 36592 2044 36604
rect 2096 36592 2102 36644
rect 6638 36632 6644 36644
rect 6599 36604 6644 36632
rect 6638 36592 6644 36604
rect 6696 36592 6702 36644
rect 6914 36592 6920 36644
rect 6972 36632 6978 36644
rect 7929 36635 7987 36641
rect 7929 36632 7941 36635
rect 6972 36604 7941 36632
rect 6972 36592 6978 36604
rect 7929 36601 7941 36604
rect 7975 36601 7987 36635
rect 7929 36595 7987 36601
rect 13081 36635 13139 36641
rect 13081 36601 13093 36635
rect 13127 36632 13139 36635
rect 13630 36632 13636 36644
rect 13127 36604 13636 36632
rect 13127 36601 13139 36604
rect 13081 36595 13139 36601
rect 13630 36592 13636 36604
rect 13688 36592 13694 36644
rect 18046 36592 18052 36644
rect 18104 36632 18110 36644
rect 18598 36632 18604 36644
rect 18104 36604 18604 36632
rect 18104 36592 18110 36604
rect 18598 36592 18604 36604
rect 18656 36632 18662 36644
rect 37550 36632 37556 36644
rect 18656 36604 37556 36632
rect 18656 36592 18662 36604
rect 37550 36592 37556 36604
rect 37608 36592 37614 36644
rect 38105 36635 38163 36641
rect 38105 36601 38117 36635
rect 38151 36632 38163 36635
rect 38562 36632 38568 36644
rect 38151 36604 38568 36632
rect 38151 36601 38163 36604
rect 38105 36595 38163 36601
rect 38562 36592 38568 36604
rect 38620 36592 38626 36644
rect 1486 36524 1492 36576
rect 1544 36564 1550 36576
rect 2593 36567 2651 36573
rect 2593 36564 2605 36567
rect 1544 36536 2605 36564
rect 1544 36524 1550 36536
rect 2593 36533 2605 36536
rect 2639 36533 2651 36567
rect 2593 36527 2651 36533
rect 6362 36524 6368 36576
rect 6420 36564 6426 36576
rect 6730 36564 6736 36576
rect 6420 36536 6736 36564
rect 6420 36524 6426 36536
rect 6730 36524 6736 36536
rect 6788 36524 6794 36576
rect 17218 36564 17224 36576
rect 17179 36536 17224 36564
rect 17218 36524 17224 36536
rect 17276 36524 17282 36576
rect 23382 36564 23388 36576
rect 23343 36536 23388 36564
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 26234 36524 26240 36576
rect 26292 36564 26298 36576
rect 26292 36536 26337 36564
rect 26292 36524 26298 36536
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 382 36320 388 36372
rect 440 36360 446 36372
rect 1489 36363 1547 36369
rect 1489 36360 1501 36363
rect 440 36332 1501 36360
rect 440 36320 446 36332
rect 1489 36329 1501 36332
rect 1535 36329 1547 36363
rect 1489 36323 1547 36329
rect 1854 36320 1860 36372
rect 1912 36360 1918 36372
rect 2225 36363 2283 36369
rect 2225 36360 2237 36363
rect 1912 36332 2237 36360
rect 1912 36320 1918 36332
rect 2225 36329 2237 36332
rect 2271 36329 2283 36363
rect 2225 36323 2283 36329
rect 2866 36320 2872 36372
rect 2924 36360 2930 36372
rect 3053 36363 3111 36369
rect 3053 36360 3065 36363
rect 2924 36332 3065 36360
rect 2924 36320 2930 36332
rect 3053 36329 3065 36332
rect 3099 36329 3111 36363
rect 3053 36323 3111 36329
rect 3878 36320 3884 36372
rect 3936 36360 3942 36372
rect 4065 36363 4123 36369
rect 4065 36360 4077 36363
rect 3936 36332 4077 36360
rect 3936 36320 3942 36332
rect 4065 36329 4077 36332
rect 4111 36329 4123 36363
rect 5350 36360 5356 36372
rect 5311 36332 5356 36360
rect 4065 36323 4123 36329
rect 5350 36320 5356 36332
rect 5408 36320 5414 36372
rect 5994 36320 6000 36372
rect 6052 36360 6058 36372
rect 6181 36363 6239 36369
rect 6181 36360 6193 36363
rect 6052 36332 6193 36360
rect 6052 36320 6058 36332
rect 6181 36329 6193 36332
rect 6227 36329 6239 36363
rect 6181 36323 6239 36329
rect 7190 36320 7196 36372
rect 7248 36360 7254 36372
rect 7285 36363 7343 36369
rect 7285 36360 7297 36363
rect 7248 36332 7297 36360
rect 7248 36320 7254 36332
rect 7285 36329 7297 36332
rect 7331 36329 7343 36363
rect 7926 36360 7932 36372
rect 7887 36332 7932 36360
rect 7285 36323 7343 36329
rect 7926 36320 7932 36332
rect 7984 36320 7990 36372
rect 8294 36320 8300 36372
rect 8352 36360 8358 36372
rect 9033 36363 9091 36369
rect 9033 36360 9045 36363
rect 8352 36332 9045 36360
rect 8352 36320 8358 36332
rect 9033 36329 9045 36332
rect 9079 36329 9091 36363
rect 9033 36323 9091 36329
rect 9858 36320 9864 36372
rect 9916 36360 9922 36372
rect 10045 36363 10103 36369
rect 10045 36360 10057 36363
rect 9916 36332 10057 36360
rect 9916 36320 9922 36332
rect 10045 36329 10057 36332
rect 10091 36329 10103 36363
rect 10045 36323 10103 36329
rect 10226 36320 10232 36372
rect 10284 36360 10290 36372
rect 10781 36363 10839 36369
rect 10781 36360 10793 36363
rect 10284 36332 10793 36360
rect 10284 36320 10290 36332
rect 10781 36329 10793 36332
rect 10827 36329 10839 36363
rect 10781 36323 10839 36329
rect 11330 36320 11336 36372
rect 11388 36360 11394 36372
rect 11517 36363 11575 36369
rect 11517 36360 11529 36363
rect 11388 36332 11529 36360
rect 11388 36320 11394 36332
rect 11517 36329 11529 36332
rect 11563 36329 11575 36363
rect 11517 36323 11575 36329
rect 12434 36320 12440 36372
rect 12492 36360 12498 36372
rect 12529 36363 12587 36369
rect 12529 36360 12541 36363
rect 12492 36332 12541 36360
rect 12492 36320 12498 36332
rect 12529 36329 12541 36332
rect 12575 36329 12587 36363
rect 12529 36323 12587 36329
rect 13446 36320 13452 36372
rect 13504 36360 13510 36372
rect 14277 36363 14335 36369
rect 14277 36360 14289 36363
rect 13504 36332 14289 36360
rect 13504 36320 13510 36332
rect 14277 36329 14289 36332
rect 14323 36329 14335 36363
rect 14277 36323 14335 36329
rect 14458 36320 14464 36372
rect 14516 36360 14522 36372
rect 15197 36363 15255 36369
rect 15197 36360 15209 36363
rect 14516 36332 15209 36360
rect 14516 36320 14522 36332
rect 15197 36329 15209 36332
rect 15243 36329 15255 36363
rect 15197 36323 15255 36329
rect 15933 36363 15991 36369
rect 15933 36329 15945 36363
rect 15979 36360 15991 36363
rect 16206 36360 16212 36372
rect 15979 36332 16212 36360
rect 15979 36329 15991 36332
rect 15933 36323 15991 36329
rect 16206 36320 16212 36332
rect 16264 36320 16270 36372
rect 16574 36320 16580 36372
rect 16632 36360 16638 36372
rect 16761 36363 16819 36369
rect 16761 36360 16773 36363
rect 16632 36332 16773 36360
rect 16632 36320 16638 36332
rect 16761 36329 16773 36332
rect 16807 36329 16819 36363
rect 16761 36323 16819 36329
rect 17586 36320 17592 36372
rect 17644 36360 17650 36372
rect 17773 36363 17831 36369
rect 17773 36360 17785 36363
rect 17644 36332 17785 36360
rect 17644 36320 17650 36332
rect 17773 36329 17785 36332
rect 17819 36329 17831 36363
rect 19334 36360 19340 36372
rect 19295 36332 19340 36360
rect 17773 36323 17831 36329
rect 19334 36320 19340 36332
rect 19392 36320 19398 36372
rect 20165 36363 20223 36369
rect 20165 36329 20177 36363
rect 20211 36360 20223 36363
rect 20530 36360 20536 36372
rect 20211 36332 20536 36360
rect 20211 36329 20223 36332
rect 20165 36323 20223 36329
rect 20530 36320 20536 36332
rect 20588 36320 20594 36372
rect 20809 36363 20867 36369
rect 20809 36329 20821 36363
rect 20855 36360 20867 36363
rect 20990 36360 20996 36372
rect 20855 36332 20996 36360
rect 20855 36329 20867 36332
rect 20809 36323 20867 36329
rect 20990 36320 20996 36332
rect 21048 36320 21054 36372
rect 21729 36363 21787 36369
rect 21729 36329 21741 36363
rect 21775 36360 21787 36363
rect 21818 36360 21824 36372
rect 21775 36332 21824 36360
rect 21775 36329 21787 36332
rect 21729 36323 21787 36329
rect 21818 36320 21824 36332
rect 21876 36320 21882 36372
rect 23750 36360 23756 36372
rect 21928 36332 23756 36360
rect 13541 36295 13599 36301
rect 13541 36261 13553 36295
rect 13587 36292 13599 36295
rect 21928 36292 21956 36332
rect 23750 36320 23756 36332
rect 23808 36320 23814 36372
rect 23934 36320 23940 36372
rect 23992 36360 23998 36372
rect 24489 36363 24547 36369
rect 24489 36360 24501 36363
rect 23992 36332 24501 36360
rect 23992 36320 23998 36332
rect 24489 36329 24501 36332
rect 24535 36329 24547 36363
rect 25314 36360 25320 36372
rect 25275 36332 25320 36360
rect 24489 36323 24547 36329
rect 25314 36320 25320 36332
rect 25372 36320 25378 36372
rect 25961 36363 26019 36369
rect 25961 36329 25973 36363
rect 26007 36360 26019 36363
rect 26418 36360 26424 36372
rect 26007 36332 26424 36360
rect 26007 36329 26019 36332
rect 25961 36323 26019 36329
rect 26418 36320 26424 36332
rect 26476 36320 26482 36372
rect 26605 36363 26663 36369
rect 26605 36329 26617 36363
rect 26651 36360 26663 36363
rect 27062 36360 27068 36372
rect 26651 36332 27068 36360
rect 26651 36329 26663 36332
rect 26605 36323 26663 36329
rect 27062 36320 27068 36332
rect 27120 36320 27126 36372
rect 27246 36360 27252 36372
rect 27207 36332 27252 36360
rect 27246 36320 27252 36332
rect 27304 36320 27310 36372
rect 28166 36360 28172 36372
rect 28127 36332 28172 36360
rect 28166 36320 28172 36332
rect 28224 36320 28230 36372
rect 28626 36360 28632 36372
rect 28587 36332 28632 36360
rect 28626 36320 28632 36332
rect 28684 36320 28690 36372
rect 28902 36320 28908 36372
rect 28960 36360 28966 36372
rect 29549 36363 29607 36369
rect 29549 36360 29561 36363
rect 28960 36332 29561 36360
rect 28960 36320 28966 36332
rect 29549 36329 29561 36332
rect 29595 36329 29607 36363
rect 29549 36323 29607 36329
rect 31294 36320 31300 36372
rect 31352 36360 31358 36372
rect 31849 36363 31907 36369
rect 31849 36360 31861 36363
rect 31352 36332 31861 36360
rect 31352 36320 31358 36332
rect 31849 36329 31861 36332
rect 31895 36329 31907 36363
rect 31849 36323 31907 36329
rect 34514 36320 34520 36372
rect 34572 36360 34578 36372
rect 34885 36363 34943 36369
rect 34885 36360 34897 36363
rect 34572 36332 34897 36360
rect 34572 36320 34578 36332
rect 34885 36329 34897 36332
rect 34931 36329 34943 36363
rect 35434 36360 35440 36372
rect 35395 36332 35440 36360
rect 34885 36323 34943 36329
rect 35434 36320 35440 36332
rect 35492 36320 35498 36372
rect 13587 36264 21956 36292
rect 22741 36295 22799 36301
rect 13587 36261 13599 36264
rect 13541 36255 13599 36261
rect 22741 36261 22753 36295
rect 22787 36292 22799 36295
rect 22830 36292 22836 36304
rect 22787 36264 22836 36292
rect 22787 36261 22799 36264
rect 22741 36255 22799 36261
rect 22830 36252 22836 36264
rect 22888 36252 22894 36304
rect 23661 36295 23719 36301
rect 23661 36261 23673 36295
rect 23707 36292 23719 36295
rect 26234 36292 26240 36304
rect 23707 36264 26240 36292
rect 23707 36261 23719 36264
rect 23661 36255 23719 36261
rect 26234 36252 26240 36264
rect 26292 36252 26298 36304
rect 27890 36252 27896 36304
rect 27948 36292 27954 36304
rect 27948 36264 35894 36292
rect 27948 36252 27954 36264
rect 15286 36184 15292 36236
rect 15344 36224 15350 36236
rect 18417 36227 18475 36233
rect 18417 36224 18429 36227
rect 15344 36196 18429 36224
rect 15344 36184 15350 36196
rect 18417 36193 18429 36196
rect 18463 36193 18475 36227
rect 18417 36187 18475 36193
rect 19260 36196 28764 36224
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 2409 36159 2467 36165
rect 2409 36125 2421 36159
rect 2455 36125 2467 36159
rect 2409 36119 2467 36125
rect 2424 36088 2452 36119
rect 3050 36116 3056 36168
rect 3108 36156 3114 36168
rect 3237 36159 3295 36165
rect 3237 36156 3249 36159
rect 3108 36128 3249 36156
rect 3108 36116 3114 36128
rect 3237 36125 3249 36128
rect 3283 36125 3295 36159
rect 3237 36119 3295 36125
rect 4249 36159 4307 36165
rect 4249 36125 4261 36159
rect 4295 36156 4307 36159
rect 4982 36156 4988 36168
rect 4295 36128 4988 36156
rect 4295 36125 4307 36128
rect 4249 36119 4307 36125
rect 4982 36116 4988 36128
rect 5040 36116 5046 36168
rect 5537 36159 5595 36165
rect 5537 36125 5549 36159
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 6365 36159 6423 36165
rect 6365 36125 6377 36159
rect 6411 36156 6423 36159
rect 7006 36156 7012 36168
rect 6411 36128 7012 36156
rect 6411 36125 6423 36128
rect 6365 36119 6423 36125
rect 3142 36088 3148 36100
rect 2424 36060 3148 36088
rect 3142 36048 3148 36060
rect 3200 36048 3206 36100
rect 4893 36091 4951 36097
rect 4893 36057 4905 36091
rect 4939 36088 4951 36091
rect 5552 36088 5580 36119
rect 7006 36116 7012 36128
rect 7064 36116 7070 36168
rect 7466 36156 7472 36168
rect 7427 36128 7472 36156
rect 7466 36116 7472 36128
rect 7524 36116 7530 36168
rect 8018 36116 8024 36168
rect 8076 36156 8082 36168
rect 8113 36159 8171 36165
rect 8113 36156 8125 36159
rect 8076 36128 8125 36156
rect 8076 36116 8082 36128
rect 8113 36125 8125 36128
rect 8159 36125 8171 36159
rect 9214 36156 9220 36168
rect 9175 36128 9220 36156
rect 8113 36119 8171 36125
rect 9214 36116 9220 36128
rect 9272 36116 9278 36168
rect 10226 36156 10232 36168
rect 10187 36128 10232 36156
rect 10226 36116 10232 36128
rect 10284 36116 10290 36168
rect 10965 36159 11023 36165
rect 10965 36125 10977 36159
rect 11011 36125 11023 36159
rect 11698 36156 11704 36168
rect 11659 36128 11704 36156
rect 10965 36119 11023 36125
rect 6454 36088 6460 36100
rect 4939 36060 6460 36088
rect 4939 36057 4951 36060
rect 4893 36051 4951 36057
rect 6454 36048 6460 36060
rect 6512 36048 6518 36100
rect 10980 36088 11008 36119
rect 11698 36116 11704 36128
rect 11756 36116 11762 36168
rect 12713 36159 12771 36165
rect 12713 36125 12725 36159
rect 12759 36125 12771 36159
rect 12713 36119 12771 36125
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36156 13415 36159
rect 13446 36156 13452 36168
rect 13403 36128 13452 36156
rect 13403 36125 13415 36128
rect 13357 36119 13415 36125
rect 12250 36088 12256 36100
rect 10980 36060 12256 36088
rect 12250 36048 12256 36060
rect 12308 36048 12314 36100
rect 12728 36088 12756 36119
rect 13446 36116 13452 36128
rect 13504 36116 13510 36168
rect 13906 36116 13912 36168
rect 13964 36156 13970 36168
rect 14093 36159 14151 36165
rect 14093 36156 14105 36159
rect 13964 36128 14105 36156
rect 13964 36116 13970 36128
rect 14093 36125 14105 36128
rect 14139 36125 14151 36159
rect 14093 36119 14151 36125
rect 14550 36116 14556 36168
rect 14608 36156 14614 36168
rect 15013 36159 15071 36165
rect 15013 36156 15025 36159
rect 14608 36128 15025 36156
rect 14608 36116 14614 36128
rect 15013 36125 15025 36128
rect 15059 36125 15071 36159
rect 15013 36119 15071 36125
rect 16117 36159 16175 36165
rect 16117 36125 16129 36159
rect 16163 36156 16175 36159
rect 16850 36156 16856 36168
rect 16163 36128 16856 36156
rect 16163 36125 16175 36128
rect 16117 36119 16175 36125
rect 16850 36116 16856 36128
rect 16908 36116 16914 36168
rect 16945 36159 17003 36165
rect 16945 36125 16957 36159
rect 16991 36156 17003 36159
rect 17126 36156 17132 36168
rect 16991 36128 17132 36156
rect 16991 36125 17003 36128
rect 16945 36119 17003 36125
rect 17126 36116 17132 36128
rect 17184 36116 17190 36168
rect 17957 36159 18015 36165
rect 17957 36125 17969 36159
rect 18003 36156 18015 36159
rect 18046 36156 18052 36168
rect 18003 36128 18052 36156
rect 18003 36125 18015 36128
rect 17957 36119 18015 36125
rect 18046 36116 18052 36128
rect 18104 36116 18110 36168
rect 12894 36088 12900 36100
rect 12728 36060 12900 36088
rect 12894 36048 12900 36060
rect 12952 36088 12958 36100
rect 19260 36088 19288 36196
rect 19521 36159 19579 36165
rect 19521 36125 19533 36159
rect 19567 36125 19579 36159
rect 19978 36156 19984 36168
rect 19939 36128 19984 36156
rect 19521 36119 19579 36125
rect 12952 36060 19288 36088
rect 19536 36088 19564 36119
rect 19978 36116 19984 36128
rect 20036 36116 20042 36168
rect 20625 36159 20683 36165
rect 20625 36125 20637 36159
rect 20671 36156 20683 36159
rect 20714 36156 20720 36168
rect 20671 36128 20720 36156
rect 20671 36125 20683 36128
rect 20625 36119 20683 36125
rect 20714 36116 20720 36128
rect 20772 36116 20778 36168
rect 21910 36156 21916 36168
rect 21871 36128 21916 36156
rect 21910 36116 21916 36128
rect 21968 36116 21974 36168
rect 24673 36159 24731 36165
rect 22020 36128 23428 36156
rect 20254 36088 20260 36100
rect 19536 36060 20260 36088
rect 12952 36048 12958 36060
rect 20254 36048 20260 36060
rect 20312 36048 20318 36100
rect 18046 35980 18052 36032
rect 18104 36020 18110 36032
rect 22020 36020 22048 36128
rect 22373 36091 22431 36097
rect 22373 36057 22385 36091
rect 22419 36088 22431 36091
rect 23106 36088 23112 36100
rect 22419 36060 23112 36088
rect 22419 36057 22431 36060
rect 22373 36051 22431 36057
rect 23106 36048 23112 36060
rect 23164 36088 23170 36100
rect 23293 36091 23351 36097
rect 23293 36088 23305 36091
rect 23164 36060 23305 36088
rect 23164 36048 23170 36060
rect 23293 36057 23305 36060
rect 23339 36057 23351 36091
rect 23400 36088 23428 36128
rect 24673 36125 24685 36159
rect 24719 36156 24731 36159
rect 24854 36156 24860 36168
rect 24719 36128 24860 36156
rect 24719 36125 24731 36128
rect 24673 36119 24731 36125
rect 24854 36116 24860 36128
rect 24912 36116 24918 36168
rect 26445 36159 26503 36165
rect 26445 36125 26457 36159
rect 26491 36156 26503 36159
rect 26602 36156 26608 36168
rect 26491 36128 26608 36156
rect 26491 36125 26503 36128
rect 26445 36119 26503 36125
rect 26602 36116 26608 36128
rect 26660 36116 26666 36168
rect 27062 36156 27068 36168
rect 27023 36128 27068 36156
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 27985 36159 28043 36165
rect 27985 36125 27997 36159
rect 28031 36125 28043 36159
rect 27985 36119 28043 36125
rect 27890 36088 27896 36100
rect 23400 36060 27896 36088
rect 23293 36051 23351 36057
rect 27890 36048 27896 36060
rect 27948 36048 27954 36100
rect 18104 35992 22048 36020
rect 22833 36023 22891 36029
rect 18104 35980 18110 35992
rect 22833 35989 22845 36023
rect 22879 36020 22891 36023
rect 23198 36020 23204 36032
rect 22879 35992 23204 36020
rect 22879 35989 22891 35992
rect 22833 35983 22891 35989
rect 23198 35980 23204 35992
rect 23256 35980 23262 36032
rect 23658 35980 23664 36032
rect 23716 36020 23722 36032
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 23716 35992 23765 36020
rect 23716 35980 23722 35992
rect 23753 35989 23765 35992
rect 23799 35989 23811 36023
rect 23753 35983 23811 35989
rect 23842 35980 23848 36032
rect 23900 36020 23906 36032
rect 28000 36020 28028 36119
rect 28736 36088 28764 36196
rect 28994 36184 29000 36236
rect 29052 36224 29058 36236
rect 30929 36227 30987 36233
rect 30929 36224 30941 36227
rect 29052 36196 30941 36224
rect 29052 36184 29058 36196
rect 30929 36193 30941 36196
rect 30975 36193 30987 36227
rect 33321 36227 33379 36233
rect 33321 36224 33333 36227
rect 30929 36187 30987 36193
rect 31036 36196 33333 36224
rect 28813 36159 28871 36165
rect 28813 36125 28825 36159
rect 28859 36156 28871 36159
rect 29546 36156 29552 36168
rect 28859 36128 29552 36156
rect 28859 36125 28871 36128
rect 28813 36119 28871 36125
rect 29546 36116 29552 36128
rect 29604 36116 29610 36168
rect 30190 36156 30196 36168
rect 30151 36128 30196 36156
rect 30190 36116 30196 36128
rect 30248 36116 30254 36168
rect 31036 36156 31064 36196
rect 33321 36193 33333 36196
rect 33367 36193 33379 36227
rect 35866 36224 35894 36264
rect 36541 36227 36599 36233
rect 36541 36224 36553 36227
rect 35866 36196 36553 36224
rect 33321 36187 33379 36193
rect 36541 36193 36553 36196
rect 36587 36193 36599 36227
rect 36541 36187 36599 36193
rect 36817 36227 36875 36233
rect 36817 36193 36829 36227
rect 36863 36224 36875 36227
rect 37458 36224 37464 36236
rect 36863 36196 37464 36224
rect 36863 36193 36875 36196
rect 36817 36187 36875 36193
rect 37458 36184 37464 36196
rect 37516 36184 37522 36236
rect 37550 36184 37556 36236
rect 37608 36224 37614 36236
rect 37608 36196 37653 36224
rect 37608 36184 37614 36196
rect 31662 36156 31668 36168
rect 30300 36128 31064 36156
rect 31623 36128 31668 36156
rect 30300 36088 30328 36128
rect 31662 36116 31668 36128
rect 31720 36116 31726 36168
rect 34698 36156 34704 36168
rect 34659 36128 34704 36156
rect 34698 36116 34704 36128
rect 34756 36116 34762 36168
rect 37277 36159 37335 36165
rect 37277 36125 37289 36159
rect 37323 36156 37335 36159
rect 38470 36156 38476 36168
rect 37323 36128 38476 36156
rect 37323 36125 37335 36128
rect 37277 36119 37335 36125
rect 38470 36116 38476 36128
rect 38528 36116 38534 36168
rect 28736 36060 30328 36088
rect 30377 36091 30435 36097
rect 30377 36057 30389 36091
rect 30423 36088 30435 36091
rect 30466 36088 30472 36100
rect 30423 36060 30472 36088
rect 30423 36057 30435 36060
rect 30377 36051 30435 36057
rect 30466 36048 30472 36060
rect 30524 36048 30530 36100
rect 30926 36048 30932 36100
rect 30984 36088 30990 36100
rect 31113 36091 31171 36097
rect 31113 36088 31125 36091
rect 30984 36060 31125 36088
rect 30984 36048 30990 36060
rect 31113 36057 31125 36060
rect 31159 36057 31171 36091
rect 31113 36051 31171 36057
rect 32585 36091 32643 36097
rect 32585 36057 32597 36091
rect 32631 36088 32643 36091
rect 32674 36088 32680 36100
rect 32631 36060 32680 36088
rect 32631 36057 32643 36060
rect 32585 36051 32643 36057
rect 32674 36048 32680 36060
rect 32732 36048 32738 36100
rect 33505 36091 33563 36097
rect 33505 36057 33517 36091
rect 33551 36088 33563 36091
rect 34057 36091 34115 36097
rect 34057 36088 34069 36091
rect 33551 36060 34069 36088
rect 33551 36057 33563 36060
rect 33505 36051 33563 36057
rect 34057 36057 34069 36060
rect 34103 36088 34115 36091
rect 34146 36088 34152 36100
rect 34103 36060 34152 36088
rect 34103 36057 34115 36060
rect 34057 36051 34115 36057
rect 34146 36048 34152 36060
rect 34204 36048 34210 36100
rect 23900 35992 28028 36020
rect 23900 35980 23906 35992
rect 28442 35980 28448 36032
rect 28500 36020 28506 36032
rect 28902 36020 28908 36032
rect 28500 35992 28908 36020
rect 28500 35980 28506 35992
rect 28902 35980 28908 35992
rect 28960 35980 28966 36032
rect 30098 35980 30104 36032
rect 30156 36020 30162 36032
rect 32493 36023 32551 36029
rect 32493 36020 32505 36023
rect 30156 35992 32505 36020
rect 30156 35980 30162 35992
rect 32493 35989 32505 35992
rect 32539 35989 32551 36023
rect 32493 35983 32551 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 750 35776 756 35828
rect 808 35816 814 35828
rect 1489 35819 1547 35825
rect 1489 35816 1501 35819
rect 808 35788 1501 35816
rect 808 35776 814 35788
rect 1489 35785 1501 35788
rect 1535 35785 1547 35819
rect 1489 35779 1547 35785
rect 2685 35819 2743 35825
rect 2685 35785 2697 35819
rect 2731 35785 2743 35819
rect 2685 35779 2743 35785
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 2700 35680 2728 35779
rect 3142 35776 3148 35828
rect 3200 35816 3206 35828
rect 3329 35819 3387 35825
rect 3329 35816 3341 35819
rect 3200 35788 3341 35816
rect 3200 35776 3206 35788
rect 3329 35785 3341 35788
rect 3375 35785 3387 35819
rect 3329 35779 3387 35785
rect 4062 35776 4068 35828
rect 4120 35816 4126 35828
rect 4525 35819 4583 35825
rect 4525 35816 4537 35819
rect 4120 35788 4537 35816
rect 4120 35776 4126 35788
rect 4525 35785 4537 35788
rect 4571 35785 4583 35819
rect 4525 35779 4583 35785
rect 5169 35819 5227 35825
rect 5169 35785 5181 35819
rect 5215 35816 5227 35819
rect 5258 35816 5264 35828
rect 5215 35788 5264 35816
rect 5215 35785 5227 35788
rect 5169 35779 5227 35785
rect 5258 35776 5264 35788
rect 5316 35776 5322 35828
rect 6641 35819 6699 35825
rect 6641 35785 6653 35819
rect 6687 35816 6699 35819
rect 7098 35816 7104 35828
rect 6687 35788 7104 35816
rect 6687 35785 6699 35788
rect 6641 35779 6699 35785
rect 7098 35776 7104 35788
rect 7156 35776 7162 35828
rect 8570 35816 8576 35828
rect 8531 35788 8576 35816
rect 8570 35776 8576 35788
rect 8628 35776 8634 35828
rect 9306 35776 9312 35828
rect 9364 35816 9370 35828
rect 9769 35819 9827 35825
rect 9769 35816 9781 35819
rect 9364 35788 9781 35816
rect 9364 35776 9370 35788
rect 9769 35785 9781 35788
rect 9815 35785 9827 35819
rect 9769 35779 9827 35785
rect 10686 35776 10692 35828
rect 10744 35816 10750 35828
rect 10781 35819 10839 35825
rect 10781 35816 10793 35819
rect 10744 35788 10793 35816
rect 10744 35776 10750 35788
rect 10781 35785 10793 35788
rect 10827 35785 10839 35819
rect 10781 35779 10839 35785
rect 11698 35776 11704 35828
rect 11756 35816 11762 35828
rect 12253 35819 12311 35825
rect 12253 35816 12265 35819
rect 11756 35788 12265 35816
rect 11756 35776 11762 35788
rect 12253 35785 12265 35788
rect 12299 35785 12311 35819
rect 12253 35779 12311 35785
rect 14185 35819 14243 35825
rect 14185 35785 14197 35819
rect 14231 35816 14243 35819
rect 14274 35816 14280 35828
rect 14231 35788 14280 35816
rect 14231 35785 14243 35788
rect 14185 35779 14243 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 14826 35816 14832 35828
rect 14787 35788 14832 35816
rect 14826 35776 14832 35788
rect 14884 35776 14890 35828
rect 15470 35776 15476 35828
rect 15528 35816 15534 35828
rect 15657 35819 15715 35825
rect 15657 35816 15669 35819
rect 15528 35788 15669 35816
rect 15528 35776 15534 35788
rect 15657 35785 15669 35788
rect 15703 35785 15715 35819
rect 16666 35816 16672 35828
rect 16627 35788 16672 35816
rect 15657 35779 15715 35785
rect 16666 35776 16672 35788
rect 16724 35776 16730 35828
rect 16850 35776 16856 35828
rect 16908 35816 16914 35828
rect 17313 35819 17371 35825
rect 17313 35816 17325 35819
rect 16908 35788 17325 35816
rect 16908 35776 16914 35788
rect 17313 35785 17325 35788
rect 17359 35785 17371 35819
rect 17313 35779 17371 35785
rect 18690 35776 18696 35828
rect 18748 35816 18754 35828
rect 19334 35816 19340 35828
rect 18748 35788 19340 35816
rect 18748 35776 18754 35788
rect 19334 35776 19340 35788
rect 19392 35776 19398 35828
rect 19705 35819 19763 35825
rect 19705 35785 19717 35819
rect 19751 35816 19763 35819
rect 20898 35816 20904 35828
rect 19751 35788 20904 35816
rect 19751 35785 19763 35788
rect 19705 35779 19763 35785
rect 20898 35776 20904 35788
rect 20956 35776 20962 35828
rect 22186 35776 22192 35828
rect 22244 35816 22250 35828
rect 22465 35819 22523 35825
rect 22465 35816 22477 35819
rect 22244 35788 22477 35816
rect 22244 35776 22250 35788
rect 22465 35785 22477 35788
rect 22511 35785 22523 35819
rect 22465 35779 22523 35785
rect 22922 35776 22928 35828
rect 22980 35816 22986 35828
rect 23201 35819 23259 35825
rect 23201 35816 23213 35819
rect 22980 35788 23213 35816
rect 22980 35776 22986 35788
rect 23201 35785 23213 35788
rect 23247 35785 23259 35819
rect 23201 35779 23259 35785
rect 23474 35776 23480 35828
rect 23532 35816 23538 35828
rect 23753 35819 23811 35825
rect 23753 35816 23765 35819
rect 23532 35788 23765 35816
rect 23532 35776 23538 35788
rect 23753 35785 23765 35788
rect 23799 35785 23811 35819
rect 24302 35816 24308 35828
rect 24263 35788 24308 35816
rect 23753 35779 23811 35785
rect 24302 35776 24308 35788
rect 24360 35776 24366 35828
rect 26421 35819 26479 35825
rect 26421 35785 26433 35819
rect 26467 35816 26479 35819
rect 26970 35816 26976 35828
rect 26467 35788 26976 35816
rect 26467 35785 26479 35788
rect 26421 35779 26479 35785
rect 26970 35776 26976 35788
rect 27028 35776 27034 35828
rect 28810 35776 28816 35828
rect 28868 35816 28874 35828
rect 29730 35816 29736 35828
rect 28868 35788 29736 35816
rect 28868 35776 28874 35788
rect 29730 35776 29736 35788
rect 29788 35776 29794 35828
rect 30282 35776 30288 35828
rect 30340 35816 30346 35828
rect 30469 35819 30527 35825
rect 30469 35816 30481 35819
rect 30340 35788 30481 35816
rect 30340 35776 30346 35788
rect 30469 35785 30481 35788
rect 30515 35785 30527 35819
rect 31202 35816 31208 35828
rect 31163 35788 31208 35816
rect 30469 35779 30527 35785
rect 31202 35776 31208 35788
rect 31260 35776 31266 35828
rect 32398 35776 32404 35828
rect 32456 35816 32462 35828
rect 33413 35819 33471 35825
rect 33413 35816 33425 35819
rect 32456 35788 33425 35816
rect 32456 35776 32462 35788
rect 33413 35785 33425 35788
rect 33459 35785 33471 35819
rect 33413 35779 33471 35785
rect 35526 35776 35532 35828
rect 35584 35816 35590 35828
rect 35805 35819 35863 35825
rect 35805 35816 35817 35819
rect 35584 35788 35817 35816
rect 35584 35776 35590 35788
rect 35805 35785 35817 35788
rect 35851 35785 35863 35819
rect 37274 35816 37280 35828
rect 37235 35788 37280 35816
rect 35805 35779 35863 35785
rect 37274 35776 37280 35788
rect 37332 35776 37338 35828
rect 27430 35708 27436 35760
rect 27488 35748 27494 35760
rect 29917 35751 29975 35757
rect 27488 35720 28396 35748
rect 27488 35708 27494 35720
rect 1719 35652 2728 35680
rect 2869 35683 2927 35689
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 2869 35649 2881 35683
rect 2915 35680 2927 35683
rect 3142 35680 3148 35692
rect 2915 35652 3148 35680
rect 2915 35649 2927 35652
rect 2869 35643 2927 35649
rect 2225 35615 2283 35621
rect 2225 35581 2237 35615
rect 2271 35612 2283 35615
rect 2884 35612 2912 35643
rect 3142 35640 3148 35652
rect 3200 35640 3206 35692
rect 3513 35683 3571 35689
rect 3513 35649 3525 35683
rect 3559 35680 3571 35683
rect 3694 35680 3700 35692
rect 3559 35652 3700 35680
rect 3559 35649 3571 35652
rect 3513 35643 3571 35649
rect 3694 35640 3700 35652
rect 3752 35640 3758 35692
rect 6457 35683 6515 35689
rect 6457 35649 6469 35683
rect 6503 35680 6515 35683
rect 8757 35683 8815 35689
rect 6503 35652 6914 35680
rect 6503 35649 6515 35652
rect 6457 35643 6515 35649
rect 2271 35584 2912 35612
rect 2271 35581 2283 35584
rect 2225 35575 2283 35581
rect 6886 35544 6914 35652
rect 8757 35649 8769 35683
rect 8803 35680 8815 35683
rect 8846 35680 8852 35692
rect 8803 35652 8852 35680
rect 8803 35649 8815 35652
rect 8757 35643 8815 35649
rect 8846 35640 8852 35652
rect 8904 35640 8910 35692
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35649 10011 35683
rect 9953 35643 10011 35649
rect 10965 35683 11023 35689
rect 10965 35649 10977 35683
rect 11011 35680 11023 35683
rect 11054 35680 11060 35692
rect 11011 35652 11060 35680
rect 11011 35649 11023 35652
rect 10965 35643 11023 35649
rect 9968 35612 9996 35643
rect 11054 35640 11060 35652
rect 11112 35640 11118 35692
rect 11517 35683 11575 35689
rect 11517 35649 11529 35683
rect 11563 35680 11575 35683
rect 11698 35680 11704 35692
rect 11563 35652 11704 35680
rect 11563 35649 11575 35652
rect 11517 35643 11575 35649
rect 11698 35640 11704 35652
rect 11756 35640 11762 35692
rect 12437 35683 12495 35689
rect 12437 35649 12449 35683
rect 12483 35680 12495 35683
rect 12618 35680 12624 35692
rect 12483 35652 12624 35680
rect 12483 35649 12495 35652
rect 12437 35643 12495 35649
rect 12618 35640 12624 35652
rect 12676 35640 12682 35692
rect 14182 35640 14188 35692
rect 14240 35680 14246 35692
rect 14369 35683 14427 35689
rect 14369 35680 14381 35683
rect 14240 35652 14381 35680
rect 14240 35640 14246 35652
rect 14369 35649 14381 35652
rect 14415 35649 14427 35683
rect 14369 35643 14427 35649
rect 14734 35640 14740 35692
rect 14792 35680 14798 35692
rect 15013 35683 15071 35689
rect 15013 35680 15025 35683
rect 14792 35652 15025 35680
rect 14792 35640 14798 35652
rect 15013 35649 15025 35652
rect 15059 35649 15071 35683
rect 15013 35643 15071 35649
rect 15841 35683 15899 35689
rect 15841 35649 15853 35683
rect 15887 35680 15899 35683
rect 15930 35680 15936 35692
rect 15887 35652 15936 35680
rect 15887 35649 15899 35652
rect 15841 35643 15899 35649
rect 15930 35640 15936 35652
rect 15988 35640 15994 35692
rect 16758 35640 16764 35692
rect 16816 35680 16822 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16816 35652 16865 35680
rect 16816 35640 16822 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 17497 35683 17555 35689
rect 17497 35649 17509 35683
rect 17543 35680 17555 35683
rect 17862 35680 17868 35692
rect 17543 35652 17868 35680
rect 17543 35649 17555 35652
rect 17497 35643 17555 35649
rect 17862 35640 17868 35652
rect 17920 35640 17926 35692
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 19521 35643 19579 35649
rect 11238 35612 11244 35624
rect 9968 35584 11244 35612
rect 11238 35572 11244 35584
rect 11296 35572 11302 35624
rect 16666 35572 16672 35624
rect 16724 35612 16730 35624
rect 18969 35615 19027 35621
rect 18969 35612 18981 35615
rect 16724 35584 18981 35612
rect 16724 35572 16730 35584
rect 18969 35581 18981 35584
rect 19015 35612 19027 35615
rect 19536 35612 19564 35643
rect 22830 35640 22836 35692
rect 22888 35680 22894 35692
rect 23017 35683 23075 35689
rect 23017 35680 23029 35683
rect 22888 35652 23029 35680
rect 22888 35640 22894 35652
rect 23017 35649 23029 35652
rect 23063 35649 23075 35683
rect 23017 35643 23075 35649
rect 26142 35640 26148 35692
rect 26200 35680 26206 35692
rect 26237 35683 26295 35689
rect 26237 35680 26249 35683
rect 26200 35652 26249 35680
rect 26200 35640 26206 35652
rect 26237 35649 26249 35652
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 26878 35640 26884 35692
rect 26936 35680 26942 35692
rect 26973 35683 27031 35689
rect 26973 35680 26985 35683
rect 26936 35652 26985 35680
rect 26936 35640 26942 35652
rect 26973 35649 26985 35652
rect 27019 35649 27031 35683
rect 26973 35643 27031 35649
rect 27154 35640 27160 35692
rect 27212 35680 27218 35692
rect 28368 35689 28396 35720
rect 29917 35717 29929 35751
rect 29963 35748 29975 35751
rect 30558 35748 30564 35760
rect 29963 35720 30564 35748
rect 29963 35717 29975 35720
rect 29917 35711 29975 35717
rect 30558 35708 30564 35720
rect 30616 35708 30622 35760
rect 27525 35683 27583 35689
rect 27525 35680 27537 35683
rect 27212 35652 27537 35680
rect 27212 35640 27218 35652
rect 27525 35649 27537 35652
rect 27571 35649 27583 35683
rect 27525 35643 27583 35649
rect 28353 35683 28411 35689
rect 28353 35649 28365 35683
rect 28399 35680 28411 35683
rect 28813 35683 28871 35689
rect 28813 35680 28825 35683
rect 28399 35652 28825 35680
rect 28399 35649 28411 35652
rect 28353 35643 28411 35649
rect 28813 35649 28825 35652
rect 28859 35649 28871 35683
rect 28813 35643 28871 35649
rect 30653 35683 30711 35689
rect 30653 35649 30665 35683
rect 30699 35680 30711 35683
rect 31294 35680 31300 35692
rect 30699 35652 31300 35680
rect 30699 35649 30711 35652
rect 30653 35643 30711 35649
rect 31294 35640 31300 35652
rect 31352 35640 31358 35692
rect 32766 35680 32772 35692
rect 32727 35652 32772 35680
rect 32766 35640 32772 35652
rect 32824 35640 32830 35692
rect 33597 35683 33655 35689
rect 33597 35649 33609 35683
rect 33643 35680 33655 35683
rect 33962 35680 33968 35692
rect 33643 35652 33968 35680
rect 33643 35649 33655 35652
rect 33597 35643 33655 35649
rect 33962 35640 33968 35652
rect 34020 35640 34026 35692
rect 34054 35640 34060 35692
rect 34112 35680 34118 35692
rect 35161 35683 35219 35689
rect 34112 35652 34157 35680
rect 34112 35640 34118 35652
rect 35161 35649 35173 35683
rect 35207 35649 35219 35683
rect 35161 35643 35219 35649
rect 19015 35584 19564 35612
rect 19015 35581 19027 35584
rect 18969 35575 19027 35581
rect 7193 35547 7251 35553
rect 7193 35544 7205 35547
rect 6886 35516 7205 35544
rect 7193 35513 7205 35516
rect 7239 35544 7251 35547
rect 8110 35544 8116 35556
rect 7239 35516 8116 35544
rect 7239 35513 7251 35516
rect 7193 35507 7251 35513
rect 8110 35504 8116 35516
rect 8168 35504 8174 35556
rect 11701 35547 11759 35553
rect 11701 35513 11713 35547
rect 11747 35544 11759 35547
rect 22554 35544 22560 35556
rect 11747 35516 22560 35544
rect 11747 35513 11759 35516
rect 11701 35507 11759 35513
rect 22554 35504 22560 35516
rect 22612 35504 22618 35556
rect 24946 35504 24952 35556
rect 25004 35544 25010 35556
rect 26896 35544 26924 35640
rect 35176 35612 35204 35643
rect 35434 35640 35440 35692
rect 35492 35680 35498 35692
rect 35621 35683 35679 35689
rect 35621 35680 35633 35683
rect 35492 35652 35633 35680
rect 35492 35640 35498 35652
rect 35621 35649 35633 35652
rect 35667 35649 35679 35683
rect 35621 35643 35679 35649
rect 36354 35640 36360 35692
rect 36412 35680 36418 35692
rect 36449 35683 36507 35689
rect 36449 35680 36461 35683
rect 36412 35652 36461 35680
rect 36412 35640 36418 35652
rect 36449 35649 36461 35652
rect 36495 35649 36507 35683
rect 36449 35643 36507 35649
rect 37826 35640 37832 35692
rect 37884 35680 37890 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37884 35652 38025 35680
rect 37884 35640 37890 35652
rect 38013 35649 38025 35652
rect 38059 35680 38071 35683
rect 39022 35680 39028 35692
rect 38059 35652 39028 35680
rect 38059 35649 38071 35652
rect 38013 35643 38071 35649
rect 39022 35640 39028 35652
rect 39080 35640 39086 35692
rect 35526 35612 35532 35624
rect 35176 35584 35532 35612
rect 35526 35572 35532 35584
rect 35584 35572 35590 35624
rect 25004 35516 26924 35544
rect 27709 35547 27767 35553
rect 25004 35504 25010 35516
rect 27709 35513 27721 35547
rect 27755 35544 27767 35547
rect 29454 35544 29460 35556
rect 27755 35516 29460 35544
rect 27755 35513 27767 35516
rect 27709 35507 27767 35513
rect 29454 35504 29460 35516
rect 29512 35504 29518 35556
rect 33410 35504 33416 35556
rect 33468 35544 33474 35556
rect 34241 35547 34299 35553
rect 34241 35544 34253 35547
rect 33468 35516 34253 35544
rect 33468 35504 33474 35516
rect 34241 35513 34253 35516
rect 34287 35513 34299 35547
rect 34241 35507 34299 35513
rect 34977 35547 35035 35553
rect 34977 35513 34989 35547
rect 35023 35544 35035 35547
rect 36538 35544 36544 35556
rect 35023 35516 36544 35544
rect 35023 35513 35035 35516
rect 34977 35507 35035 35513
rect 36538 35504 36544 35516
rect 36596 35504 36602 35556
rect 36633 35547 36691 35553
rect 36633 35513 36645 35547
rect 36679 35544 36691 35547
rect 37366 35544 37372 35556
rect 36679 35516 37372 35544
rect 36679 35513 36691 35516
rect 36633 35507 36691 35513
rect 37366 35504 37372 35516
rect 37424 35504 37430 35556
rect 3694 35436 3700 35488
rect 3752 35476 3758 35488
rect 3973 35479 4031 35485
rect 3973 35476 3985 35479
rect 3752 35448 3985 35476
rect 3752 35436 3758 35448
rect 3973 35445 3985 35448
rect 4019 35445 4031 35479
rect 5718 35476 5724 35488
rect 5679 35448 5724 35476
rect 3973 35439 4031 35445
rect 5718 35436 5724 35448
rect 5776 35436 5782 35488
rect 8018 35476 8024 35488
rect 7979 35448 8024 35476
rect 8018 35436 8024 35448
rect 8076 35436 8082 35488
rect 12618 35436 12624 35488
rect 12676 35476 12682 35488
rect 12897 35479 12955 35485
rect 12897 35476 12909 35479
rect 12676 35448 12909 35476
rect 12676 35436 12682 35448
rect 12897 35445 12909 35448
rect 12943 35445 12955 35479
rect 13446 35476 13452 35488
rect 13407 35448 13452 35476
rect 12897 35439 12955 35445
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 17862 35436 17868 35488
rect 17920 35476 17926 35488
rect 17957 35479 18015 35485
rect 17957 35476 17969 35479
rect 17920 35448 17969 35476
rect 17920 35436 17926 35448
rect 17957 35445 17969 35448
rect 18003 35445 18015 35479
rect 17957 35439 18015 35445
rect 19978 35436 19984 35488
rect 20036 35476 20042 35488
rect 20165 35479 20223 35485
rect 20165 35476 20177 35479
rect 20036 35448 20177 35476
rect 20036 35436 20042 35448
rect 20165 35445 20177 35448
rect 20211 35445 20223 35479
rect 20714 35476 20720 35488
rect 20675 35448 20720 35476
rect 20165 35439 20223 35445
rect 20714 35436 20720 35448
rect 20772 35436 20778 35488
rect 21910 35476 21916 35488
rect 21871 35448 21916 35476
rect 21910 35436 21916 35448
rect 21968 35436 21974 35488
rect 24854 35476 24860 35488
rect 24815 35448 24860 35476
rect 24854 35436 24860 35448
rect 24912 35436 24918 35488
rect 25406 35476 25412 35488
rect 25367 35448 25412 35476
rect 25406 35436 25412 35448
rect 25464 35436 25470 35488
rect 28166 35476 28172 35488
rect 28127 35448 28172 35476
rect 28166 35436 28172 35448
rect 28224 35436 28230 35488
rect 29638 35436 29644 35488
rect 29696 35476 29702 35488
rect 32677 35479 32735 35485
rect 32677 35476 32689 35479
rect 29696 35448 32689 35476
rect 29696 35436 29702 35448
rect 32677 35445 32689 35448
rect 32723 35445 32735 35479
rect 32677 35439 32735 35445
rect 37921 35479 37979 35485
rect 37921 35445 37933 35479
rect 37967 35476 37979 35479
rect 38746 35476 38752 35488
rect 37967 35448 38752 35476
rect 37967 35445 37979 35448
rect 37921 35439 37979 35445
rect 38746 35436 38752 35448
rect 38804 35436 38810 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1578 35272 1584 35284
rect 1539 35244 1584 35272
rect 1578 35232 1584 35244
rect 1636 35232 1642 35284
rect 1762 35232 1768 35284
rect 1820 35272 1826 35284
rect 2133 35275 2191 35281
rect 2133 35272 2145 35275
rect 1820 35244 2145 35272
rect 1820 35232 1826 35244
rect 2133 35241 2145 35244
rect 2179 35241 2191 35275
rect 6178 35272 6184 35284
rect 6139 35244 6184 35272
rect 2133 35235 2191 35241
rect 6178 35232 6184 35244
rect 6236 35232 6242 35284
rect 6730 35272 6736 35284
rect 6691 35244 6736 35272
rect 6730 35232 6736 35244
rect 6788 35232 6794 35284
rect 7466 35232 7472 35284
rect 7524 35272 7530 35284
rect 7837 35275 7895 35281
rect 7837 35272 7849 35275
rect 7524 35244 7849 35272
rect 7524 35232 7530 35244
rect 7837 35241 7849 35244
rect 7883 35241 7895 35275
rect 7837 35235 7895 35241
rect 9582 35232 9588 35284
rect 9640 35272 9646 35284
rect 9953 35275 10011 35281
rect 9953 35272 9965 35275
rect 9640 35244 9965 35272
rect 9640 35232 9646 35244
rect 9953 35241 9965 35244
rect 9999 35272 10011 35275
rect 10134 35272 10140 35284
rect 9999 35244 10140 35272
rect 9999 35241 10011 35244
rect 9953 35235 10011 35241
rect 10134 35232 10140 35244
rect 10192 35232 10198 35284
rect 10226 35232 10232 35284
rect 10284 35272 10290 35284
rect 10413 35275 10471 35281
rect 10413 35272 10425 35275
rect 10284 35244 10425 35272
rect 10284 35232 10290 35244
rect 10413 35241 10425 35244
rect 10459 35241 10471 35275
rect 12158 35272 12164 35284
rect 12119 35244 12164 35272
rect 10413 35235 10471 35241
rect 12158 35232 12164 35244
rect 12216 35232 12222 35284
rect 12710 35272 12716 35284
rect 12671 35244 12716 35272
rect 12710 35232 12716 35244
rect 12768 35232 12774 35284
rect 15289 35275 15347 35281
rect 15289 35241 15301 35275
rect 15335 35272 15347 35275
rect 15378 35272 15384 35284
rect 15335 35244 15384 35272
rect 15335 35241 15347 35244
rect 15289 35235 15347 35241
rect 15378 35232 15384 35244
rect 15436 35232 15442 35284
rect 17494 35272 17500 35284
rect 17455 35244 17500 35272
rect 17494 35232 17500 35244
rect 17552 35232 17558 35284
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18049 35275 18107 35281
rect 18049 35272 18061 35275
rect 18012 35244 18061 35272
rect 18012 35232 18018 35244
rect 18049 35241 18061 35244
rect 18095 35241 18107 35275
rect 18598 35272 18604 35284
rect 18559 35244 18604 35272
rect 18049 35235 18107 35241
rect 18598 35232 18604 35244
rect 18656 35232 18662 35284
rect 19242 35272 19248 35284
rect 19203 35244 19248 35272
rect 19242 35232 19248 35244
rect 19300 35232 19306 35284
rect 20070 35272 20076 35284
rect 20031 35244 20076 35272
rect 20070 35232 20076 35244
rect 20128 35232 20134 35284
rect 29546 35272 29552 35284
rect 29507 35244 29552 35272
rect 29546 35232 29552 35244
rect 29604 35232 29610 35284
rect 33502 35272 33508 35284
rect 33463 35244 33508 35272
rect 33502 35232 33508 35244
rect 33560 35232 33566 35284
rect 35345 35275 35403 35281
rect 35345 35241 35357 35275
rect 35391 35272 35403 35275
rect 35618 35272 35624 35284
rect 35391 35244 35624 35272
rect 35391 35241 35403 35244
rect 35345 35235 35403 35241
rect 35618 35232 35624 35244
rect 35676 35232 35682 35284
rect 38013 35275 38071 35281
rect 38013 35241 38025 35275
rect 38059 35272 38071 35275
rect 38286 35272 38292 35284
rect 38059 35244 38292 35272
rect 38059 35241 38071 35244
rect 38013 35235 38071 35241
rect 38286 35232 38292 35244
rect 38344 35232 38350 35284
rect 1670 35164 1676 35216
rect 1728 35204 1734 35216
rect 2685 35207 2743 35213
rect 2685 35204 2697 35207
rect 1728 35176 2697 35204
rect 1728 35164 1734 35176
rect 2685 35173 2697 35176
rect 2731 35173 2743 35207
rect 2685 35167 2743 35173
rect 15933 35207 15991 35213
rect 15933 35173 15945 35207
rect 15979 35204 15991 35207
rect 26329 35207 26387 35213
rect 15979 35176 16574 35204
rect 15979 35173 15991 35176
rect 15933 35167 15991 35173
rect 16546 35136 16574 35176
rect 26329 35173 26341 35207
rect 26375 35204 26387 35207
rect 28166 35204 28172 35216
rect 26375 35176 28172 35204
rect 26375 35173 26387 35176
rect 26329 35167 26387 35173
rect 28166 35164 28172 35176
rect 28224 35164 28230 35216
rect 25498 35136 25504 35148
rect 16546 35108 25504 35136
rect 25498 35096 25504 35108
rect 25556 35096 25562 35148
rect 28442 35096 28448 35148
rect 28500 35136 28506 35148
rect 30101 35139 30159 35145
rect 30101 35136 30113 35139
rect 28500 35108 30113 35136
rect 28500 35096 28506 35108
rect 30101 35105 30113 35108
rect 30147 35105 30159 35139
rect 30101 35099 30159 35105
rect 32968 35108 36124 35136
rect 2869 35071 2927 35077
rect 2869 35037 2881 35071
rect 2915 35068 2927 35071
rect 10594 35068 10600 35080
rect 2915 35040 3924 35068
rect 10555 35040 10600 35068
rect 2915 35037 2927 35040
rect 2869 35031 2927 35037
rect 3896 34944 3924 35040
rect 10594 35028 10600 35040
rect 10652 35028 10658 35080
rect 15102 35068 15108 35080
rect 15063 35040 15108 35068
rect 15102 35028 15108 35040
rect 15160 35028 15166 35080
rect 15746 35068 15752 35080
rect 15707 35040 15752 35068
rect 15746 35028 15752 35040
rect 15804 35068 15810 35080
rect 16393 35071 16451 35077
rect 16393 35068 16405 35071
rect 15804 35040 16405 35068
rect 15804 35028 15810 35040
rect 16393 35037 16405 35040
rect 16439 35037 16451 35071
rect 29638 35068 29644 35080
rect 16393 35031 16451 35037
rect 16546 35040 29644 35068
rect 13354 35000 13360 35012
rect 13267 34972 13360 35000
rect 13354 34960 13360 34972
rect 13412 35000 13418 35012
rect 16546 35000 16574 35040
rect 29638 35028 29644 35040
rect 29696 35028 29702 35080
rect 30009 35071 30067 35077
rect 30009 35037 30021 35071
rect 30055 35068 30067 35071
rect 32968 35068 32996 35108
rect 36096 35080 36124 35108
rect 30055 35040 32996 35068
rect 35529 35071 35587 35077
rect 30055 35037 30067 35040
rect 30009 35031 30067 35037
rect 35529 35037 35541 35071
rect 35575 35068 35587 35071
rect 35986 35068 35992 35080
rect 35575 35040 35894 35068
rect 35947 35040 35992 35068
rect 35575 35037 35587 35040
rect 35529 35031 35587 35037
rect 13412 34972 16574 35000
rect 13412 34960 13418 34972
rect 20438 34960 20444 35012
rect 20496 35000 20502 35012
rect 25961 35003 26019 35009
rect 20496 34972 21128 35000
rect 20496 34960 20502 34972
rect 21100 34944 21128 34972
rect 25961 34969 25973 35003
rect 26007 35000 26019 35003
rect 26234 35000 26240 35012
rect 26007 34972 26240 35000
rect 26007 34969 26019 34972
rect 25961 34963 26019 34969
rect 26234 34960 26240 34972
rect 26292 34960 26298 35012
rect 30558 34960 30564 35012
rect 30616 35000 30622 35012
rect 31389 35003 31447 35009
rect 31389 35000 31401 35003
rect 30616 34972 31401 35000
rect 30616 34960 30622 34972
rect 31389 34969 31401 34972
rect 31435 35000 31447 35003
rect 31662 35000 31668 35012
rect 31435 34972 31668 35000
rect 31435 34969 31447 34972
rect 31389 34963 31447 34969
rect 31662 34960 31668 34972
rect 31720 34960 31726 35012
rect 3878 34932 3884 34944
rect 3839 34904 3884 34932
rect 3878 34892 3884 34904
rect 3936 34892 3942 34944
rect 4433 34935 4491 34941
rect 4433 34901 4445 34935
rect 4479 34932 4491 34935
rect 4706 34932 4712 34944
rect 4479 34904 4712 34932
rect 4479 34901 4491 34904
rect 4433 34895 4491 34901
rect 4706 34892 4712 34904
rect 4764 34892 4770 34944
rect 4985 34935 5043 34941
rect 4985 34901 4997 34935
rect 5031 34932 5043 34935
rect 5074 34932 5080 34944
rect 5031 34904 5080 34932
rect 5031 34901 5043 34904
rect 4985 34895 5043 34901
rect 5074 34892 5080 34904
rect 5132 34892 5138 34944
rect 5534 34932 5540 34944
rect 5495 34904 5540 34932
rect 5534 34892 5540 34904
rect 5592 34892 5598 34944
rect 7098 34892 7104 34944
rect 7156 34932 7162 34944
rect 7285 34935 7343 34941
rect 7285 34932 7297 34935
rect 7156 34904 7297 34932
rect 7156 34892 7162 34904
rect 7285 34901 7297 34904
rect 7331 34901 7343 34935
rect 7285 34895 7343 34901
rect 8846 34892 8852 34944
rect 8904 34932 8910 34944
rect 8941 34935 8999 34941
rect 8941 34932 8953 34935
rect 8904 34904 8953 34932
rect 8904 34892 8910 34904
rect 8941 34901 8953 34904
rect 8987 34901 8999 34935
rect 11054 34932 11060 34944
rect 11015 34904 11060 34932
rect 8941 34895 8999 34901
rect 11054 34892 11060 34904
rect 11112 34892 11118 34944
rect 11698 34932 11704 34944
rect 11659 34904 11704 34932
rect 11698 34892 11704 34904
rect 11756 34892 11762 34944
rect 14182 34892 14188 34944
rect 14240 34932 14246 34944
rect 14461 34935 14519 34941
rect 14461 34932 14473 34935
rect 14240 34904 14473 34932
rect 14240 34892 14246 34904
rect 14461 34901 14473 34904
rect 14507 34901 14519 34935
rect 14461 34895 14519 34901
rect 16758 34892 16764 34944
rect 16816 34932 16822 34944
rect 16945 34935 17003 34941
rect 16945 34932 16957 34935
rect 16816 34904 16957 34932
rect 16816 34892 16822 34904
rect 16945 34901 16957 34904
rect 16991 34901 17003 34935
rect 16945 34895 17003 34901
rect 19426 34892 19432 34944
rect 19484 34932 19490 34944
rect 20530 34932 20536 34944
rect 19484 34904 20536 34932
rect 19484 34892 19490 34904
rect 20530 34892 20536 34904
rect 20588 34892 20594 34944
rect 21082 34932 21088 34944
rect 21043 34904 21088 34932
rect 21082 34892 21088 34904
rect 21140 34892 21146 34944
rect 22186 34892 22192 34944
rect 22244 34932 22250 34944
rect 22830 34932 22836 34944
rect 22244 34904 22836 34932
rect 22244 34892 22250 34904
rect 22830 34892 22836 34904
rect 22888 34892 22894 34944
rect 26326 34892 26332 34944
rect 26384 34932 26390 34944
rect 26421 34935 26479 34941
rect 26421 34932 26433 34935
rect 26384 34904 26433 34932
rect 26384 34892 26390 34904
rect 26421 34901 26433 34904
rect 26467 34901 26479 34935
rect 26421 34895 26479 34901
rect 28997 34935 29055 34941
rect 28997 34901 29009 34935
rect 29043 34932 29055 34935
rect 29914 34932 29920 34944
rect 29043 34904 29920 34932
rect 29043 34901 29055 34904
rect 28997 34895 29055 34901
rect 29914 34892 29920 34904
rect 29972 34892 29978 34944
rect 30374 34892 30380 34944
rect 30432 34932 30438 34944
rect 30837 34935 30895 34941
rect 30837 34932 30849 34935
rect 30432 34904 30849 34932
rect 30432 34892 30438 34904
rect 30837 34901 30849 34904
rect 30883 34932 30895 34935
rect 31018 34932 31024 34944
rect 30883 34904 31024 34932
rect 30883 34901 30895 34904
rect 30837 34895 30895 34901
rect 31018 34892 31024 34904
rect 31076 34892 31082 34944
rect 31938 34932 31944 34944
rect 31899 34904 31944 34932
rect 31938 34892 31944 34904
rect 31996 34892 32002 34944
rect 32766 34892 32772 34944
rect 32824 34932 32830 34944
rect 32953 34935 33011 34941
rect 32953 34932 32965 34935
rect 32824 34904 32965 34932
rect 32824 34892 32830 34904
rect 32953 34901 32965 34904
rect 32999 34901 33011 34935
rect 32953 34895 33011 34901
rect 33226 34892 33232 34944
rect 33284 34932 33290 34944
rect 34057 34935 34115 34941
rect 34057 34932 34069 34935
rect 33284 34904 34069 34932
rect 33284 34892 33290 34904
rect 34057 34901 34069 34904
rect 34103 34932 34115 34935
rect 34238 34932 34244 34944
rect 34103 34904 34244 34932
rect 34103 34901 34115 34904
rect 34057 34895 34115 34901
rect 34238 34892 34244 34904
rect 34296 34892 34302 34944
rect 34698 34932 34704 34944
rect 34659 34904 34704 34932
rect 34698 34892 34704 34904
rect 34756 34892 34762 34944
rect 35866 34932 35894 35040
rect 35986 35028 35992 35040
rect 36044 35028 36050 35080
rect 36078 35028 36084 35080
rect 36136 35028 36142 35080
rect 37274 35028 37280 35080
rect 37332 35068 37338 35080
rect 37829 35071 37887 35077
rect 37829 35068 37841 35071
rect 37332 35040 37841 35068
rect 37332 35028 37338 35040
rect 37829 35037 37841 35040
rect 37875 35068 37887 35071
rect 38286 35068 38292 35080
rect 37875 35040 38292 35068
rect 37875 35037 37887 35040
rect 37829 35031 37887 35037
rect 38286 35028 38292 35040
rect 38344 35028 38350 35080
rect 36256 35003 36314 35009
rect 36256 34969 36268 35003
rect 36302 35000 36314 35003
rect 36446 35000 36452 35012
rect 36302 34972 36452 35000
rect 36302 34969 36314 34972
rect 36256 34963 36314 34969
rect 36446 34960 36452 34972
rect 36504 34960 36510 35012
rect 37369 34935 37427 34941
rect 37369 34932 37381 34935
rect 35866 34904 37381 34932
rect 37369 34901 37381 34904
rect 37415 34901 37427 34935
rect 37369 34895 37427 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2590 34728 2596 34740
rect 2551 34700 2596 34728
rect 2590 34688 2596 34700
rect 2648 34688 2654 34740
rect 9214 34728 9220 34740
rect 9175 34700 9220 34728
rect 9214 34688 9220 34700
rect 9272 34688 9278 34740
rect 12161 34731 12219 34737
rect 12161 34697 12173 34731
rect 12207 34728 12219 34731
rect 12250 34728 12256 34740
rect 12207 34700 12256 34728
rect 12207 34697 12219 34700
rect 12161 34691 12219 34697
rect 12250 34688 12256 34700
rect 12308 34688 12314 34740
rect 12894 34728 12900 34740
rect 12855 34700 12900 34728
rect 12894 34688 12900 34700
rect 12952 34688 12958 34740
rect 15102 34688 15108 34740
rect 15160 34728 15166 34740
rect 15657 34731 15715 34737
rect 15657 34728 15669 34731
rect 15160 34700 15669 34728
rect 15160 34688 15166 34700
rect 15657 34697 15669 34700
rect 15703 34697 15715 34731
rect 16942 34728 16948 34740
rect 16903 34700 16948 34728
rect 15657 34691 15715 34697
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 20254 34688 20260 34740
rect 20312 34728 20318 34740
rect 23293 34731 23351 34737
rect 20312 34700 20576 34728
rect 20312 34688 20318 34700
rect 3050 34620 3056 34672
rect 3108 34660 3114 34672
rect 3605 34663 3663 34669
rect 3605 34660 3617 34663
rect 3108 34632 3617 34660
rect 3108 34620 3114 34632
rect 3605 34629 3617 34632
rect 3651 34629 3663 34663
rect 6365 34663 6423 34669
rect 6365 34660 6377 34663
rect 3605 34623 3663 34629
rect 4448 34632 6377 34660
rect 2866 34484 2872 34536
rect 2924 34524 2930 34536
rect 3053 34527 3111 34533
rect 3053 34524 3065 34527
rect 2924 34496 3065 34524
rect 2924 34484 2930 34496
rect 3053 34493 3065 34496
rect 3099 34524 3111 34527
rect 3234 34524 3240 34536
rect 3099 34496 3240 34524
rect 3099 34493 3111 34496
rect 3053 34487 3111 34493
rect 3234 34484 3240 34496
rect 3292 34484 3298 34536
rect 4154 34484 4160 34536
rect 4212 34524 4218 34536
rect 4448 34533 4476 34632
rect 6365 34629 6377 34632
rect 6411 34660 6423 34663
rect 9490 34660 9496 34672
rect 6411 34632 9496 34660
rect 6411 34629 6423 34632
rect 6365 34623 6423 34629
rect 9490 34620 9496 34632
rect 9548 34620 9554 34672
rect 19058 34620 19064 34672
rect 19116 34660 19122 34672
rect 19978 34660 19984 34672
rect 19116 34632 19984 34660
rect 19116 34620 19122 34632
rect 19978 34620 19984 34632
rect 20036 34620 20042 34672
rect 4700 34595 4758 34601
rect 4700 34561 4712 34595
rect 4746 34592 4758 34595
rect 5258 34592 5264 34604
rect 4746 34564 5264 34592
rect 4746 34561 4758 34564
rect 4700 34555 4758 34561
rect 5258 34552 5264 34564
rect 5316 34552 5322 34604
rect 13906 34592 13912 34604
rect 13867 34564 13912 34592
rect 13906 34552 13912 34564
rect 13964 34552 13970 34604
rect 14274 34552 14280 34604
rect 14332 34592 14338 34604
rect 14550 34592 14556 34604
rect 14332 34564 14556 34592
rect 14332 34552 14338 34564
rect 14550 34552 14556 34564
rect 14608 34552 14614 34604
rect 14734 34552 14740 34604
rect 14792 34592 14798 34604
rect 18322 34601 18328 34604
rect 15105 34595 15163 34601
rect 15105 34592 15117 34595
rect 14792 34564 15117 34592
rect 14792 34552 14798 34564
rect 15105 34561 15117 34564
rect 15151 34561 15163 34595
rect 15105 34555 15163 34561
rect 18316 34555 18328 34601
rect 18380 34592 18386 34604
rect 18380 34564 18416 34592
rect 18322 34552 18328 34555
rect 18380 34552 18386 34564
rect 4433 34527 4491 34533
rect 4433 34524 4445 34527
rect 4212 34496 4445 34524
rect 4212 34484 4218 34496
rect 4433 34493 4445 34496
rect 4479 34493 4491 34527
rect 9766 34524 9772 34536
rect 9727 34496 9772 34524
rect 4433 34487 4491 34493
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 10594 34484 10600 34536
rect 10652 34524 10658 34536
rect 10689 34527 10747 34533
rect 10689 34524 10701 34527
rect 10652 34496 10701 34524
rect 10652 34484 10658 34496
rect 10689 34493 10701 34496
rect 10735 34493 10747 34527
rect 10689 34487 10747 34493
rect 11238 34484 11244 34536
rect 11296 34524 11302 34536
rect 11517 34527 11575 34533
rect 11517 34524 11529 34527
rect 11296 34496 11529 34524
rect 11296 34484 11302 34496
rect 11517 34493 11529 34496
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 13722 34484 13728 34536
rect 13780 34524 13786 34536
rect 17497 34527 17555 34533
rect 17497 34524 17509 34527
rect 13780 34496 17509 34524
rect 13780 34484 13786 34496
rect 17497 34493 17509 34496
rect 17543 34524 17555 34527
rect 18049 34527 18107 34533
rect 18049 34524 18061 34527
rect 17543 34496 18061 34524
rect 17543 34493 17555 34496
rect 17497 34487 17555 34493
rect 18049 34493 18061 34496
rect 18095 34493 18107 34527
rect 18049 34487 18107 34493
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20254 34524 20260 34536
rect 20027 34496 20260 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 20254 34484 20260 34496
rect 20312 34484 20318 34536
rect 20548 34533 20576 34700
rect 23293 34697 23305 34731
rect 23339 34728 23351 34731
rect 23842 34728 23848 34740
rect 23339 34700 23848 34728
rect 23339 34697 23351 34700
rect 23293 34691 23351 34697
rect 23842 34688 23848 34700
rect 23900 34688 23906 34740
rect 24213 34731 24271 34737
rect 24213 34697 24225 34731
rect 24259 34728 24271 34731
rect 27154 34728 27160 34740
rect 24259 34700 27160 34728
rect 24259 34697 24271 34700
rect 24213 34691 24271 34697
rect 27154 34688 27160 34700
rect 27212 34688 27218 34740
rect 35802 34688 35808 34740
rect 35860 34728 35866 34740
rect 36541 34731 36599 34737
rect 36541 34728 36553 34731
rect 35860 34700 36553 34728
rect 35860 34688 35866 34700
rect 36541 34697 36553 34700
rect 36587 34697 36599 34731
rect 37274 34728 37280 34740
rect 36541 34691 36599 34697
rect 37108 34700 37280 34728
rect 22833 34663 22891 34669
rect 22833 34629 22845 34663
rect 22879 34660 22891 34663
rect 23106 34660 23112 34672
rect 22879 34632 23112 34660
rect 22879 34629 22891 34632
rect 22833 34623 22891 34629
rect 23106 34620 23112 34632
rect 23164 34660 23170 34672
rect 23753 34663 23811 34669
rect 23753 34660 23765 34663
rect 23164 34632 23765 34660
rect 23164 34620 23170 34632
rect 23753 34629 23765 34632
rect 23799 34660 23811 34663
rect 26234 34660 26240 34672
rect 23799 34632 26240 34660
rect 23799 34629 23811 34632
rect 23753 34623 23811 34629
rect 26234 34620 26240 34632
rect 26292 34660 26298 34672
rect 27522 34660 27528 34672
rect 26292 34632 27528 34660
rect 26292 34620 26298 34632
rect 27522 34620 27528 34632
rect 27580 34620 27586 34672
rect 34793 34663 34851 34669
rect 34793 34629 34805 34663
rect 34839 34660 34851 34663
rect 37108 34660 37136 34700
rect 37274 34688 37280 34700
rect 37332 34688 37338 34740
rect 37369 34731 37427 34737
rect 37369 34697 37381 34731
rect 37415 34728 37427 34731
rect 37918 34728 37924 34740
rect 37415 34700 37924 34728
rect 37415 34697 37427 34700
rect 37369 34691 37427 34697
rect 37918 34688 37924 34700
rect 37976 34688 37982 34740
rect 38013 34731 38071 34737
rect 38013 34697 38025 34731
rect 38059 34728 38071 34731
rect 39390 34728 39396 34740
rect 38059 34700 39396 34728
rect 38059 34697 38071 34700
rect 38013 34691 38071 34697
rect 39390 34688 39396 34700
rect 39448 34688 39454 34740
rect 34839 34632 37136 34660
rect 34839 34629 34851 34632
rect 34793 34623 34851 34629
rect 37182 34620 37188 34672
rect 37240 34660 37246 34672
rect 39758 34660 39764 34672
rect 37240 34632 39764 34660
rect 37240 34620 37246 34632
rect 39758 34620 39764 34632
rect 39816 34620 39822 34672
rect 35250 34592 35256 34604
rect 35211 34564 35256 34592
rect 35250 34552 35256 34564
rect 35308 34592 35314 34604
rect 36170 34592 36176 34604
rect 35308 34564 36176 34592
rect 35308 34552 35314 34564
rect 36170 34552 36176 34564
rect 36228 34552 36234 34604
rect 36725 34595 36783 34601
rect 36725 34561 36737 34595
rect 36771 34592 36783 34595
rect 37550 34592 37556 34604
rect 36771 34564 37556 34592
rect 36771 34561 36783 34564
rect 36725 34555 36783 34561
rect 37550 34552 37556 34564
rect 37608 34552 37614 34604
rect 37829 34595 37887 34601
rect 37829 34561 37841 34595
rect 37875 34561 37887 34595
rect 37829 34555 37887 34561
rect 20533 34527 20591 34533
rect 20533 34493 20545 34527
rect 20579 34524 20591 34527
rect 25498 34524 25504 34536
rect 20579 34496 25504 34524
rect 20579 34493 20591 34496
rect 20533 34487 20591 34493
rect 25498 34484 25504 34496
rect 25556 34484 25562 34536
rect 32950 34524 32956 34536
rect 32911 34496 32956 34524
rect 32950 34484 32956 34496
rect 33008 34484 33014 34536
rect 33781 34527 33839 34533
rect 33781 34493 33793 34527
rect 33827 34524 33839 34527
rect 33962 34524 33968 34536
rect 33827 34496 33968 34524
rect 33827 34493 33839 34496
rect 33781 34487 33839 34493
rect 33962 34484 33968 34496
rect 34020 34484 34026 34536
rect 36906 34484 36912 34536
rect 36964 34524 36970 34536
rect 37844 34524 37872 34555
rect 36964 34496 37872 34524
rect 36964 34484 36970 34496
rect 23109 34459 23167 34465
rect 23109 34425 23121 34459
rect 23155 34425 23167 34459
rect 23109 34419 23167 34425
rect 5810 34388 5816 34400
rect 5771 34360 5816 34388
rect 5810 34348 5816 34360
rect 5868 34348 5874 34400
rect 19426 34388 19432 34400
rect 19387 34360 19432 34388
rect 19426 34348 19432 34360
rect 19484 34348 19490 34400
rect 22370 34388 22376 34400
rect 22331 34360 22376 34388
rect 22370 34348 22376 34360
rect 22428 34388 22434 34400
rect 23124 34388 23152 34419
rect 23934 34416 23940 34468
rect 23992 34456 23998 34468
rect 24029 34459 24087 34465
rect 24029 34456 24041 34459
rect 23992 34428 24041 34456
rect 23992 34416 23998 34428
rect 24029 34425 24041 34428
rect 24075 34425 24087 34459
rect 24029 34419 24087 34425
rect 22428 34360 23152 34388
rect 22428 34348 22434 34360
rect 35802 34348 35808 34400
rect 35860 34388 35866 34400
rect 35989 34391 36047 34397
rect 35989 34388 36001 34391
rect 35860 34360 36001 34388
rect 35860 34348 35866 34360
rect 35989 34357 36001 34360
rect 36035 34357 36047 34391
rect 35989 34351 36047 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 18046 34184 18052 34196
rect 18007 34156 18052 34184
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 31294 34184 31300 34196
rect 31255 34156 31300 34184
rect 31294 34144 31300 34156
rect 31352 34144 31358 34196
rect 35897 34187 35955 34193
rect 35897 34153 35909 34187
rect 35943 34184 35955 34187
rect 35986 34184 35992 34196
rect 35943 34156 35992 34184
rect 35943 34153 35955 34156
rect 35897 34147 35955 34153
rect 35986 34144 35992 34156
rect 36044 34144 36050 34196
rect 36078 34144 36084 34196
rect 36136 34184 36142 34196
rect 36357 34187 36415 34193
rect 36357 34184 36369 34187
rect 36136 34156 36369 34184
rect 36136 34144 36142 34156
rect 36357 34153 36369 34156
rect 36403 34153 36415 34187
rect 37182 34184 37188 34196
rect 37143 34156 37188 34184
rect 36357 34147 36415 34153
rect 37182 34144 37188 34156
rect 37240 34144 37246 34196
rect 37642 34144 37648 34196
rect 37700 34184 37706 34196
rect 37921 34187 37979 34193
rect 37921 34184 37933 34187
rect 37700 34156 37933 34184
rect 37700 34144 37706 34156
rect 37921 34153 37933 34156
rect 37967 34153 37979 34187
rect 37921 34147 37979 34153
rect 36722 34048 36728 34060
rect 36556 34020 36728 34048
rect 9401 33983 9459 33989
rect 9401 33949 9413 33983
rect 9447 33980 9459 33983
rect 9490 33980 9496 33992
rect 9447 33952 9496 33980
rect 9447 33949 9459 33952
rect 9401 33943 9459 33949
rect 9490 33940 9496 33952
rect 9548 33980 9554 33992
rect 31481 33983 31539 33989
rect 9548 33952 11376 33980
rect 9548 33940 9554 33952
rect 9668 33915 9726 33921
rect 9668 33881 9680 33915
rect 9714 33912 9726 33915
rect 10134 33912 10140 33924
rect 9714 33884 10140 33912
rect 9714 33881 9726 33884
rect 9668 33875 9726 33881
rect 10134 33872 10140 33884
rect 10192 33872 10198 33924
rect 10778 33844 10784 33856
rect 10739 33816 10784 33844
rect 10778 33804 10784 33816
rect 10836 33804 10842 33856
rect 11348 33853 11376 33952
rect 31481 33949 31493 33983
rect 31527 33980 31539 33983
rect 32122 33980 32128 33992
rect 31527 33952 32128 33980
rect 31527 33949 31539 33952
rect 31481 33943 31539 33949
rect 32122 33940 32128 33952
rect 32180 33940 32186 33992
rect 36556 33989 36584 34020
rect 36722 34008 36728 34020
rect 36780 34008 36786 34060
rect 36541 33983 36599 33989
rect 36541 33949 36553 33983
rect 36587 33949 36599 33983
rect 36541 33943 36599 33949
rect 36630 33940 36636 33992
rect 36688 33980 36694 33992
rect 37001 33983 37059 33989
rect 37001 33980 37013 33983
rect 36688 33952 37013 33980
rect 36688 33940 36694 33952
rect 37001 33949 37013 33952
rect 37047 33949 37059 33983
rect 37734 33980 37740 33992
rect 37695 33952 37740 33980
rect 37001 33943 37059 33949
rect 37734 33940 37740 33952
rect 37792 33940 37798 33992
rect 11333 33847 11391 33853
rect 11333 33813 11345 33847
rect 11379 33844 11391 33847
rect 13722 33844 13728 33856
rect 11379 33816 13728 33844
rect 11379 33813 11391 33816
rect 11333 33807 11391 33813
rect 13722 33804 13728 33816
rect 13780 33804 13786 33856
rect 15930 33844 15936 33856
rect 15891 33816 15936 33844
rect 15930 33804 15936 33816
rect 15988 33804 15994 33856
rect 17126 33844 17132 33856
rect 17087 33816 17132 33844
rect 17126 33804 17132 33816
rect 17184 33804 17190 33856
rect 23661 33847 23719 33853
rect 23661 33813 23673 33847
rect 23707 33844 23719 33847
rect 23934 33844 23940 33856
rect 23707 33816 23940 33844
rect 23707 33813 23719 33816
rect 23661 33807 23719 33813
rect 23934 33804 23940 33816
rect 23992 33804 23998 33856
rect 33594 33804 33600 33856
rect 33652 33844 33658 33856
rect 33873 33847 33931 33853
rect 33873 33844 33885 33847
rect 33652 33816 33885 33844
rect 33652 33804 33658 33816
rect 33873 33813 33885 33816
rect 33919 33844 33931 33847
rect 34054 33844 34060 33856
rect 33919 33816 34060 33844
rect 33919 33813 33931 33816
rect 33873 33807 33931 33813
rect 34054 33804 34060 33816
rect 34112 33804 34118 33856
rect 34606 33804 34612 33856
rect 34664 33844 34670 33856
rect 34701 33847 34759 33853
rect 34701 33844 34713 33847
rect 34664 33816 34713 33844
rect 34664 33804 34670 33816
rect 34701 33813 34713 33816
rect 34747 33813 34759 33847
rect 34701 33807 34759 33813
rect 35345 33847 35403 33853
rect 35345 33813 35357 33847
rect 35391 33844 35403 33847
rect 35434 33844 35440 33856
rect 35391 33816 35440 33844
rect 35391 33813 35403 33816
rect 35345 33807 35403 33813
rect 35434 33804 35440 33816
rect 35492 33804 35498 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 5258 33640 5264 33652
rect 5219 33612 5264 33640
rect 5258 33600 5264 33612
rect 5316 33600 5322 33652
rect 10134 33640 10140 33652
rect 10095 33612 10140 33640
rect 10134 33600 10140 33612
rect 10192 33600 10198 33652
rect 10778 33600 10784 33652
rect 10836 33640 10842 33652
rect 11609 33643 11667 33649
rect 11609 33640 11621 33643
rect 10836 33612 11621 33640
rect 10836 33600 10842 33612
rect 11609 33609 11621 33612
rect 11655 33640 11667 33643
rect 11790 33640 11796 33652
rect 11655 33612 11796 33640
rect 11655 33609 11667 33612
rect 11609 33603 11667 33609
rect 11790 33600 11796 33612
rect 11848 33600 11854 33652
rect 18322 33600 18328 33652
rect 18380 33640 18386 33652
rect 18417 33643 18475 33649
rect 18417 33640 18429 33643
rect 18380 33612 18429 33640
rect 18380 33600 18386 33612
rect 18417 33609 18429 33612
rect 18463 33609 18475 33643
rect 29362 33640 29368 33652
rect 29323 33612 29368 33640
rect 18417 33603 18475 33609
rect 29362 33600 29368 33612
rect 29420 33600 29426 33652
rect 36722 33640 36728 33652
rect 36683 33612 36728 33640
rect 36722 33600 36728 33612
rect 36780 33600 36786 33652
rect 37369 33643 37427 33649
rect 37369 33609 37381 33643
rect 37415 33640 37427 33643
rect 37826 33640 37832 33652
rect 37415 33612 37832 33640
rect 37415 33609 37427 33612
rect 37369 33603 37427 33609
rect 37826 33600 37832 33612
rect 37884 33600 37890 33652
rect 38013 33643 38071 33649
rect 38013 33609 38025 33643
rect 38059 33640 38071 33643
rect 38654 33640 38660 33652
rect 38059 33612 38660 33640
rect 38059 33609 38071 33612
rect 38013 33603 38071 33609
rect 38654 33600 38660 33612
rect 38712 33600 38718 33652
rect 10244 33544 11560 33572
rect 5445 33507 5503 33513
rect 5445 33473 5457 33507
rect 5491 33504 5503 33507
rect 6822 33504 6828 33516
rect 5491 33476 6828 33504
rect 5491 33473 5503 33476
rect 5445 33467 5503 33473
rect 6822 33464 6828 33476
rect 6880 33464 6886 33516
rect 4890 33396 4896 33448
rect 4948 33436 4954 33448
rect 5166 33436 5172 33448
rect 4948 33408 5172 33436
rect 4948 33396 4954 33408
rect 5166 33396 5172 33408
rect 5224 33396 5230 33448
rect 5721 33439 5779 33445
rect 5721 33405 5733 33439
rect 5767 33436 5779 33439
rect 5810 33436 5816 33448
rect 5767 33408 5816 33436
rect 5767 33405 5779 33408
rect 5721 33399 5779 33405
rect 5810 33396 5816 33408
rect 5868 33436 5874 33448
rect 6362 33436 6368 33448
rect 5868 33408 6368 33436
rect 5868 33396 5874 33408
rect 6362 33396 6368 33408
rect 6420 33396 6426 33448
rect 4798 33260 4804 33312
rect 4856 33300 4862 33312
rect 5629 33303 5687 33309
rect 5629 33300 5641 33303
rect 4856 33272 5641 33300
rect 4856 33260 4862 33272
rect 5629 33269 5641 33272
rect 5675 33269 5687 33303
rect 5629 33263 5687 33269
rect 7650 33260 7656 33312
rect 7708 33300 7714 33312
rect 10244 33300 10272 33544
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33473 10379 33507
rect 10321 33467 10379 33473
rect 10597 33507 10655 33513
rect 10597 33473 10609 33507
rect 10643 33504 10655 33507
rect 10778 33504 10784 33516
rect 10643 33476 10784 33504
rect 10643 33473 10655 33476
rect 10597 33467 10655 33473
rect 10336 33368 10364 33467
rect 10778 33464 10784 33476
rect 10836 33464 10842 33516
rect 11532 33513 11560 33544
rect 11517 33507 11575 33513
rect 11517 33473 11529 33507
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 11793 33507 11851 33513
rect 11793 33473 11805 33507
rect 11839 33504 11851 33507
rect 18601 33507 18659 33513
rect 11839 33476 12388 33504
rect 11839 33473 11851 33476
rect 11793 33467 11851 33473
rect 12360 33377 12388 33476
rect 18601 33473 18613 33507
rect 18647 33504 18659 33507
rect 19518 33504 19524 33516
rect 18647 33476 19524 33504
rect 18647 33473 18659 33476
rect 18601 33467 18659 33473
rect 19518 33464 19524 33476
rect 19576 33464 19582 33516
rect 27522 33504 27528 33516
rect 27483 33476 27528 33504
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 29178 33504 29184 33516
rect 29139 33476 29184 33504
rect 29178 33464 29184 33476
rect 29236 33464 29242 33516
rect 37826 33504 37832 33516
rect 37787 33476 37832 33504
rect 37826 33464 37832 33476
rect 37884 33464 37890 33516
rect 18877 33439 18935 33445
rect 18877 33405 18889 33439
rect 18923 33436 18935 33439
rect 19426 33436 19432 33448
rect 18923 33408 19432 33436
rect 18923 33405 18935 33408
rect 18877 33399 18935 33405
rect 19426 33396 19432 33408
rect 19484 33396 19490 33448
rect 27798 33436 27804 33448
rect 27759 33408 27804 33436
rect 27798 33396 27804 33408
rect 27856 33396 27862 33448
rect 11793 33371 11851 33377
rect 11793 33368 11805 33371
rect 10336 33340 11805 33368
rect 11793 33337 11805 33340
rect 11839 33337 11851 33371
rect 11793 33331 11851 33337
rect 12345 33371 12403 33377
rect 12345 33337 12357 33371
rect 12391 33368 12403 33371
rect 19334 33368 19340 33380
rect 12391 33340 19340 33368
rect 12391 33337 12403 33340
rect 12345 33331 12403 33337
rect 19334 33328 19340 33340
rect 19392 33328 19398 33380
rect 10505 33303 10563 33309
rect 10505 33300 10517 33303
rect 7708 33272 10517 33300
rect 7708 33260 7714 33272
rect 10505 33269 10517 33272
rect 10551 33269 10563 33303
rect 10505 33263 10563 33269
rect 18785 33303 18843 33309
rect 18785 33269 18797 33303
rect 18831 33300 18843 33303
rect 19242 33300 19248 33312
rect 18831 33272 19248 33300
rect 18831 33269 18843 33272
rect 18785 33263 18843 33269
rect 19242 33260 19248 33272
rect 19300 33260 19306 33312
rect 35345 33303 35403 33309
rect 35345 33269 35357 33303
rect 35391 33300 35403 33303
rect 35526 33300 35532 33312
rect 35391 33272 35532 33300
rect 35391 33269 35403 33272
rect 35345 33263 35403 33269
rect 35526 33260 35532 33272
rect 35584 33260 35590 33312
rect 36173 33303 36231 33309
rect 36173 33269 36185 33303
rect 36219 33300 36231 33303
rect 36354 33300 36360 33312
rect 36219 33272 36360 33300
rect 36219 33269 36231 33272
rect 36173 33263 36231 33269
rect 36354 33260 36360 33272
rect 36412 33260 36418 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 19518 33096 19524 33108
rect 19479 33068 19524 33096
rect 19518 33056 19524 33068
rect 19576 33056 19582 33108
rect 28442 33028 28448 33040
rect 28403 33000 28448 33028
rect 28442 32988 28448 33000
rect 28500 32988 28506 33040
rect 19242 32892 19248 32904
rect 19203 32864 19248 32892
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 19337 32895 19395 32901
rect 19337 32861 19349 32895
rect 19383 32892 19395 32895
rect 19426 32892 19432 32904
rect 19383 32864 19432 32892
rect 19383 32861 19395 32864
rect 19337 32855 19395 32861
rect 19426 32852 19432 32864
rect 19484 32852 19490 32904
rect 27798 32852 27804 32904
rect 27856 32892 27862 32904
rect 28261 32895 28319 32901
rect 28261 32892 28273 32895
rect 27856 32864 28273 32892
rect 27856 32852 27862 32864
rect 28261 32861 28273 32864
rect 28307 32892 28319 32895
rect 32858 32892 32864 32904
rect 28307 32864 32864 32892
rect 28307 32861 28319 32864
rect 28261 32855 28319 32861
rect 32858 32852 32864 32864
rect 32916 32892 32922 32904
rect 37829 32895 37887 32901
rect 37829 32892 37841 32895
rect 32916 32864 37841 32892
rect 32916 32852 32922 32864
rect 37829 32861 37841 32864
rect 37875 32861 37887 32895
rect 38102 32892 38108 32904
rect 38063 32864 38108 32892
rect 37829 32855 37887 32861
rect 38102 32852 38108 32864
rect 38160 32852 38166 32904
rect 19521 32827 19579 32833
rect 19521 32793 19533 32827
rect 19567 32793 19579 32827
rect 19521 32787 19579 32793
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 19536 32756 19564 32787
rect 19978 32756 19984 32768
rect 19392 32728 19984 32756
rect 19392 32716 19398 32728
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 36265 32759 36323 32765
rect 36265 32725 36277 32759
rect 36311 32756 36323 32759
rect 36538 32756 36544 32768
rect 36311 32728 36544 32756
rect 36311 32725 36323 32728
rect 36265 32719 36323 32725
rect 36538 32716 36544 32728
rect 36596 32716 36602 32768
rect 36817 32759 36875 32765
rect 36817 32725 36829 32759
rect 36863 32756 36875 32759
rect 36906 32756 36912 32768
rect 36863 32728 36912 32756
rect 36863 32725 36875 32728
rect 36817 32719 36875 32725
rect 36906 32716 36912 32728
rect 36964 32716 36970 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 6822 32552 6828 32564
rect 6783 32524 6828 32552
rect 6822 32512 6828 32524
rect 6880 32512 6886 32564
rect 26142 32552 26148 32564
rect 26103 32524 26148 32552
rect 26142 32512 26148 32524
rect 26200 32512 26206 32564
rect 32122 32552 32128 32564
rect 32083 32524 32128 32552
rect 32122 32512 32128 32524
rect 32180 32512 32186 32564
rect 38102 32484 38108 32496
rect 38063 32456 38108 32484
rect 38102 32444 38108 32456
rect 38160 32444 38166 32496
rect 6733 32419 6791 32425
rect 6733 32385 6745 32419
rect 6779 32385 6791 32419
rect 6733 32379 6791 32385
rect 6917 32419 6975 32425
rect 6917 32385 6929 32419
rect 6963 32416 6975 32419
rect 7650 32416 7656 32428
rect 6963 32388 7656 32416
rect 6963 32385 6975 32388
rect 6917 32379 6975 32385
rect 6748 32348 6776 32379
rect 7650 32376 7656 32388
rect 7708 32376 7714 32428
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32416 13691 32419
rect 13722 32416 13728 32428
rect 13679 32388 13728 32416
rect 13679 32385 13691 32388
rect 13633 32379 13691 32385
rect 13722 32376 13728 32388
rect 13780 32416 13786 32428
rect 14366 32425 14372 32428
rect 14093 32419 14151 32425
rect 14093 32416 14105 32419
rect 13780 32388 14105 32416
rect 13780 32376 13786 32388
rect 14093 32385 14105 32388
rect 14139 32385 14151 32419
rect 14093 32379 14151 32385
rect 14360 32379 14372 32425
rect 14424 32416 14430 32428
rect 14424 32388 14460 32416
rect 14366 32376 14372 32379
rect 14424 32376 14430 32388
rect 25314 32376 25320 32428
rect 25372 32416 25378 32428
rect 25777 32419 25835 32425
rect 25777 32416 25789 32419
rect 25372 32388 25789 32416
rect 25372 32376 25378 32388
rect 25777 32385 25789 32388
rect 25823 32385 25835 32419
rect 25777 32379 25835 32385
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32416 26019 32419
rect 26234 32416 26240 32428
rect 26007 32388 26240 32416
rect 26007 32385 26019 32388
rect 25961 32379 26019 32385
rect 26234 32376 26240 32388
rect 26292 32376 26298 32428
rect 32493 32419 32551 32425
rect 32493 32416 32505 32419
rect 31496 32388 32505 32416
rect 6748 32320 6914 32348
rect 6886 32212 6914 32320
rect 18782 32240 18788 32292
rect 18840 32280 18846 32292
rect 31496 32289 31524 32388
rect 32493 32385 32505 32388
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32585 32419 32643 32425
rect 32585 32385 32597 32419
rect 32631 32416 32643 32419
rect 34238 32416 34244 32428
rect 32631 32388 34244 32416
rect 32631 32385 32643 32388
rect 32585 32379 32643 32385
rect 34238 32376 34244 32388
rect 34296 32376 34302 32428
rect 32769 32351 32827 32357
rect 32769 32317 32781 32351
rect 32815 32348 32827 32351
rect 32858 32348 32864 32360
rect 32815 32320 32864 32348
rect 32815 32317 32827 32320
rect 32769 32311 32827 32317
rect 32858 32308 32864 32320
rect 32916 32308 32922 32360
rect 31481 32283 31539 32289
rect 31481 32280 31493 32283
rect 18840 32252 31493 32280
rect 18840 32240 18846 32252
rect 31481 32249 31493 32252
rect 31527 32249 31539 32283
rect 31481 32243 31539 32249
rect 7466 32212 7472 32224
rect 6886 32184 7472 32212
rect 7466 32172 7472 32184
rect 7524 32172 7530 32224
rect 15194 32172 15200 32224
rect 15252 32212 15258 32224
rect 15473 32215 15531 32221
rect 15473 32212 15485 32215
rect 15252 32184 15485 32212
rect 15252 32172 15258 32184
rect 15473 32181 15485 32184
rect 15519 32181 15531 32215
rect 25314 32212 25320 32224
rect 25275 32184 25320 32212
rect 15473 32175 15531 32181
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 37553 32215 37611 32221
rect 37553 32181 37565 32215
rect 37599 32212 37611 32215
rect 37734 32212 37740 32224
rect 37599 32184 37740 32212
rect 37599 32181 37611 32184
rect 37553 32175 37611 32181
rect 37734 32172 37740 32184
rect 37792 32212 37798 32224
rect 38654 32212 38660 32224
rect 37792 32184 38660 32212
rect 37792 32172 37798 32184
rect 38654 32172 38660 32184
rect 38712 32172 38718 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 26513 32011 26571 32017
rect 26513 31977 26525 32011
rect 26559 32008 26571 32011
rect 26602 32008 26608 32020
rect 26559 31980 26608 32008
rect 26559 31977 26571 31980
rect 26513 31971 26571 31977
rect 26602 31968 26608 31980
rect 26660 31968 26666 32020
rect 28353 32011 28411 32017
rect 28353 31977 28365 32011
rect 28399 32008 28411 32011
rect 29178 32008 29184 32020
rect 28399 31980 29184 32008
rect 28399 31977 28411 31980
rect 28353 31971 28411 31977
rect 29178 31968 29184 31980
rect 29236 31968 29242 32020
rect 26234 31832 26240 31884
rect 26292 31872 26298 31884
rect 27522 31872 27528 31884
rect 26292 31844 27528 31872
rect 26292 31832 26298 31844
rect 25685 31807 25743 31813
rect 25685 31773 25697 31807
rect 25731 31804 25743 31807
rect 25866 31804 25872 31816
rect 25731 31776 25872 31804
rect 25731 31773 25743 31776
rect 25685 31767 25743 31773
rect 25866 31764 25872 31776
rect 25924 31804 25930 31816
rect 26344 31813 26372 31844
rect 27522 31832 27528 31844
rect 27580 31872 27586 31884
rect 27580 31844 28212 31872
rect 27580 31832 27586 31844
rect 26145 31807 26203 31813
rect 26145 31804 26157 31807
rect 25924 31776 26157 31804
rect 25924 31764 25930 31776
rect 26145 31773 26157 31776
rect 26191 31773 26203 31807
rect 26145 31767 26203 31773
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31773 26387 31807
rect 26329 31767 26387 31773
rect 26694 31764 26700 31816
rect 26752 31804 26758 31816
rect 28184 31813 28212 31844
rect 27433 31807 27491 31813
rect 27433 31804 27445 31807
rect 26752 31776 27445 31804
rect 26752 31764 26758 31776
rect 27433 31773 27445 31776
rect 27479 31804 27491 31807
rect 27985 31807 28043 31813
rect 27985 31804 27997 31807
rect 27479 31776 27997 31804
rect 27479 31773 27491 31776
rect 27433 31767 27491 31773
rect 27985 31773 27997 31776
rect 28031 31773 28043 31807
rect 27985 31767 28043 31773
rect 28169 31807 28227 31813
rect 28169 31773 28181 31807
rect 28215 31804 28227 31807
rect 28442 31804 28448 31816
rect 28215 31776 28448 31804
rect 28215 31773 28227 31776
rect 28169 31767 28227 31773
rect 28442 31764 28448 31776
rect 28500 31764 28506 31816
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 34885 31467 34943 31473
rect 34885 31433 34897 31467
rect 34931 31433 34943 31467
rect 34885 31427 34943 31433
rect 33042 31288 33048 31340
rect 33100 31328 33106 31340
rect 34701 31331 34759 31337
rect 34701 31328 34713 31331
rect 33100 31300 34713 31328
rect 33100 31288 33106 31300
rect 34701 31297 34713 31300
rect 34747 31297 34759 31331
rect 34900 31328 34928 31427
rect 35986 31356 35992 31408
rect 36044 31396 36050 31408
rect 36044 31368 36768 31396
rect 36044 31356 36050 31368
rect 36446 31328 36452 31340
rect 36504 31337 36510 31340
rect 36740 31337 36768 31368
rect 34900 31300 36452 31328
rect 34701 31291 34759 31297
rect 36446 31288 36452 31300
rect 36504 31291 36516 31337
rect 36725 31331 36783 31337
rect 36725 31297 36737 31331
rect 36771 31297 36783 31331
rect 36725 31291 36783 31297
rect 37461 31331 37519 31337
rect 37461 31297 37473 31331
rect 37507 31328 37519 31331
rect 38102 31328 38108 31340
rect 37507 31300 38108 31328
rect 37507 31297 37519 31300
rect 37461 31291 37519 31297
rect 36504 31288 36510 31291
rect 38102 31288 38108 31300
rect 38160 31288 38166 31340
rect 34238 31152 34244 31204
rect 34296 31192 34302 31204
rect 34296 31164 35848 31192
rect 34296 31152 34302 31164
rect 33134 31084 33140 31136
rect 33192 31124 33198 31136
rect 35345 31127 35403 31133
rect 35345 31124 35357 31127
rect 33192 31096 35357 31124
rect 33192 31084 33198 31096
rect 35345 31093 35357 31096
rect 35391 31093 35403 31127
rect 35820 31124 35848 31164
rect 37921 31127 37979 31133
rect 37921 31124 37933 31127
rect 35820 31096 37933 31124
rect 35345 31087 35403 31093
rect 37921 31093 37933 31096
rect 37967 31093 37979 31127
rect 37921 31087 37979 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 27062 30920 27068 30932
rect 27023 30892 27068 30920
rect 27062 30880 27068 30892
rect 27120 30880 27126 30932
rect 33042 30920 33048 30932
rect 33003 30892 33048 30920
rect 33042 30880 33048 30892
rect 33100 30880 33106 30932
rect 34422 30880 34428 30932
rect 34480 30920 34486 30932
rect 35253 30923 35311 30929
rect 35253 30920 35265 30923
rect 34480 30892 35265 30920
rect 34480 30880 34486 30892
rect 35253 30889 35265 30892
rect 35299 30920 35311 30923
rect 35986 30920 35992 30932
rect 35299 30892 35992 30920
rect 35299 30889 35311 30892
rect 35253 30883 35311 30889
rect 35986 30880 35992 30892
rect 36044 30880 36050 30932
rect 27522 30812 27528 30864
rect 27580 30812 27586 30864
rect 32858 30852 32864 30864
rect 32819 30824 32864 30852
rect 32858 30812 32864 30824
rect 32916 30812 32922 30864
rect 27540 30784 27568 30812
rect 27617 30787 27675 30793
rect 27617 30784 27629 30787
rect 27540 30756 27629 30784
rect 27617 30753 27629 30756
rect 27663 30753 27675 30787
rect 27617 30747 27675 30753
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 1903 30688 3801 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 3789 30685 3801 30688
rect 3835 30716 3847 30719
rect 4062 30716 4068 30728
rect 3835 30688 4068 30716
rect 3835 30685 3847 30688
rect 3789 30679 3847 30685
rect 4062 30676 4068 30688
rect 4120 30676 4126 30728
rect 4798 30716 4804 30728
rect 4759 30688 4804 30716
rect 4798 30676 4804 30688
rect 4856 30676 4862 30728
rect 4985 30719 5043 30725
rect 4985 30685 4997 30719
rect 5031 30716 5043 30719
rect 23661 30719 23719 30725
rect 5031 30688 5580 30716
rect 5031 30685 5043 30688
rect 4985 30679 5043 30685
rect 2124 30651 2182 30657
rect 2124 30617 2136 30651
rect 2170 30648 2182 30651
rect 3602 30648 3608 30660
rect 2170 30620 3608 30648
rect 2170 30617 2182 30620
rect 2124 30611 2182 30617
rect 3602 30608 3608 30620
rect 3660 30608 3666 30660
rect 3237 30583 3295 30589
rect 3237 30549 3249 30583
rect 3283 30580 3295 30583
rect 4062 30580 4068 30592
rect 3283 30552 4068 30580
rect 3283 30549 3295 30552
rect 3237 30543 3295 30549
rect 4062 30540 4068 30552
rect 4120 30540 4126 30592
rect 4890 30580 4896 30592
rect 4851 30552 4896 30580
rect 4890 30540 4896 30552
rect 4948 30540 4954 30592
rect 5552 30589 5580 30688
rect 23661 30685 23673 30719
rect 23707 30716 23719 30719
rect 27525 30719 27583 30725
rect 23707 30688 24532 30716
rect 23707 30685 23719 30688
rect 23661 30679 23719 30685
rect 22738 30608 22744 30660
rect 22796 30648 22802 30660
rect 24504 30657 24532 30688
rect 27525 30685 27537 30719
rect 27571 30716 27583 30719
rect 37182 30716 37188 30728
rect 27571 30688 37188 30716
rect 27571 30685 27583 30688
rect 27525 30679 27583 30685
rect 37182 30676 37188 30688
rect 37240 30676 37246 30728
rect 23394 30651 23452 30657
rect 23394 30648 23406 30651
rect 22796 30620 23406 30648
rect 22796 30608 22802 30620
rect 23394 30617 23406 30620
rect 23440 30617 23452 30651
rect 23394 30611 23452 30617
rect 24489 30651 24547 30657
rect 24489 30617 24501 30651
rect 24535 30648 24547 30651
rect 27154 30648 27160 30660
rect 24535 30620 27160 30648
rect 24535 30617 24547 30620
rect 24489 30611 24547 30617
rect 27154 30608 27160 30620
rect 27212 30608 27218 30660
rect 32582 30648 32588 30660
rect 32543 30620 32588 30648
rect 32582 30608 32588 30620
rect 32640 30608 32646 30660
rect 5537 30583 5595 30589
rect 5537 30549 5549 30583
rect 5583 30580 5595 30583
rect 6914 30580 6920 30592
rect 5583 30552 6920 30580
rect 5583 30549 5595 30552
rect 5537 30543 5595 30549
rect 6914 30540 6920 30552
rect 6972 30580 6978 30592
rect 7466 30580 7472 30592
rect 6972 30552 7472 30580
rect 6972 30540 6978 30552
rect 7466 30540 7472 30552
rect 7524 30580 7530 30592
rect 8202 30580 8208 30592
rect 7524 30552 8208 30580
rect 7524 30540 7530 30552
rect 8202 30540 8208 30552
rect 8260 30540 8266 30592
rect 22278 30580 22284 30592
rect 22239 30552 22284 30580
rect 22278 30540 22284 30552
rect 22336 30540 22342 30592
rect 26605 30583 26663 30589
rect 26605 30549 26617 30583
rect 26651 30580 26663 30583
rect 27338 30580 27344 30592
rect 26651 30552 27344 30580
rect 26651 30549 26663 30552
rect 26605 30543 26663 30549
rect 27338 30540 27344 30552
rect 27396 30580 27402 30592
rect 27433 30583 27491 30589
rect 27433 30580 27445 30583
rect 27396 30552 27445 30580
rect 27396 30540 27402 30552
rect 27433 30549 27445 30552
rect 27479 30549 27491 30583
rect 27433 30543 27491 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 4798 30336 4804 30388
rect 4856 30376 4862 30388
rect 4985 30379 5043 30385
rect 4985 30376 4997 30379
rect 4856 30348 4997 30376
rect 4856 30336 4862 30348
rect 4985 30345 4997 30348
rect 5031 30345 5043 30379
rect 4985 30339 5043 30345
rect 5276 30348 5488 30376
rect 3602 30308 3608 30320
rect 3563 30280 3608 30308
rect 3602 30268 3608 30280
rect 3660 30268 3666 30320
rect 5153 30311 5211 30317
rect 5153 30277 5165 30311
rect 5199 30308 5211 30311
rect 5276 30308 5304 30348
rect 5199 30280 5304 30308
rect 5353 30311 5411 30317
rect 5199 30277 5211 30280
rect 5153 30271 5211 30277
rect 5353 30277 5365 30311
rect 5399 30277 5411 30311
rect 5460 30308 5488 30348
rect 6196 30348 6500 30376
rect 5626 30308 5632 30320
rect 5460 30280 5632 30308
rect 5353 30271 5411 30277
rect 1578 30200 1584 30252
rect 1636 30240 1642 30252
rect 1857 30243 1915 30249
rect 1857 30240 1869 30243
rect 1636 30212 1869 30240
rect 1636 30200 1642 30212
rect 1857 30209 1869 30212
rect 1903 30209 1915 30243
rect 1857 30203 1915 30209
rect 3789 30243 3847 30249
rect 3789 30209 3801 30243
rect 3835 30240 3847 30243
rect 4890 30240 4896 30252
rect 3835 30212 4896 30240
rect 3835 30209 3847 30212
rect 3789 30203 3847 30209
rect 4890 30200 4896 30212
rect 4948 30200 4954 30252
rect 5368 30240 5396 30271
rect 5626 30268 5632 30280
rect 5684 30308 5690 30320
rect 6196 30308 6224 30348
rect 6362 30308 6368 30320
rect 5684 30280 6224 30308
rect 6323 30280 6368 30308
rect 5684 30268 5690 30280
rect 6362 30268 6368 30280
rect 6420 30268 6426 30320
rect 6472 30308 6500 30348
rect 11440 30348 11744 30376
rect 6733 30311 6791 30317
rect 6733 30308 6745 30311
rect 6472 30280 6745 30308
rect 6733 30277 6745 30280
rect 6779 30277 6791 30311
rect 6733 30271 6791 30277
rect 7650 30268 7656 30320
rect 7708 30308 7714 30320
rect 8021 30311 8079 30317
rect 8021 30308 8033 30311
rect 7708 30280 8033 30308
rect 7708 30268 7714 30280
rect 8021 30277 8033 30280
rect 8067 30308 8079 30311
rect 10962 30308 10968 30320
rect 8067 30280 10968 30308
rect 8067 30277 8079 30280
rect 8021 30271 8079 30277
rect 10962 30268 10968 30280
rect 11020 30308 11026 30320
rect 11440 30308 11468 30348
rect 11020 30280 11468 30308
rect 11020 30268 11026 30280
rect 11514 30268 11520 30320
rect 11572 30308 11578 30320
rect 11716 30317 11744 30348
rect 11882 30336 11888 30388
rect 11940 30376 11946 30388
rect 12897 30379 12955 30385
rect 12897 30376 12909 30379
rect 11940 30348 12909 30376
rect 11940 30336 11946 30348
rect 12897 30345 12909 30348
rect 12943 30345 12955 30379
rect 12897 30339 12955 30345
rect 15378 30336 15384 30388
rect 15436 30376 15442 30388
rect 16025 30379 16083 30385
rect 16025 30376 16037 30379
rect 15436 30348 16037 30376
rect 15436 30336 15442 30348
rect 16025 30345 16037 30348
rect 16071 30345 16083 30379
rect 22738 30376 22744 30388
rect 22699 30348 22744 30376
rect 16025 30339 16083 30345
rect 22738 30336 22744 30348
rect 22796 30336 22802 30388
rect 32398 30376 32404 30388
rect 32359 30348 32404 30376
rect 32398 30336 32404 30348
rect 32456 30336 32462 30388
rect 32582 30336 32588 30388
rect 32640 30376 32646 30388
rect 32769 30379 32827 30385
rect 32769 30376 32781 30379
rect 32640 30348 32781 30376
rect 32640 30336 32646 30348
rect 32769 30345 32781 30348
rect 32815 30345 32827 30379
rect 32769 30339 32827 30345
rect 11716 30311 11775 30317
rect 11572 30280 11617 30308
rect 11716 30280 11729 30311
rect 11572 30268 11578 30280
rect 11717 30277 11729 30280
rect 11763 30277 11775 30311
rect 12989 30311 13047 30317
rect 12989 30308 13001 30311
rect 11717 30271 11775 30277
rect 11808 30280 13001 30308
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 5368 30212 6561 30240
rect 4062 30172 4068 30184
rect 4023 30144 4068 30172
rect 4062 30132 4068 30144
rect 4120 30172 4126 30184
rect 5368 30172 5396 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 6641 30243 6699 30249
rect 6641 30209 6653 30243
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30240 6975 30243
rect 7837 30243 7895 30249
rect 7837 30240 7849 30243
rect 6963 30212 7849 30240
rect 6963 30209 6975 30212
rect 6917 30203 6975 30209
rect 7837 30209 7849 30212
rect 7883 30240 7895 30243
rect 11808 30240 11836 30280
rect 12989 30277 13001 30280
rect 13035 30277 13047 30311
rect 14366 30308 14372 30320
rect 14327 30280 14372 30308
rect 12989 30271 13047 30277
rect 14366 30268 14372 30280
rect 14424 30268 14430 30320
rect 15473 30311 15531 30317
rect 15473 30308 15485 30311
rect 14568 30280 15485 30308
rect 14568 30249 14596 30280
rect 15473 30277 15485 30280
rect 15519 30277 15531 30311
rect 19137 30311 19195 30317
rect 19137 30308 19149 30311
rect 15473 30271 15531 30277
rect 18248 30280 19149 30308
rect 12805 30243 12863 30249
rect 12805 30240 12817 30243
rect 7883 30212 11836 30240
rect 11900 30212 12817 30240
rect 7883 30209 7895 30212
rect 7837 30203 7895 30209
rect 4120 30144 5396 30172
rect 4120 30132 4126 30144
rect 2133 30107 2191 30113
rect 2133 30073 2145 30107
rect 2179 30104 2191 30107
rect 6178 30104 6184 30116
rect 2179 30076 6184 30104
rect 2179 30073 2191 30076
rect 2133 30067 2191 30073
rect 6178 30064 6184 30076
rect 6236 30064 6242 30116
rect 3973 30039 4031 30045
rect 3973 30005 3985 30039
rect 4019 30036 4031 30039
rect 4798 30036 4804 30048
rect 4019 30008 4804 30036
rect 4019 30005 4031 30008
rect 3973 29999 4031 30005
rect 4798 29996 4804 30008
rect 4856 29996 4862 30048
rect 4890 29996 4896 30048
rect 4948 30036 4954 30048
rect 5169 30039 5227 30045
rect 5169 30036 5181 30039
rect 4948 30008 5181 30036
rect 4948 29996 4954 30008
rect 5169 30005 5181 30008
rect 5215 30036 5227 30039
rect 6656 30036 6684 30203
rect 11422 30132 11428 30184
rect 11480 30172 11486 30184
rect 11900 30172 11928 30212
rect 12805 30209 12817 30212
rect 12851 30209 12863 30243
rect 12805 30203 12863 30209
rect 14553 30243 14611 30249
rect 14553 30209 14565 30243
rect 14599 30209 14611 30243
rect 14553 30203 14611 30209
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30240 14887 30243
rect 15194 30240 15200 30252
rect 14875 30212 15200 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 14737 30175 14795 30181
rect 14737 30172 14749 30175
rect 11480 30144 11928 30172
rect 12406 30144 14749 30172
rect 11480 30132 11486 30144
rect 11606 30064 11612 30116
rect 11664 30104 11670 30116
rect 11885 30107 11943 30113
rect 11885 30104 11897 30107
rect 11664 30076 11897 30104
rect 11664 30064 11670 30076
rect 11885 30073 11897 30076
rect 11931 30104 11943 30107
rect 12406 30104 12434 30144
rect 14737 30141 14749 30144
rect 14783 30141 14795 30175
rect 14737 30135 14795 30141
rect 11931 30076 12434 30104
rect 12621 30107 12679 30113
rect 11931 30073 11943 30076
rect 11885 30067 11943 30073
rect 12621 30073 12633 30107
rect 12667 30104 12679 30107
rect 14844 30104 14872 30203
rect 15194 30200 15200 30212
rect 15252 30200 15258 30252
rect 15378 30240 15384 30252
rect 15339 30212 15384 30240
rect 15378 30200 15384 30212
rect 15436 30200 15442 30252
rect 18248 30249 18276 30280
rect 19137 30277 19149 30280
rect 19183 30308 19195 30311
rect 19242 30308 19248 30320
rect 19183 30280 19248 30308
rect 19183 30277 19195 30280
rect 19137 30271 19195 30277
rect 19242 30268 19248 30280
rect 19300 30268 19306 30320
rect 19337 30311 19395 30317
rect 19337 30277 19349 30311
rect 19383 30277 19395 30311
rect 19337 30271 19395 30277
rect 15577 30246 15635 30249
rect 15577 30243 15700 30246
rect 15577 30209 15589 30243
rect 15623 30240 15700 30243
rect 17221 30243 17279 30249
rect 17221 30240 17233 30243
rect 15623 30218 17233 30240
rect 15623 30209 15635 30218
rect 15672 30212 17233 30218
rect 15577 30203 15635 30209
rect 17221 30209 17233 30212
rect 17267 30240 17279 30243
rect 18233 30243 18291 30249
rect 18233 30240 18245 30243
rect 17267 30212 18245 30240
rect 17267 30209 17279 30212
rect 17221 30203 17279 30209
rect 18233 30209 18245 30212
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18325 30243 18383 30249
rect 18325 30209 18337 30243
rect 18371 30209 18383 30243
rect 18325 30203 18383 30209
rect 18509 30243 18567 30249
rect 18509 30209 18521 30243
rect 18555 30240 18567 30243
rect 18690 30240 18696 30252
rect 18555 30212 18696 30240
rect 18555 30209 18567 30212
rect 18509 30203 18567 30209
rect 15470 30132 15476 30184
rect 15528 30172 15534 30184
rect 17494 30172 17500 30184
rect 15528 30144 17500 30172
rect 15528 30132 15534 30144
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 18340 30172 18368 30203
rect 18690 30200 18696 30212
rect 18748 30240 18754 30252
rect 19352 30240 19380 30271
rect 19426 30268 19432 30320
rect 19484 30308 19490 30320
rect 20073 30311 20131 30317
rect 20073 30308 20085 30311
rect 19484 30280 20085 30308
rect 19484 30268 19490 30280
rect 20073 30277 20085 30280
rect 20119 30277 20131 30311
rect 20073 30271 20131 30277
rect 32030 30268 32036 30320
rect 32088 30308 32094 30320
rect 32217 30311 32275 30317
rect 32217 30308 32229 30311
rect 32088 30280 32229 30308
rect 32088 30268 32094 30280
rect 32217 30277 32229 30280
rect 32263 30308 32275 30311
rect 33134 30308 33140 30320
rect 32263 30280 33140 30308
rect 32263 30277 32275 30280
rect 32217 30271 32275 30277
rect 33134 30268 33140 30280
rect 33192 30268 33198 30320
rect 19981 30243 20039 30249
rect 19981 30240 19993 30243
rect 18748 30212 19993 30240
rect 18748 30200 18754 30212
rect 19981 30209 19993 30212
rect 20027 30209 20039 30243
rect 20162 30240 20168 30252
rect 20123 30212 20168 30240
rect 19981 30203 20039 30209
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 22557 30243 22615 30249
rect 22557 30209 22569 30243
rect 22603 30240 22615 30243
rect 22922 30240 22928 30252
rect 22603 30212 22928 30240
rect 22603 30209 22615 30212
rect 22557 30203 22615 30209
rect 22922 30200 22928 30212
rect 22980 30200 22986 30252
rect 30282 30200 30288 30252
rect 30340 30240 30346 30252
rect 32493 30243 32551 30249
rect 32493 30240 32505 30243
rect 30340 30212 32505 30240
rect 30340 30200 30346 30212
rect 32493 30209 32505 30212
rect 32539 30209 32551 30243
rect 32493 30203 32551 30209
rect 19426 30172 19432 30184
rect 18340 30144 19432 30172
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 19797 30175 19855 30181
rect 19797 30141 19809 30175
rect 19843 30172 19855 30175
rect 22278 30172 22284 30184
rect 19843 30144 22284 30172
rect 19843 30141 19855 30144
rect 19797 30135 19855 30141
rect 22278 30132 22284 30144
rect 22336 30132 22342 30184
rect 32122 30172 32128 30184
rect 32083 30144 32128 30172
rect 32122 30132 32128 30144
rect 32180 30132 32186 30184
rect 32585 30175 32643 30181
rect 32585 30141 32597 30175
rect 32631 30141 32643 30175
rect 32585 30135 32643 30141
rect 12667 30076 14872 30104
rect 12667 30073 12679 30076
rect 12621 30067 12679 30073
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 18969 30107 19027 30113
rect 18969 30104 18981 30107
rect 18380 30076 18981 30104
rect 18380 30064 18386 30076
rect 18969 30073 18981 30076
rect 19015 30104 19027 30107
rect 22373 30107 22431 30113
rect 22373 30104 22385 30107
rect 19015 30076 22385 30104
rect 19015 30073 19027 30076
rect 18969 30067 19027 30073
rect 22373 30073 22385 30076
rect 22419 30073 22431 30107
rect 32600 30104 32628 30135
rect 22373 30067 22431 30073
rect 31496 30076 32628 30104
rect 5215 30008 6684 30036
rect 11701 30039 11759 30045
rect 5215 30005 5227 30008
rect 5169 29999 5227 30005
rect 11701 30005 11713 30039
rect 11747 30036 11759 30039
rect 11790 30036 11796 30048
rect 11747 30008 11796 30036
rect 11747 30005 11759 30008
rect 11701 29999 11759 30005
rect 11790 29996 11796 30008
rect 11848 29996 11854 30048
rect 13173 30039 13231 30045
rect 13173 30005 13185 30039
rect 13219 30036 13231 30039
rect 15470 30036 15476 30048
rect 13219 30008 15476 30036
rect 13219 30005 13231 30008
rect 13173 29999 13231 30005
rect 15470 29996 15476 30008
rect 15528 29996 15534 30048
rect 18414 29996 18420 30048
rect 18472 30036 18478 30048
rect 18509 30039 18567 30045
rect 18509 30036 18521 30039
rect 18472 30008 18521 30036
rect 18472 29996 18478 30008
rect 18509 30005 18521 30008
rect 18555 30005 18567 30039
rect 18509 29999 18567 30005
rect 19153 30039 19211 30045
rect 19153 30005 19165 30039
rect 19199 30036 19211 30039
rect 19426 30036 19432 30048
rect 19199 30008 19432 30036
rect 19199 30005 19211 30008
rect 19153 29999 19211 30005
rect 19426 29996 19432 30008
rect 19484 29996 19490 30048
rect 20349 30039 20407 30045
rect 20349 30005 20361 30039
rect 20395 30036 20407 30039
rect 22278 30036 22284 30048
rect 20395 30008 22284 30036
rect 20395 30005 20407 30008
rect 20349 29999 20407 30005
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 30834 29996 30840 30048
rect 30892 30036 30898 30048
rect 31496 30045 31524 30076
rect 31481 30039 31539 30045
rect 31481 30036 31493 30039
rect 30892 30008 31493 30036
rect 30892 29996 30898 30008
rect 31481 30005 31493 30008
rect 31527 30005 31539 30039
rect 31481 29999 31539 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 8202 29792 8208 29844
rect 8260 29832 8266 29844
rect 15378 29832 15384 29844
rect 8260 29804 15384 29832
rect 8260 29792 8266 29804
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 17494 29792 17500 29844
rect 17552 29832 17558 29844
rect 20162 29832 20168 29844
rect 17552 29804 20168 29832
rect 17552 29792 17558 29804
rect 20162 29792 20168 29804
rect 20220 29792 20226 29844
rect 32677 29835 32735 29841
rect 32677 29801 32689 29835
rect 32723 29832 32735 29835
rect 32858 29832 32864 29844
rect 32723 29804 32864 29832
rect 32723 29801 32735 29804
rect 32677 29795 32735 29801
rect 32858 29792 32864 29804
rect 32916 29792 32922 29844
rect 37182 29792 37188 29844
rect 37240 29832 37246 29844
rect 37921 29835 37979 29841
rect 37921 29832 37933 29835
rect 37240 29804 37933 29832
rect 37240 29792 37246 29804
rect 37921 29801 37933 29804
rect 37967 29801 37979 29835
rect 37921 29795 37979 29801
rect 9490 29724 9496 29776
rect 9548 29764 9554 29776
rect 9861 29767 9919 29773
rect 9861 29764 9873 29767
rect 9548 29736 9873 29764
rect 9548 29724 9554 29736
rect 9861 29733 9873 29736
rect 9907 29733 9919 29767
rect 9861 29727 9919 29733
rect 11333 29767 11391 29773
rect 11333 29733 11345 29767
rect 11379 29764 11391 29767
rect 11514 29764 11520 29776
rect 11379 29736 11520 29764
rect 11379 29733 11391 29736
rect 11333 29727 11391 29733
rect 11514 29724 11520 29736
rect 11572 29724 11578 29776
rect 32309 29699 32367 29705
rect 32309 29696 32321 29699
rect 31726 29668 32321 29696
rect 10962 29588 10968 29640
rect 11020 29628 11026 29640
rect 11057 29631 11115 29637
rect 11057 29628 11069 29631
rect 11020 29600 11069 29628
rect 11020 29588 11026 29600
rect 11057 29597 11069 29600
rect 11103 29597 11115 29631
rect 11057 29591 11115 29597
rect 11149 29631 11207 29637
rect 11149 29597 11161 29631
rect 11195 29628 11207 29631
rect 11790 29628 11796 29640
rect 11195 29600 11796 29628
rect 11195 29597 11207 29600
rect 11149 29591 11207 29597
rect 11790 29588 11796 29600
rect 11848 29588 11854 29640
rect 22278 29588 22284 29640
rect 22336 29628 22342 29640
rect 25409 29631 25467 29637
rect 25409 29628 25421 29631
rect 22336 29600 25421 29628
rect 22336 29588 22342 29600
rect 25409 29597 25421 29600
rect 25455 29628 25467 29631
rect 25455 29600 26234 29628
rect 25455 29597 25467 29600
rect 25409 29591 25467 29597
rect 10045 29563 10103 29569
rect 10045 29529 10057 29563
rect 10091 29560 10103 29563
rect 10134 29560 10140 29572
rect 10091 29532 10140 29560
rect 10091 29529 10103 29532
rect 10045 29523 10103 29529
rect 10134 29520 10140 29532
rect 10192 29520 10198 29572
rect 11330 29560 11336 29572
rect 11291 29532 11336 29560
rect 11330 29520 11336 29532
rect 11388 29520 11394 29572
rect 25222 29560 25228 29572
rect 25183 29532 25228 29560
rect 25222 29520 25228 29532
rect 25280 29520 25286 29572
rect 26206 29560 26234 29600
rect 31570 29588 31576 29640
rect 31628 29628 31634 29640
rect 31726 29628 31754 29668
rect 32309 29665 32321 29668
rect 32355 29665 32367 29699
rect 32309 29659 32367 29665
rect 32398 29656 32404 29708
rect 32456 29696 32462 29708
rect 32582 29696 32588 29708
rect 32456 29668 32588 29696
rect 32456 29656 32462 29668
rect 32582 29656 32588 29668
rect 32640 29656 32646 29708
rect 31628 29600 31754 29628
rect 31628 29588 31634 29600
rect 32030 29588 32036 29640
rect 32088 29628 32094 29640
rect 32217 29631 32275 29637
rect 32217 29628 32229 29631
rect 32088 29600 32229 29628
rect 32088 29588 32094 29600
rect 32217 29597 32229 29600
rect 32263 29597 32275 29631
rect 32217 29591 32275 29597
rect 32493 29631 32551 29637
rect 32493 29597 32505 29631
rect 32539 29597 32551 29631
rect 32493 29591 32551 29597
rect 37461 29631 37519 29637
rect 37461 29597 37473 29631
rect 37507 29628 37519 29631
rect 38102 29628 38108 29640
rect 37507 29600 38108 29628
rect 37507 29597 37519 29600
rect 37461 29591 37519 29597
rect 32122 29560 32128 29572
rect 26206 29532 32128 29560
rect 32122 29520 32128 29532
rect 32180 29560 32186 29572
rect 32508 29560 32536 29591
rect 38102 29588 38108 29600
rect 38160 29588 38166 29640
rect 32180 29532 32536 29560
rect 32180 29520 32186 29532
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 9490 29248 9496 29300
rect 9548 29288 9554 29300
rect 10505 29291 10563 29297
rect 10505 29288 10517 29291
rect 9548 29260 10517 29288
rect 9548 29248 9554 29260
rect 10505 29257 10517 29260
rect 10551 29257 10563 29291
rect 10505 29251 10563 29257
rect 11517 29291 11575 29297
rect 11517 29257 11529 29291
rect 11563 29257 11575 29291
rect 22922 29288 22928 29300
rect 22883 29260 22928 29288
rect 11517 29251 11575 29257
rect 9508 29220 9536 29248
rect 11532 29220 11560 29251
rect 22922 29248 22928 29260
rect 22980 29248 22986 29300
rect 23477 29223 23535 29229
rect 23477 29220 23489 29223
rect 8680 29192 9536 29220
rect 10244 29192 11560 29220
rect 22848 29192 23489 29220
rect 8386 29112 8392 29164
rect 8444 29152 8450 29164
rect 8680 29161 8708 29192
rect 8665 29155 8723 29161
rect 8665 29152 8677 29155
rect 8444 29124 8677 29152
rect 8444 29112 8450 29124
rect 8665 29121 8677 29124
rect 8711 29121 8723 29155
rect 8665 29115 8723 29121
rect 8932 29155 8990 29161
rect 8932 29121 8944 29155
rect 8978 29152 8990 29155
rect 10244 29152 10272 29192
rect 11514 29152 11520 29164
rect 8978 29124 10272 29152
rect 11475 29124 11520 29152
rect 8978 29121 8990 29124
rect 8932 29115 8990 29121
rect 11514 29112 11520 29124
rect 11572 29112 11578 29164
rect 11606 29112 11612 29164
rect 11664 29152 11670 29164
rect 11664 29124 11709 29152
rect 11664 29112 11670 29124
rect 15378 29112 15384 29164
rect 15436 29152 15442 29164
rect 22848 29161 22876 29192
rect 23477 29189 23489 29192
rect 23523 29189 23535 29223
rect 23477 29183 23535 29189
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 15436 29124 22845 29152
rect 15436 29112 15442 29124
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 23017 29155 23075 29161
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 25222 29152 25228 29164
rect 23063 29124 25228 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 25222 29112 25228 29124
rect 25280 29112 25286 29164
rect 30282 29112 30288 29164
rect 30340 29152 30346 29164
rect 31113 29155 31171 29161
rect 31113 29152 31125 29155
rect 30340 29124 31125 29152
rect 30340 29112 30346 29124
rect 31113 29121 31125 29124
rect 31159 29121 31171 29155
rect 31113 29115 31171 29121
rect 11793 29087 11851 29093
rect 11793 29053 11805 29087
rect 11839 29084 11851 29087
rect 12253 29087 12311 29093
rect 12253 29084 12265 29087
rect 11839 29056 12265 29084
rect 11839 29053 11851 29056
rect 11793 29047 11851 29053
rect 12253 29053 12265 29056
rect 12299 29084 12311 29087
rect 13078 29084 13084 29096
rect 12299 29056 13084 29084
rect 12299 29053 12311 29056
rect 12253 29047 12311 29053
rect 13078 29044 13084 29056
rect 13136 29044 13142 29096
rect 10045 29019 10103 29025
rect 10045 28985 10057 29019
rect 10091 29016 10103 29019
rect 11330 29016 11336 29028
rect 10091 28988 11336 29016
rect 10091 28985 10103 28988
rect 10045 28979 10103 28985
rect 11330 28976 11336 28988
rect 11388 28976 11394 29028
rect 31297 29019 31355 29025
rect 31297 28985 31309 29019
rect 31343 29016 31355 29019
rect 31570 29016 31576 29028
rect 31343 28988 31576 29016
rect 31343 28985 31355 28988
rect 31297 28979 31355 28985
rect 31570 28976 31576 28988
rect 31628 28976 31634 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 6178 28744 6184 28756
rect 6139 28716 6184 28744
rect 6178 28704 6184 28716
rect 6236 28704 6242 28756
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 6972 28716 7017 28744
rect 6972 28704 6978 28716
rect 18322 28676 18328 28688
rect 18283 28648 18328 28676
rect 18322 28636 18328 28648
rect 18380 28636 18386 28688
rect 6178 28500 6184 28552
rect 6236 28540 6242 28552
rect 6730 28540 6736 28552
rect 6236 28512 6736 28540
rect 6236 28500 6242 28512
rect 6730 28500 6736 28512
rect 6788 28500 6794 28552
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 18472 28512 18517 28540
rect 18472 28500 18478 28512
rect 18141 28475 18199 28481
rect 18141 28441 18153 28475
rect 18187 28441 18199 28475
rect 18141 28435 18199 28441
rect 17586 28404 17592 28416
rect 17547 28376 17592 28404
rect 17586 28364 17592 28376
rect 17644 28404 17650 28416
rect 18156 28404 18184 28435
rect 28994 28432 29000 28484
rect 29052 28472 29058 28484
rect 30653 28475 30711 28481
rect 30653 28472 30665 28475
rect 29052 28444 30665 28472
rect 29052 28432 29058 28444
rect 30653 28441 30665 28444
rect 30699 28441 30711 28475
rect 30653 28435 30711 28441
rect 18414 28404 18420 28416
rect 17644 28376 18184 28404
rect 18375 28376 18420 28404
rect 17644 28364 17650 28376
rect 18414 28364 18420 28376
rect 18472 28364 18478 28416
rect 26418 28364 26424 28416
rect 26476 28404 26482 28416
rect 26513 28407 26571 28413
rect 26513 28404 26525 28407
rect 26476 28376 26525 28404
rect 26476 28364 26482 28376
rect 26513 28373 26525 28376
rect 26559 28373 26571 28407
rect 30742 28404 30748 28416
rect 30703 28376 30748 28404
rect 26513 28367 26571 28373
rect 30742 28364 30748 28376
rect 30800 28364 30806 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 28537 28203 28595 28209
rect 28537 28169 28549 28203
rect 28583 28200 28595 28203
rect 30282 28200 30288 28212
rect 28583 28172 30288 28200
rect 28583 28169 28595 28172
rect 28537 28163 28595 28169
rect 30282 28160 30288 28172
rect 30340 28160 30346 28212
rect 31570 28160 31576 28212
rect 31628 28200 31634 28212
rect 32217 28203 32275 28209
rect 32217 28200 32229 28203
rect 31628 28172 32229 28200
rect 31628 28160 31634 28172
rect 32217 28169 32229 28172
rect 32263 28169 32275 28203
rect 32217 28163 32275 28169
rect 28997 28135 29055 28141
rect 28997 28132 29009 28135
rect 27172 28104 29009 28132
rect 27172 28076 27200 28104
rect 28997 28101 29009 28104
rect 29043 28132 29055 28135
rect 30742 28132 30748 28144
rect 29043 28104 30748 28132
rect 29043 28101 29055 28104
rect 28997 28095 29055 28101
rect 30742 28092 30748 28104
rect 30800 28132 30806 28144
rect 34422 28132 34428 28144
rect 30800 28104 34428 28132
rect 30800 28092 30806 28104
rect 34422 28092 34428 28104
rect 34480 28092 34486 28144
rect 25222 28024 25228 28076
rect 25280 28064 25286 28076
rect 26142 28064 26148 28076
rect 25280 28036 26148 28064
rect 25280 28024 25286 28036
rect 26142 28024 26148 28036
rect 26200 28024 26206 28076
rect 26234 28024 26240 28076
rect 26292 28064 26298 28076
rect 26418 28064 26424 28076
rect 26292 28036 26337 28064
rect 26379 28036 26424 28064
rect 26292 28024 26298 28036
rect 26418 28024 26424 28036
rect 26476 28024 26482 28076
rect 27154 28064 27160 28076
rect 27115 28036 27160 28064
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27430 28073 27436 28076
rect 27424 28027 27436 28073
rect 27488 28064 27494 28076
rect 27488 28036 27524 28064
rect 27430 28024 27436 28027
rect 27488 28024 27494 28036
rect 31754 28024 31760 28076
rect 31812 28064 31818 28076
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31812 28036 32137 28064
rect 31812 28024 31818 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 32401 28067 32459 28073
rect 32401 28033 32413 28067
rect 32447 28064 32459 28067
rect 32582 28064 32588 28076
rect 32447 28036 32588 28064
rect 32447 28033 32459 28036
rect 32401 28027 32459 28033
rect 32582 28024 32588 28036
rect 32640 28024 32646 28076
rect 37461 28067 37519 28073
rect 37461 28033 37473 28067
rect 37507 28064 37519 28067
rect 38102 28064 38108 28076
rect 37507 28036 38108 28064
rect 37507 28033 37519 28036
rect 37461 28027 37519 28033
rect 38102 28024 38108 28036
rect 38160 28024 38166 28076
rect 26421 27863 26479 27869
rect 26421 27829 26433 27863
rect 26467 27860 26479 27863
rect 27062 27860 27068 27872
rect 26467 27832 27068 27860
rect 26467 27829 26479 27832
rect 26421 27823 26479 27829
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 32398 27860 32404 27872
rect 32359 27832 32404 27860
rect 32398 27820 32404 27832
rect 32456 27820 32462 27872
rect 34790 27820 34796 27872
rect 34848 27860 34854 27872
rect 37921 27863 37979 27869
rect 37921 27860 37933 27863
rect 34848 27832 37933 27860
rect 34848 27820 34854 27832
rect 37921 27829 37933 27832
rect 37967 27829 37979 27863
rect 37921 27823 37979 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 27341 27659 27399 27665
rect 27341 27625 27353 27659
rect 27387 27656 27399 27659
rect 27430 27656 27436 27668
rect 27387 27628 27436 27656
rect 27387 27625 27399 27628
rect 27341 27619 27399 27625
rect 27430 27616 27436 27628
rect 27488 27616 27494 27668
rect 31754 27656 31760 27668
rect 31588 27628 31760 27656
rect 4798 27588 4804 27600
rect 4759 27560 4804 27588
rect 4798 27548 4804 27560
rect 4856 27548 4862 27600
rect 5997 27591 6055 27597
rect 5997 27557 6009 27591
rect 6043 27588 6055 27591
rect 6914 27588 6920 27600
rect 6043 27560 6920 27588
rect 6043 27557 6055 27560
rect 5997 27551 6055 27557
rect 5626 27520 5632 27532
rect 4632 27492 5632 27520
rect 4632 27461 4660 27492
rect 5626 27480 5632 27492
rect 5684 27480 5690 27532
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27421 4583 27455
rect 4525 27415 4583 27421
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27421 4675 27455
rect 4617 27415 4675 27421
rect 4540 27384 4568 27415
rect 4798 27412 4804 27464
rect 4856 27452 4862 27464
rect 5261 27455 5319 27461
rect 5261 27452 5273 27455
rect 4856 27424 5273 27452
rect 4856 27412 4862 27424
rect 5261 27421 5273 27424
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 5445 27455 5503 27461
rect 5445 27421 5457 27455
rect 5491 27452 5503 27455
rect 6012 27452 6040 27551
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 18690 27588 18696 27600
rect 18651 27560 18696 27588
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 26142 27548 26148 27600
rect 26200 27588 26206 27600
rect 26200 27548 26234 27588
rect 26206 27520 26234 27548
rect 26973 27523 27031 27529
rect 26973 27520 26985 27523
rect 26206 27492 26985 27520
rect 26973 27489 26985 27492
rect 27019 27520 27031 27523
rect 31588 27520 31616 27628
rect 31754 27616 31760 27628
rect 31812 27616 31818 27668
rect 32582 27588 32588 27600
rect 31680 27560 32588 27588
rect 31680 27529 31708 27560
rect 32582 27548 32588 27560
rect 32640 27548 32646 27600
rect 34422 27548 34428 27600
rect 34480 27588 34486 27600
rect 35621 27591 35679 27597
rect 35621 27588 35633 27591
rect 34480 27560 35633 27588
rect 34480 27548 34486 27560
rect 35621 27557 35633 27560
rect 35667 27557 35679 27591
rect 37550 27588 37556 27600
rect 37511 27560 37556 27588
rect 35621 27551 35679 27557
rect 27019 27492 31616 27520
rect 31665 27523 31723 27529
rect 27019 27489 27031 27492
rect 26973 27483 27031 27489
rect 31665 27489 31677 27523
rect 31711 27489 31723 27523
rect 31665 27483 31723 27489
rect 31754 27480 31760 27532
rect 31812 27520 31818 27532
rect 31941 27523 31999 27529
rect 31812 27492 31857 27520
rect 31812 27480 31818 27492
rect 31941 27489 31953 27523
rect 31987 27520 31999 27523
rect 35636 27520 35664 27551
rect 37550 27548 37556 27560
rect 37608 27548 37614 27600
rect 35710 27520 35716 27532
rect 31987 27492 32628 27520
rect 35623 27492 35716 27520
rect 31987 27489 31999 27492
rect 31941 27483 31999 27489
rect 17313 27455 17371 27461
rect 17313 27452 17325 27455
rect 5491 27424 6040 27452
rect 16776 27424 17325 27452
rect 5491 27421 5503 27424
rect 5445 27415 5503 27421
rect 4890 27384 4896 27396
rect 4540 27356 4896 27384
rect 4890 27344 4896 27356
rect 4948 27344 4954 27396
rect 5350 27316 5356 27328
rect 5311 27288 5356 27316
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 15470 27276 15476 27328
rect 15528 27316 15534 27328
rect 16776 27325 16804 27424
rect 17313 27421 17325 27424
rect 17359 27421 17371 27455
rect 17313 27415 17371 27421
rect 17580 27455 17638 27461
rect 17580 27421 17592 27455
rect 17626 27452 17638 27455
rect 18414 27452 18420 27464
rect 17626 27424 18420 27452
rect 17626 27421 17638 27424
rect 17580 27415 17638 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 26234 27412 26240 27464
rect 26292 27452 26298 27464
rect 26881 27455 26939 27461
rect 26881 27452 26893 27455
rect 26292 27424 26893 27452
rect 26292 27412 26298 27424
rect 26881 27421 26893 27424
rect 26927 27421 26939 27455
rect 26881 27415 26939 27421
rect 26896 27384 26924 27415
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27157 27455 27215 27461
rect 27157 27452 27169 27455
rect 27120 27424 27169 27452
rect 27120 27412 27126 27424
rect 27157 27421 27169 27424
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 30834 27412 30840 27464
rect 30892 27452 30898 27464
rect 31481 27455 31539 27461
rect 31481 27452 31493 27455
rect 30892 27424 31493 27452
rect 30892 27412 30898 27424
rect 31481 27421 31493 27424
rect 31527 27421 31539 27455
rect 31481 27415 31539 27421
rect 31570 27412 31576 27464
rect 31628 27452 31634 27464
rect 32398 27452 32404 27464
rect 31628 27424 31721 27452
rect 32359 27424 32404 27452
rect 31628 27412 31634 27424
rect 32398 27412 32404 27424
rect 32456 27412 32462 27464
rect 32600 27461 32628 27492
rect 35710 27480 35716 27492
rect 35768 27520 35774 27532
rect 36173 27523 36231 27529
rect 36173 27520 36185 27523
rect 35768 27492 36185 27520
rect 35768 27480 35774 27492
rect 36173 27489 36185 27492
rect 36219 27489 36231 27523
rect 36173 27483 36231 27489
rect 32585 27455 32643 27461
rect 32585 27421 32597 27455
rect 32631 27421 32643 27455
rect 32585 27415 32643 27421
rect 31588 27384 31616 27412
rect 26896 27356 31616 27384
rect 36262 27344 36268 27396
rect 36320 27384 36326 27396
rect 36418 27387 36476 27393
rect 36418 27384 36430 27387
rect 36320 27356 36430 27384
rect 36320 27344 36326 27356
rect 36418 27353 36430 27356
rect 36464 27353 36476 27387
rect 36418 27347 36476 27353
rect 16761 27319 16819 27325
rect 16761 27316 16773 27319
rect 15528 27288 16773 27316
rect 15528 27276 15534 27288
rect 16761 27285 16773 27288
rect 16807 27285 16819 27319
rect 30834 27316 30840 27328
rect 30795 27288 30840 27316
rect 16761 27279 16819 27285
rect 30834 27276 30840 27288
rect 30892 27276 30898 27328
rect 32490 27316 32496 27328
rect 32451 27288 32496 27316
rect 32490 27276 32496 27288
rect 32548 27276 32554 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 33873 27115 33931 27121
rect 33873 27081 33885 27115
rect 33919 27112 33931 27115
rect 34422 27112 34428 27124
rect 33919 27084 34428 27112
rect 33919 27081 33931 27084
rect 33873 27075 33931 27081
rect 34422 27072 34428 27084
rect 34480 27072 34486 27124
rect 32490 27004 32496 27056
rect 32548 27044 32554 27056
rect 35446 27047 35504 27053
rect 35446 27044 35458 27047
rect 32548 27016 35458 27044
rect 32548 27004 32554 27016
rect 35446 27013 35458 27016
rect 35492 27044 35504 27047
rect 36262 27044 36268 27056
rect 35492 27016 36268 27044
rect 35492 27013 35504 27016
rect 35446 27007 35504 27013
rect 36262 27004 36268 27016
rect 36320 27004 36326 27056
rect 15013 26979 15071 26985
rect 15013 26945 15025 26979
rect 15059 26976 15071 26979
rect 15838 26976 15844 26988
rect 15059 26948 15844 26976
rect 15059 26945 15071 26948
rect 15013 26939 15071 26945
rect 15838 26936 15844 26948
rect 15896 26936 15902 26988
rect 35710 26976 35716 26988
rect 35671 26948 35716 26976
rect 35710 26936 35716 26948
rect 35768 26936 35774 26988
rect 16574 26868 16580 26920
rect 16632 26908 16638 26920
rect 16758 26908 16764 26920
rect 16632 26880 16764 26908
rect 16632 26868 16638 26880
rect 16758 26868 16764 26880
rect 16816 26868 16822 26920
rect 17586 26840 17592 26852
rect 15212 26812 17592 26840
rect 13078 26732 13084 26784
rect 13136 26772 13142 26784
rect 15212 26781 15240 26812
rect 17586 26800 17592 26812
rect 17644 26800 17650 26852
rect 32582 26800 32588 26852
rect 32640 26840 32646 26852
rect 34333 26843 34391 26849
rect 34333 26840 34345 26843
rect 32640 26812 34345 26840
rect 32640 26800 32646 26812
rect 34333 26809 34345 26812
rect 34379 26809 34391 26843
rect 34333 26803 34391 26809
rect 15197 26775 15255 26781
rect 15197 26772 15209 26775
rect 13136 26744 15209 26772
rect 13136 26732 13142 26744
rect 15197 26741 15209 26744
rect 15243 26741 15255 26775
rect 15838 26772 15844 26784
rect 15799 26744 15844 26772
rect 15197 26735 15255 26741
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 4157 26571 4215 26577
rect 4157 26537 4169 26571
rect 4203 26568 4215 26571
rect 5626 26568 5632 26580
rect 4203 26540 5632 26568
rect 4203 26537 4215 26540
rect 4157 26531 4215 26537
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 15838 26528 15844 26580
rect 15896 26568 15902 26580
rect 30834 26568 30840 26580
rect 15896 26540 30840 26568
rect 15896 26528 15902 26540
rect 30834 26528 30840 26540
rect 30892 26528 30898 26580
rect 5350 26432 5356 26444
rect 3988 26404 5356 26432
rect 3988 26373 4016 26404
rect 5350 26392 5356 26404
rect 5408 26392 5414 26444
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4246 26324 4252 26376
rect 4304 26364 4310 26376
rect 4890 26364 4896 26376
rect 4304 26336 4896 26364
rect 4304 26324 4310 26336
rect 4890 26324 4896 26336
rect 4948 26324 4954 26376
rect 3786 26228 3792 26240
rect 3747 26200 3792 26228
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 3697 26027 3755 26033
rect 3697 25993 3709 26027
rect 3743 26024 3755 26027
rect 4154 26024 4160 26036
rect 3743 25996 4160 26024
rect 3743 25993 3755 25996
rect 3697 25987 3755 25993
rect 4154 25984 4160 25996
rect 4212 25984 4218 26036
rect 4249 26027 4307 26033
rect 4249 25993 4261 26027
rect 4295 26024 4307 26027
rect 8386 26024 8392 26036
rect 4295 25996 8392 26024
rect 4295 25993 4307 25996
rect 4249 25987 4307 25993
rect 4264 25956 4292 25987
rect 8386 25984 8392 25996
rect 8444 25984 8450 26036
rect 26418 25984 26424 26036
rect 26476 26024 26482 26036
rect 27065 26027 27123 26033
rect 27065 26024 27077 26027
rect 26476 25996 27077 26024
rect 26476 25984 26482 25996
rect 27065 25993 27077 25996
rect 27111 25993 27123 26027
rect 30834 26024 30840 26036
rect 30795 25996 30840 26024
rect 27065 25987 27123 25993
rect 30834 25984 30840 25996
rect 30892 25984 30898 26036
rect 23753 25959 23811 25965
rect 23753 25956 23765 25959
rect 2332 25928 4292 25956
rect 21836 25928 23765 25956
rect 2332 25897 2360 25928
rect 2317 25891 2375 25897
rect 2317 25857 2329 25891
rect 2363 25857 2375 25891
rect 2317 25851 2375 25857
rect 2584 25891 2642 25897
rect 2584 25857 2596 25891
rect 2630 25888 2642 25891
rect 3786 25888 3792 25900
rect 2630 25860 3792 25888
rect 2630 25857 2642 25860
rect 2584 25851 2642 25857
rect 3786 25848 3792 25860
rect 3844 25848 3850 25900
rect 21836 25897 21864 25928
rect 23753 25925 23765 25928
rect 23799 25956 23811 25959
rect 27154 25956 27160 25968
rect 23799 25928 27160 25956
rect 23799 25925 23811 25928
rect 23753 25919 23811 25925
rect 27154 25916 27160 25928
rect 27212 25916 27218 25968
rect 30193 25959 30251 25965
rect 30193 25956 30205 25959
rect 27264 25928 30205 25956
rect 22094 25897 22100 25900
rect 21821 25891 21879 25897
rect 21821 25857 21833 25891
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 22088 25851 22100 25897
rect 22152 25888 22158 25900
rect 27264 25897 27292 25928
rect 30193 25925 30205 25928
rect 30239 25956 30251 25959
rect 30742 25956 30748 25968
rect 30239 25928 30748 25956
rect 30239 25925 30251 25928
rect 30193 25919 30251 25925
rect 30742 25916 30748 25928
rect 30800 25916 30806 25968
rect 26421 25891 26479 25897
rect 26421 25888 26433 25891
rect 22152 25860 22188 25888
rect 26206 25860 26433 25888
rect 22094 25848 22100 25851
rect 22152 25848 22158 25860
rect 8386 25712 8392 25764
rect 8444 25752 8450 25764
rect 8481 25755 8539 25761
rect 8481 25752 8493 25755
rect 8444 25724 8493 25752
rect 8444 25712 8450 25724
rect 8481 25721 8493 25724
rect 8527 25752 8539 25755
rect 13909 25755 13967 25761
rect 13909 25752 13921 25755
rect 8527 25724 13921 25752
rect 8527 25721 8539 25724
rect 8481 25715 8539 25721
rect 13909 25721 13921 25724
rect 13955 25752 13967 25755
rect 15470 25752 15476 25764
rect 13955 25724 15476 25752
rect 13955 25721 13967 25724
rect 13909 25715 13967 25721
rect 15470 25712 15476 25724
rect 15528 25712 15534 25764
rect 26206 25752 26234 25860
rect 26421 25857 26433 25860
rect 26467 25888 26479 25891
rect 27249 25891 27307 25897
rect 27249 25888 27261 25891
rect 26467 25860 27261 25888
rect 26467 25857 26479 25860
rect 26421 25851 26479 25857
rect 27249 25857 27261 25860
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 38102 25752 38108 25764
rect 22756 25724 26234 25752
rect 38063 25724 38108 25752
rect 14458 25644 14464 25696
rect 14516 25684 14522 25696
rect 22756 25684 22784 25724
rect 38102 25712 38108 25724
rect 38160 25712 38166 25764
rect 14516 25656 22784 25684
rect 14516 25644 14522 25656
rect 23106 25644 23112 25696
rect 23164 25684 23170 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 23164 25656 23213 25684
rect 23164 25644 23170 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 13078 25480 13084 25492
rect 9876 25452 11652 25480
rect 13039 25452 13084 25480
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 8386 25276 8392 25288
rect 6963 25248 8392 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 9876 25285 9904 25452
rect 11514 25412 11520 25424
rect 10152 25384 11520 25412
rect 10152 25285 10180 25384
rect 11514 25372 11520 25384
rect 11572 25372 11578 25424
rect 11624 25412 11652 25452
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 22005 25483 22063 25489
rect 22005 25449 22017 25483
rect 22051 25480 22063 25483
rect 22094 25480 22100 25492
rect 22051 25452 22100 25480
rect 22051 25449 22063 25452
rect 22005 25443 22063 25449
rect 22094 25440 22100 25452
rect 22152 25440 22158 25492
rect 22373 25483 22431 25489
rect 22373 25449 22385 25483
rect 22419 25480 22431 25483
rect 22419 25452 23244 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 14458 25412 14464 25424
rect 11624 25384 14464 25412
rect 14458 25372 14464 25384
rect 14516 25372 14522 25424
rect 22925 25415 22983 25421
rect 22925 25381 22937 25415
rect 22971 25381 22983 25415
rect 22925 25375 22983 25381
rect 15470 25344 15476 25356
rect 15431 25316 15476 25344
rect 15470 25304 15476 25316
rect 15528 25304 15534 25356
rect 22940 25344 22968 25375
rect 22204 25316 22968 25344
rect 22204 25285 22232 25316
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25276 9275 25279
rect 9861 25279 9919 25285
rect 9861 25276 9873 25279
rect 9263 25248 9873 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 9861 25245 9873 25248
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25245 10379 25279
rect 10321 25239 10379 25245
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 22465 25279 22523 25285
rect 22465 25245 22477 25279
rect 22511 25276 22523 25279
rect 23106 25276 23112 25288
rect 22511 25248 23112 25276
rect 22511 25245 22523 25248
rect 22465 25239 22523 25245
rect 7184 25211 7242 25217
rect 7184 25177 7196 25211
rect 7230 25208 7242 25211
rect 7926 25208 7932 25220
rect 7230 25180 7932 25208
rect 7230 25177 7242 25180
rect 7184 25171 7242 25177
rect 7926 25168 7932 25180
rect 7984 25168 7990 25220
rect 9232 25208 9260 25239
rect 10336 25208 10364 25239
rect 10962 25208 10968 25220
rect 8220 25180 9260 25208
rect 9508 25180 10968 25208
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 8220 25140 8248 25180
rect 6788 25112 8248 25140
rect 8297 25143 8355 25149
rect 6788 25100 6794 25112
rect 8297 25109 8309 25143
rect 8343 25140 8355 25143
rect 9508 25140 9536 25180
rect 10962 25168 10968 25180
rect 11020 25168 11026 25220
rect 12986 25168 12992 25220
rect 13044 25208 13050 25220
rect 15206 25211 15264 25217
rect 15206 25208 15218 25211
rect 13044 25180 15218 25208
rect 13044 25168 13050 25180
rect 15206 25177 15218 25180
rect 15252 25177 15264 25211
rect 15206 25171 15264 25177
rect 22002 25168 22008 25220
rect 22060 25208 22066 25220
rect 22480 25208 22508 25239
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23216 25285 23244 25452
rect 30926 25440 30932 25492
rect 30984 25480 30990 25492
rect 31021 25483 31079 25489
rect 31021 25480 31033 25483
rect 30984 25452 31033 25480
rect 30984 25440 30990 25452
rect 31021 25449 31033 25452
rect 31067 25449 31079 25483
rect 31021 25443 31079 25449
rect 31386 25304 31392 25356
rect 31444 25344 31450 25356
rect 31573 25347 31631 25353
rect 31573 25344 31585 25347
rect 31444 25316 31585 25344
rect 31444 25304 31450 25316
rect 31573 25313 31585 25316
rect 31619 25313 31631 25347
rect 31573 25307 31631 25313
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23290 25276 23296 25288
rect 23247 25248 23296 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23290 25236 23296 25248
rect 23348 25236 23354 25288
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25276 31539 25279
rect 34790 25276 34796 25288
rect 31527 25248 34796 25276
rect 31527 25245 31539 25248
rect 31481 25239 31539 25245
rect 34790 25236 34796 25248
rect 34848 25236 34854 25288
rect 22060 25180 22508 25208
rect 22925 25211 22983 25217
rect 22060 25168 22066 25180
rect 22925 25177 22937 25211
rect 22971 25177 22983 25211
rect 22925 25171 22983 25177
rect 28813 25211 28871 25217
rect 28813 25177 28825 25211
rect 28859 25177 28871 25211
rect 28994 25208 29000 25220
rect 28955 25180 29000 25208
rect 28813 25171 28871 25177
rect 9674 25140 9680 25152
rect 8343 25112 9536 25140
rect 9635 25112 9680 25140
rect 8343 25109 8355 25112
rect 8297 25103 8355 25109
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 14090 25140 14096 25152
rect 14051 25112 14096 25140
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 22940 25140 22968 25171
rect 23661 25143 23719 25149
rect 23661 25140 23673 25143
rect 20036 25112 23673 25140
rect 20036 25100 20042 25112
rect 23661 25109 23673 25112
rect 23707 25140 23719 25143
rect 25682 25140 25688 25152
rect 23707 25112 25688 25140
rect 23707 25109 23719 25112
rect 23661 25103 23719 25109
rect 25682 25100 25688 25112
rect 25740 25140 25746 25152
rect 26418 25140 26424 25152
rect 25740 25112 26424 25140
rect 25740 25100 25746 25112
rect 26418 25100 26424 25112
rect 26476 25100 26482 25152
rect 28166 25140 28172 25152
rect 28127 25112 28172 25140
rect 28166 25100 28172 25112
rect 28224 25140 28230 25152
rect 28828 25140 28856 25171
rect 28994 25168 29000 25180
rect 29052 25168 29058 25220
rect 31389 25211 31447 25217
rect 31389 25177 31401 25211
rect 31435 25208 31447 25211
rect 31570 25208 31576 25220
rect 31435 25180 31576 25208
rect 31435 25177 31447 25180
rect 31389 25171 31447 25177
rect 31570 25168 31576 25180
rect 31628 25208 31634 25220
rect 32217 25211 32275 25217
rect 32217 25208 32229 25211
rect 31628 25180 32229 25208
rect 31628 25168 31634 25180
rect 32217 25177 32229 25180
rect 32263 25177 32275 25211
rect 32217 25171 32275 25177
rect 28224 25112 28856 25140
rect 28224 25100 28230 25112
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7926 24936 7932 24948
rect 7887 24908 7932 24936
rect 7926 24896 7932 24908
rect 7984 24896 7990 24948
rect 11514 24896 11520 24948
rect 11572 24936 11578 24948
rect 12986 24936 12992 24948
rect 11572 24908 12388 24936
rect 12947 24908 12992 24936
rect 11572 24896 11578 24908
rect 12360 24880 12388 24908
rect 12986 24896 12992 24908
rect 13044 24896 13050 24948
rect 9674 24828 9680 24880
rect 9732 24828 9738 24880
rect 11348 24840 11652 24868
rect 8113 24803 8171 24809
rect 8113 24769 8125 24803
rect 8159 24800 8171 24803
rect 9309 24803 9367 24809
rect 9309 24800 9321 24803
rect 8159 24772 9321 24800
rect 8159 24769 8171 24772
rect 8113 24763 8171 24769
rect 9309 24769 9321 24772
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24800 9551 24803
rect 9692 24800 9720 24828
rect 9539 24772 9720 24800
rect 10321 24803 10379 24809
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 10367 24772 10916 24800
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 10888 24741 10916 24772
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 11348 24800 11376 24840
rect 11514 24800 11520 24812
rect 11020 24772 11376 24800
rect 11475 24772 11520 24800
rect 11020 24760 11026 24772
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 11624 24800 11652 24840
rect 12342 24828 12348 24880
rect 12400 24868 12406 24880
rect 12400 24840 12664 24868
rect 12400 24828 12406 24840
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11624 24772 11713 24800
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 12526 24800 12532 24812
rect 12487 24772 12532 24800
rect 11701 24763 11759 24769
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 12636 24809 12664 24840
rect 12621 24803 12679 24809
rect 12621 24769 12633 24803
rect 12667 24769 12679 24803
rect 12621 24763 12679 24769
rect 12713 24803 12771 24809
rect 12713 24769 12725 24803
rect 12759 24769 12771 24803
rect 12713 24763 12771 24769
rect 12897 24803 12955 24809
rect 12897 24769 12909 24803
rect 12943 24769 12955 24803
rect 12897 24763 12955 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24800 13047 24803
rect 13078 24800 13084 24812
rect 13035 24772 13084 24800
rect 13035 24769 13047 24772
rect 12989 24763 13047 24769
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24701 9735 24735
rect 9677 24695 9735 24701
rect 10873 24735 10931 24741
rect 10873 24701 10885 24735
rect 10919 24732 10931 24735
rect 12434 24732 12440 24744
rect 10919 24704 12440 24732
rect 10919 24701 10931 24704
rect 10873 24695 10931 24701
rect 9692 24596 9720 24695
rect 12434 24692 12440 24704
rect 12492 24692 12498 24744
rect 10134 24664 10140 24676
rect 10095 24636 10140 24664
rect 10134 24624 10140 24636
rect 10192 24624 10198 24676
rect 11609 24599 11667 24605
rect 11609 24596 11621 24599
rect 9692 24568 11621 24596
rect 11609 24565 11621 24568
rect 11655 24596 11667 24599
rect 12728 24596 12756 24763
rect 12912 24732 12940 24763
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 14090 24800 14096 24812
rect 13679 24772 14096 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 20898 24760 20904 24812
rect 20956 24800 20962 24812
rect 28166 24800 28172 24812
rect 20956 24772 28172 24800
rect 20956 24760 20962 24772
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 12912 24704 13553 24732
rect 13541 24701 13553 24704
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 11655 24568 12756 24596
rect 11655 24565 11667 24568
rect 11609 24559 11667 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 20898 24392 20904 24404
rect 12492 24364 20904 24392
rect 12492 24352 12498 24364
rect 20898 24352 20904 24364
rect 20956 24352 20962 24404
rect 25682 24392 25688 24404
rect 25643 24364 25688 24392
rect 25682 24352 25688 24364
rect 25740 24352 25746 24404
rect 8846 24284 8852 24336
rect 8904 24324 8910 24336
rect 30377 24327 30435 24333
rect 30377 24324 30389 24327
rect 8904 24296 30389 24324
rect 8904 24284 8910 24296
rect 30377 24293 30389 24296
rect 30423 24293 30435 24327
rect 30377 24287 30435 24293
rect 8018 24216 8024 24268
rect 8076 24256 8082 24268
rect 29549 24259 29607 24265
rect 29549 24256 29561 24259
rect 8076 24228 29561 24256
rect 8076 24216 8082 24228
rect 29549 24225 29561 24228
rect 29595 24225 29607 24259
rect 29549 24219 29607 24225
rect 10962 24148 10968 24200
rect 11020 24188 11026 24200
rect 12621 24191 12679 24197
rect 12621 24188 12633 24191
rect 11020 24160 12633 24188
rect 11020 24148 11026 24160
rect 12621 24157 12633 24160
rect 12667 24157 12679 24191
rect 12621 24151 12679 24157
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 14090 24188 14096 24200
rect 12851 24160 14096 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 23348 24160 25053 24188
rect 23348 24148 23354 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 25225 24191 25283 24197
rect 25225 24157 25237 24191
rect 25271 24188 25283 24191
rect 25682 24188 25688 24200
rect 25271 24160 25688 24188
rect 25271 24157 25283 24160
rect 25225 24151 25283 24157
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24188 29791 24191
rect 30561 24191 30619 24197
rect 30561 24188 30573 24191
rect 29779 24160 30573 24188
rect 29779 24157 29791 24160
rect 29733 24151 29791 24157
rect 30561 24157 30573 24160
rect 30607 24188 30619 24191
rect 31386 24188 31392 24200
rect 30607 24160 31392 24188
rect 30607 24157 30619 24160
rect 30561 24151 30619 24157
rect 31386 24148 31392 24160
rect 31444 24148 31450 24200
rect 19426 24080 19432 24132
rect 19484 24120 19490 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 19484 24092 19625 24120
rect 19484 24080 19490 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 29917 24123 29975 24129
rect 29917 24089 29929 24123
rect 29963 24120 29975 24123
rect 30098 24120 30104 24132
rect 29963 24092 30104 24120
rect 29963 24089 29975 24092
rect 29917 24083 29975 24089
rect 30098 24080 30104 24092
rect 30156 24080 30162 24132
rect 30745 24123 30803 24129
rect 30745 24089 30757 24123
rect 30791 24120 30803 24123
rect 30834 24120 30840 24132
rect 30791 24092 30840 24120
rect 30791 24089 30803 24092
rect 30745 24083 30803 24089
rect 30834 24080 30840 24092
rect 30892 24120 30898 24132
rect 31205 24123 31263 24129
rect 31205 24120 31217 24123
rect 30892 24092 31217 24120
rect 30892 24080 30898 24092
rect 31205 24089 31217 24092
rect 31251 24089 31263 24123
rect 31205 24083 31263 24089
rect 37369 24123 37427 24129
rect 37369 24089 37381 24123
rect 37415 24120 37427 24123
rect 38010 24120 38016 24132
rect 37415 24092 38016 24120
rect 37415 24089 37427 24092
rect 37369 24083 37427 24089
rect 38010 24080 38016 24092
rect 38068 24080 38074 24132
rect 12437 24055 12495 24061
rect 12437 24021 12449 24055
rect 12483 24052 12495 24055
rect 12526 24052 12532 24064
rect 12483 24024 12532 24052
rect 12483 24021 12495 24024
rect 12437 24015 12495 24021
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 25130 24052 25136 24064
rect 25091 24024 25136 24052
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 37918 24052 37924 24064
rect 37879 24024 37924 24052
rect 37918 24012 37924 24024
rect 37976 24012 37982 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 37277 23851 37335 23857
rect 37277 23817 37289 23851
rect 37323 23848 37335 23851
rect 37458 23848 37464 23860
rect 37323 23820 37464 23848
rect 37323 23817 37335 23820
rect 37277 23811 37335 23817
rect 37458 23808 37464 23820
rect 37516 23808 37522 23860
rect 37550 23808 37556 23860
rect 37608 23848 37614 23860
rect 37737 23851 37795 23857
rect 37737 23848 37749 23851
rect 37608 23820 37749 23848
rect 37608 23808 37614 23820
rect 37737 23817 37749 23820
rect 37783 23817 37795 23851
rect 37737 23811 37795 23817
rect 10594 23740 10600 23792
rect 10652 23780 10658 23792
rect 31205 23783 31263 23789
rect 31205 23780 31217 23783
rect 10652 23752 31217 23780
rect 10652 23740 10658 23752
rect 31205 23749 31217 23752
rect 31251 23749 31263 23783
rect 31386 23780 31392 23792
rect 31347 23752 31392 23780
rect 31205 23743 31263 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 17580 23715 17638 23721
rect 17580 23681 17592 23715
rect 17626 23712 17638 23715
rect 18046 23712 18052 23724
rect 17626 23684 18052 23712
rect 17626 23681 17638 23684
rect 17580 23675 17638 23681
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23712 31631 23715
rect 37642 23712 37648 23724
rect 31619 23684 31754 23712
rect 37603 23684 37648 23712
rect 31619 23681 31631 23684
rect 31573 23675 31631 23681
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 16776 23616 17325 23644
rect 16776 23520 16804 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 18693 23579 18751 23585
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 20622 23576 20628 23588
rect 18739 23548 20628 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 16758 23508 16764 23520
rect 16719 23480 16764 23508
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 19426 23508 19432 23520
rect 19387 23480 19432 23508
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 30098 23508 30104 23520
rect 30059 23480 30104 23508
rect 30098 23468 30104 23480
rect 30156 23468 30162 23520
rect 31726 23508 31754 23684
rect 37642 23672 37648 23684
rect 37700 23672 37706 23724
rect 35894 23604 35900 23656
rect 35952 23644 35958 23656
rect 37829 23647 37887 23653
rect 37829 23644 37841 23647
rect 35952 23616 37841 23644
rect 35952 23604 35958 23616
rect 37829 23613 37841 23616
rect 37875 23613 37887 23647
rect 37829 23607 37887 23613
rect 32217 23511 32275 23517
rect 32217 23508 32229 23511
rect 31726 23480 32229 23508
rect 32217 23477 32229 23480
rect 32263 23508 32275 23511
rect 32306 23508 32312 23520
rect 32263 23480 32312 23508
rect 32263 23477 32275 23480
rect 32217 23471 32275 23477
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 17313 23307 17371 23313
rect 17313 23273 17325 23307
rect 17359 23304 17371 23307
rect 17586 23304 17592 23316
rect 17359 23276 17592 23304
rect 17359 23273 17371 23276
rect 17313 23267 17371 23273
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 18046 23304 18052 23316
rect 18007 23276 18052 23304
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 17604 23168 17632 23264
rect 20993 23239 21051 23245
rect 20993 23205 21005 23239
rect 21039 23205 21051 23239
rect 20993 23199 21051 23205
rect 17678 23168 17684 23180
rect 17591 23140 17684 23168
rect 17678 23128 17684 23140
rect 17736 23168 17742 23180
rect 17773 23171 17831 23177
rect 17773 23168 17785 23171
rect 17736 23140 17785 23168
rect 17736 23128 17742 23140
rect 17773 23137 17785 23140
rect 17819 23137 17831 23171
rect 17773 23131 17831 23137
rect 17954 23100 17960 23112
rect 17915 23072 17960 23100
rect 17954 23060 17960 23072
rect 18012 23060 18018 23112
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 21008 23100 21036 23199
rect 31386 23128 31392 23180
rect 31444 23168 31450 23180
rect 32493 23171 32551 23177
rect 32493 23168 32505 23171
rect 31444 23140 32505 23168
rect 31444 23128 31450 23140
rect 32493 23137 32505 23140
rect 32539 23137 32551 23171
rect 32493 23131 32551 23137
rect 21266 23100 21272 23112
rect 18095 23072 21036 23100
rect 21227 23072 21272 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23100 25835 23103
rect 27617 23103 27675 23109
rect 27617 23100 27629 23103
rect 25823 23072 27629 23100
rect 25823 23069 25835 23072
rect 25777 23063 25835 23069
rect 27617 23069 27629 23072
rect 27663 23100 27675 23103
rect 28258 23100 28264 23112
rect 27663 23072 28264 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 32217 23103 32275 23109
rect 32217 23069 32229 23103
rect 32263 23100 32275 23103
rect 32398 23100 32404 23112
rect 32263 23072 32404 23100
rect 32263 23069 32275 23072
rect 32217 23063 32275 23069
rect 32398 23060 32404 23072
rect 32456 23060 32462 23112
rect 20622 22992 20628 23044
rect 20680 23032 20686 23044
rect 20993 23035 21051 23041
rect 20993 23032 21005 23035
rect 20680 23004 21005 23032
rect 20680 22992 20686 23004
rect 20993 23001 21005 23004
rect 21039 23001 21051 23035
rect 20993 22995 21051 23001
rect 21177 23035 21235 23041
rect 21177 23001 21189 23035
rect 21223 23032 21235 23035
rect 22002 23032 22008 23044
rect 21223 23004 22008 23032
rect 21223 23001 21235 23004
rect 21177 22995 21235 23001
rect 22002 22992 22008 23004
rect 22060 22992 22066 23044
rect 26050 23041 26056 23044
rect 26044 22995 26056 23041
rect 26108 23032 26114 23044
rect 26108 23004 26144 23032
rect 26050 22992 26056 22995
rect 26108 22992 26114 23004
rect 27157 22967 27215 22973
rect 27157 22933 27169 22967
rect 27203 22964 27215 22967
rect 27246 22964 27252 22976
rect 27203 22936 27252 22964
rect 27203 22933 27215 22936
rect 27157 22927 27215 22933
rect 27246 22924 27252 22936
rect 27304 22924 27310 22976
rect 37550 22964 37556 22976
rect 37511 22936 37556 22964
rect 37550 22924 37556 22936
rect 37608 22924 37614 22976
rect 37642 22924 37648 22976
rect 37700 22964 37706 22976
rect 38013 22967 38071 22973
rect 38013 22964 38025 22967
rect 37700 22936 38025 22964
rect 37700 22924 37706 22936
rect 38013 22933 38025 22936
rect 38059 22933 38071 22967
rect 38013 22927 38071 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 25961 22763 26019 22769
rect 20588 22732 22324 22760
rect 20588 22720 20594 22732
rect 20622 22652 20628 22704
rect 20680 22692 20686 22704
rect 22296 22692 22324 22732
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26050 22760 26056 22772
rect 26007 22732 26056 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 26050 22720 26056 22732
rect 26108 22720 26114 22772
rect 32674 22720 32680 22772
rect 32732 22760 32738 22772
rect 33229 22763 33287 22769
rect 33229 22760 33241 22763
rect 32732 22732 33241 22760
rect 32732 22720 32738 22732
rect 33229 22729 33241 22732
rect 33275 22729 33287 22763
rect 33229 22723 33287 22729
rect 35621 22695 35679 22701
rect 20680 22664 22140 22692
rect 22296 22664 34928 22692
rect 20680 22652 20686 22664
rect 22002 22624 22008 22636
rect 21963 22596 22008 22624
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 22112 22633 22140 22664
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 25188 22596 26157 22624
rect 25188 22584 25194 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 32674 22584 32680 22636
rect 32732 22624 32738 22636
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 32732 22596 33609 22624
rect 32732 22584 32738 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22624 33747 22627
rect 34790 22624 34796 22636
rect 33735 22596 34796 22624
rect 33735 22593 33747 22596
rect 33689 22587 33747 22593
rect 34790 22584 34796 22596
rect 34848 22584 34854 22636
rect 34900 22624 34928 22664
rect 35621 22661 35633 22695
rect 35667 22692 35679 22695
rect 35894 22692 35900 22704
rect 35667 22664 35900 22692
rect 35667 22661 35679 22664
rect 35621 22655 35679 22661
rect 35894 22652 35900 22664
rect 35952 22652 35958 22704
rect 37550 22652 37556 22704
rect 37608 22692 37614 22704
rect 37829 22695 37887 22701
rect 37829 22692 37841 22695
rect 37608 22664 37841 22692
rect 37608 22652 37614 22664
rect 37829 22661 37841 22664
rect 37875 22692 37887 22695
rect 38194 22692 38200 22704
rect 37875 22664 38200 22692
rect 37875 22661 37887 22664
rect 37829 22655 37887 22661
rect 38194 22652 38200 22664
rect 38252 22652 38258 22704
rect 37645 22627 37703 22633
rect 37645 22624 37657 22627
rect 34900 22596 37657 22624
rect 37645 22593 37657 22596
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 26421 22559 26479 22565
rect 26421 22525 26433 22559
rect 26467 22556 26479 22559
rect 27246 22556 27252 22568
rect 26467 22528 27252 22556
rect 26467 22525 26479 22528
rect 26421 22519 26479 22525
rect 27246 22516 27252 22528
rect 27304 22516 27310 22568
rect 32122 22516 32128 22568
rect 32180 22556 32186 22568
rect 32398 22556 32404 22568
rect 32180 22528 32404 22556
rect 32180 22516 32186 22528
rect 32398 22516 32404 22528
rect 32456 22556 32462 22568
rect 33873 22559 33931 22565
rect 33873 22556 33885 22559
rect 32456 22528 33885 22556
rect 32456 22516 32462 22528
rect 33873 22525 33885 22528
rect 33919 22556 33931 22559
rect 37918 22556 37924 22568
rect 33919 22528 37924 22556
rect 33919 22525 33931 22528
rect 33873 22519 33931 22525
rect 37918 22516 37924 22528
rect 37976 22516 37982 22568
rect 17218 22448 17224 22500
rect 17276 22488 17282 22500
rect 35069 22491 35127 22497
rect 35069 22488 35081 22491
rect 17276 22460 35081 22488
rect 17276 22448 17282 22460
rect 35069 22457 35081 22460
rect 35115 22488 35127 22491
rect 35897 22491 35955 22497
rect 35897 22488 35909 22491
rect 35115 22460 35909 22488
rect 35115 22457 35127 22460
rect 35069 22451 35127 22457
rect 35897 22457 35909 22460
rect 35943 22457 35955 22491
rect 35897 22451 35955 22457
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21048 22392 21833 22420
rect 21048 22380 21054 22392
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 26329 22423 26387 22429
rect 26329 22389 26341 22423
rect 26375 22420 26387 22423
rect 26418 22420 26424 22432
rect 26375 22392 26424 22420
rect 26375 22389 26387 22392
rect 26329 22383 26387 22389
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 32030 22380 32036 22432
rect 32088 22420 32094 22432
rect 32674 22420 32680 22432
rect 32088 22392 32680 22420
rect 32088 22380 32094 22392
rect 32674 22380 32680 22392
rect 32732 22380 32738 22432
rect 36078 22420 36084 22432
rect 36039 22392 36084 22420
rect 36078 22380 36084 22392
rect 36136 22380 36142 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 5997 22151 6055 22157
rect 5997 22117 6009 22151
rect 6043 22117 6055 22151
rect 31386 22148 31392 22160
rect 5997 22111 6055 22117
rect 31220 22120 31392 22148
rect 6012 22080 6040 22111
rect 6914 22080 6920 22092
rect 6012 22052 6920 22080
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 17954 22040 17960 22092
rect 18012 22080 18018 22092
rect 20809 22083 20867 22089
rect 20809 22080 20821 22083
rect 18012 22052 20821 22080
rect 18012 22040 18018 22052
rect 20809 22049 20821 22052
rect 20855 22049 20867 22083
rect 20809 22043 20867 22049
rect 21177 22083 21235 22089
rect 21177 22049 21189 22083
rect 21223 22080 21235 22083
rect 21266 22080 21272 22092
rect 21223 22052 21272 22080
rect 21223 22049 21235 22052
rect 21177 22043 21235 22049
rect 21266 22040 21272 22052
rect 21324 22080 21330 22092
rect 23290 22080 23296 22092
rect 21324 22052 23296 22080
rect 21324 22040 21330 22052
rect 23290 22040 23296 22052
rect 23348 22040 23354 22092
rect 31220 22089 31248 22120
rect 31386 22108 31392 22120
rect 31444 22108 31450 22160
rect 31205 22083 31263 22089
rect 31205 22049 31217 22083
rect 31251 22080 31263 22083
rect 31251 22052 31285 22080
rect 31251 22049 31263 22052
rect 31205 22043 31263 22049
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 22012 4675 22015
rect 4663 21984 6592 22012
rect 4663 21981 4675 21984
rect 4617 21975 4675 21981
rect 4884 21947 4942 21953
rect 4884 21913 4896 21947
rect 4930 21944 4942 21947
rect 6362 21944 6368 21956
rect 4930 21916 6368 21944
rect 4930 21913 4942 21916
rect 4884 21907 4942 21913
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 6564 21888 6592 21984
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 20990 22012 20996 22024
rect 20680 21984 20996 22012
rect 20680 21972 20686 21984
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 37461 22015 37519 22021
rect 37461 21981 37473 22015
rect 37507 22012 37519 22015
rect 38102 22012 38108 22024
rect 37507 21984 38108 22012
rect 37507 21981 37519 21984
rect 37461 21975 37519 21981
rect 38102 21972 38108 21984
rect 38160 21972 38166 22024
rect 30929 21947 30987 21953
rect 30929 21944 30941 21947
rect 30300 21916 30941 21944
rect 30300 21888 30328 21916
rect 30929 21913 30941 21916
rect 30975 21913 30987 21947
rect 30929 21907 30987 21913
rect 34790 21904 34796 21956
rect 34848 21944 34854 21956
rect 34848 21916 37964 21944
rect 34848 21904 34854 21916
rect 6546 21876 6552 21888
rect 6507 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 30101 21879 30159 21885
rect 30101 21845 30113 21879
rect 30147 21876 30159 21879
rect 30282 21876 30288 21888
rect 30147 21848 30288 21876
rect 30147 21845 30159 21848
rect 30101 21839 30159 21845
rect 30282 21836 30288 21848
rect 30340 21836 30346 21888
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 30561 21879 30619 21885
rect 30561 21876 30573 21879
rect 30524 21848 30573 21876
rect 30524 21836 30530 21848
rect 30561 21845 30573 21848
rect 30607 21845 30619 21879
rect 30561 21839 30619 21845
rect 31021 21879 31079 21885
rect 31021 21845 31033 21879
rect 31067 21876 31079 21879
rect 33042 21876 33048 21888
rect 31067 21848 33048 21876
rect 31067 21845 31079 21848
rect 31021 21839 31079 21845
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 37936 21885 37964 21916
rect 37921 21879 37979 21885
rect 37921 21845 37933 21879
rect 37967 21845 37979 21879
rect 37921 21839 37979 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 3421 21675 3479 21681
rect 3421 21641 3433 21675
rect 3467 21672 3479 21675
rect 4614 21672 4620 21684
rect 3467 21644 4620 21672
rect 3467 21641 3479 21644
rect 3421 21635 3479 21641
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 2056 21576 4016 21604
rect 2056 21545 2084 21576
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21505 2099 21539
rect 2041 21499 2099 21505
rect 2308 21539 2366 21545
rect 2308 21505 2320 21539
rect 2354 21536 2366 21539
rect 2774 21536 2780 21548
rect 2354 21508 2780 21536
rect 2354 21505 2366 21508
rect 2308 21499 2366 21505
rect 2774 21496 2780 21508
rect 2832 21496 2838 21548
rect 3988 21341 4016 21576
rect 23290 21564 23296 21616
rect 23348 21604 23354 21616
rect 23385 21607 23443 21613
rect 23385 21604 23397 21607
rect 23348 21576 23397 21604
rect 23348 21564 23354 21576
rect 23385 21573 23397 21576
rect 23431 21573 23443 21607
rect 23385 21567 23443 21573
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 23658 21536 23664 21548
rect 23615 21508 23664 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 3973 21335 4031 21341
rect 3973 21301 3985 21335
rect 4019 21332 4031 21335
rect 6546 21332 6552 21344
rect 4019 21304 6552 21332
rect 4019 21301 4031 21304
rect 3973 21295 4031 21301
rect 6546 21292 6552 21304
rect 6604 21332 6610 21344
rect 10410 21332 10416 21344
rect 6604 21304 10416 21332
rect 6604 21292 6610 21304
rect 10410 21292 10416 21304
rect 10468 21292 10474 21344
rect 33134 21292 33140 21344
rect 33192 21332 33198 21344
rect 34698 21332 34704 21344
rect 33192 21304 34704 21332
rect 33192 21292 33198 21304
rect 34698 21292 34704 21304
rect 34756 21292 34762 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 6362 21128 6368 21140
rect 6323 21100 6368 21128
rect 6362 21088 6368 21100
rect 6420 21088 6426 21140
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 6546 20992 6552 21004
rect 5684 20964 6552 20992
rect 5684 20952 5690 20964
rect 6546 20952 6552 20964
rect 6604 20952 6610 21004
rect 6641 20995 6699 21001
rect 6641 20961 6653 20995
rect 6687 20992 6699 20995
rect 7285 20995 7343 21001
rect 7285 20992 7297 20995
rect 6687 20964 7297 20992
rect 6687 20961 6699 20964
rect 6641 20955 6699 20961
rect 7285 20961 7297 20964
rect 7331 20992 7343 20995
rect 10226 20992 10232 21004
rect 7331 20964 10232 20992
rect 7331 20961 7343 20964
rect 7285 20955 7343 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 36078 20952 36084 21004
rect 36136 20992 36142 21004
rect 37001 20995 37059 21001
rect 37001 20992 37013 20995
rect 36136 20964 37013 20992
rect 36136 20952 36142 20964
rect 37001 20961 37013 20964
rect 37047 20961 37059 20995
rect 37001 20955 37059 20961
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 6788 20896 6833 20924
rect 10428 20896 10977 20924
rect 6788 20884 6794 20896
rect 10428 20800 10456 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 37090 20884 37096 20936
rect 37148 20924 37154 20936
rect 37277 20927 37335 20933
rect 37277 20924 37289 20927
rect 37148 20896 37289 20924
rect 37148 20884 37154 20896
rect 37277 20893 37289 20896
rect 37323 20893 37335 20927
rect 37277 20887 37335 20893
rect 11054 20816 11060 20868
rect 11112 20856 11118 20868
rect 11210 20859 11268 20865
rect 11210 20856 11222 20859
rect 11112 20828 11222 20856
rect 11112 20816 11118 20828
rect 11210 20825 11222 20828
rect 11256 20825 11268 20859
rect 11210 20819 11268 20825
rect 10410 20788 10416 20800
rect 10371 20760 10416 20788
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 12345 20791 12403 20797
rect 12345 20757 12357 20791
rect 12391 20788 12403 20791
rect 13078 20788 13084 20800
rect 12391 20760 13084 20788
rect 12391 20757 12403 20760
rect 12345 20751 12403 20757
rect 13078 20748 13084 20760
rect 13136 20748 13142 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 6733 20587 6791 20593
rect 6733 20553 6745 20587
rect 6779 20584 6791 20587
rect 7006 20584 7012 20596
rect 6779 20556 7012 20584
rect 6779 20553 6791 20556
rect 6733 20547 6791 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 11054 20584 11060 20596
rect 10183 20556 11060 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 33042 20544 33048 20596
rect 33100 20584 33106 20596
rect 37921 20587 37979 20593
rect 37921 20584 37933 20587
rect 33100 20556 37933 20584
rect 33100 20544 33106 20556
rect 37921 20553 37933 20556
rect 37967 20553 37979 20587
rect 37921 20547 37979 20553
rect 4614 20476 4620 20528
rect 4672 20516 4678 20528
rect 6917 20519 6975 20525
rect 6917 20516 6929 20519
rect 4672 20488 6929 20516
rect 4672 20476 4678 20488
rect 6917 20485 6929 20488
rect 6963 20485 6975 20519
rect 6917 20479 6975 20485
rect 28445 20519 28503 20525
rect 28445 20485 28457 20519
rect 28491 20516 28503 20519
rect 28994 20516 29000 20528
rect 28491 20488 29000 20516
rect 28491 20485 28503 20488
rect 28445 20479 28503 20485
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20448 6883 20451
rect 7466 20448 7472 20460
rect 6871 20420 7472 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 10226 20408 10232 20460
rect 10284 20448 10290 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10284 20420 10425 20448
rect 10284 20408 10290 20420
rect 10413 20417 10425 20420
rect 10459 20448 10471 20451
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 10459 20420 11529 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 11517 20417 11529 20420
rect 11563 20448 11575 20451
rect 15194 20448 15200 20460
rect 11563 20420 12434 20448
rect 15155 20420 15200 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7101 20383 7159 20389
rect 7101 20380 7113 20383
rect 6972 20352 7113 20380
rect 6972 20340 6978 20352
rect 7101 20349 7113 20352
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 7432 20352 10333 20380
rect 7432 20340 7438 20352
rect 10321 20349 10333 20352
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20380 10563 20383
rect 12250 20380 12256 20392
rect 10551 20352 12256 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 12406 20312 12434 20420
rect 15194 20408 15200 20420
rect 15252 20448 15258 20460
rect 15838 20448 15844 20460
rect 15252 20420 15844 20448
rect 15252 20408 15258 20420
rect 15838 20408 15844 20420
rect 15896 20448 15902 20460
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 15896 20420 15945 20448
rect 15896 20408 15902 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 37461 20451 37519 20457
rect 37461 20417 37473 20451
rect 37507 20448 37519 20451
rect 38102 20448 38108 20460
rect 37507 20420 38108 20448
rect 37507 20417 37519 20420
rect 37461 20411 37519 20417
rect 38102 20408 38108 20420
rect 38160 20408 38166 20460
rect 15381 20315 15439 20321
rect 15381 20312 15393 20315
rect 12406 20284 15393 20312
rect 15381 20281 15393 20284
rect 15427 20312 15439 20315
rect 25590 20312 25596 20324
rect 15427 20284 25596 20312
rect 15427 20281 15439 20284
rect 15381 20275 15439 20281
rect 25590 20272 25596 20284
rect 25648 20272 25654 20324
rect 28258 20312 28264 20324
rect 28219 20284 28264 20312
rect 28258 20272 28264 20284
rect 28316 20272 28322 20324
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 6730 20000 6736 20052
rect 6788 20040 6794 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6788 20012 6837 20040
rect 6788 20000 6794 20012
rect 6825 20009 6837 20012
rect 6871 20009 6883 20043
rect 6825 20003 6883 20009
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10410 20040 10416 20052
rect 10100 20012 10416 20040
rect 10100 20000 10106 20012
rect 10410 20000 10416 20012
rect 10468 20040 10474 20052
rect 10468 20012 15516 20040
rect 10468 20000 10474 20012
rect 6914 19932 6920 19984
rect 6972 19972 6978 19984
rect 6972 19944 7328 19972
rect 6972 19932 6978 19944
rect 4157 19907 4215 19913
rect 4157 19873 4169 19907
rect 4203 19904 4215 19907
rect 4798 19904 4804 19916
rect 4203 19876 4804 19904
rect 4203 19873 4215 19876
rect 4157 19867 4215 19873
rect 4798 19864 4804 19876
rect 4856 19904 4862 19916
rect 7300 19913 7328 19944
rect 7466 19932 7472 19984
rect 7524 19972 7530 19984
rect 8202 19972 8208 19984
rect 7524 19944 8208 19972
rect 7524 19932 7530 19944
rect 8202 19932 8208 19944
rect 8260 19972 8266 19984
rect 12529 19975 12587 19981
rect 12529 19972 12541 19975
rect 8260 19944 12541 19972
rect 8260 19932 8266 19944
rect 12529 19941 12541 19944
rect 12575 19941 12587 19975
rect 13078 19972 13084 19984
rect 13039 19944 13084 19972
rect 12529 19935 12587 19941
rect 13078 19932 13084 19944
rect 13136 19932 13142 19984
rect 7193 19907 7251 19913
rect 7193 19904 7205 19907
rect 4856 19876 7205 19904
rect 4856 19864 4862 19876
rect 7193 19873 7205 19876
rect 7239 19873 7251 19907
rect 7193 19867 7251 19873
rect 7285 19907 7343 19913
rect 7285 19873 7297 19907
rect 7331 19873 7343 19907
rect 7285 19867 7343 19873
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 4614 19836 4620 19848
rect 4387 19808 4620 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 7006 19836 7012 19848
rect 6919 19808 7012 19836
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7374 19836 7380 19848
rect 7147 19808 7380 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 10134 19836 10140 19848
rect 10095 19808 10140 19836
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 15488 19845 15516 20012
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 18012 20012 18153 20040
rect 18012 20000 18018 20012
rect 18141 20009 18153 20012
rect 18187 20009 18199 20043
rect 18141 20003 18199 20009
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 26697 20043 26755 20049
rect 26697 20040 26709 20043
rect 23716 20012 26709 20040
rect 23716 20000 23722 20012
rect 26697 20009 26709 20012
rect 26743 20009 26755 20043
rect 26697 20003 26755 20009
rect 17313 19975 17371 19981
rect 17313 19941 17325 19975
rect 17359 19972 17371 19975
rect 23017 19975 23075 19981
rect 17359 19944 18276 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 18248 19913 18276 19944
rect 23017 19941 23029 19975
rect 23063 19972 23075 19975
rect 23290 19972 23296 19984
rect 23063 19944 23296 19972
rect 23063 19941 23075 19944
rect 23017 19935 23075 19941
rect 23290 19932 23296 19944
rect 23348 19932 23354 19984
rect 27246 19972 27252 19984
rect 27207 19944 27252 19972
rect 27246 19932 27252 19944
rect 27304 19932 27310 19984
rect 30024 19944 30972 19972
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 19978 19904 19984 19916
rect 18279 19876 19984 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 25590 19864 25596 19916
rect 25648 19904 25654 19916
rect 30024 19904 30052 19944
rect 25648 19876 30052 19904
rect 30116 19876 30880 19904
rect 25648 19864 25654 19876
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12584 19808 12725 19836
rect 12584 19796 12590 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19836 15531 19839
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15519 19808 15945 19836
rect 15519 19805 15531 19808
rect 15473 19799 15531 19805
rect 15933 19805 15945 19808
rect 15979 19836 15991 19839
rect 16758 19836 16764 19848
rect 15979 19808 16764 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 23106 19796 23112 19848
rect 23164 19836 23170 19848
rect 23293 19839 23351 19845
rect 23293 19836 23305 19839
rect 23164 19808 23305 19836
rect 23164 19796 23170 19808
rect 23293 19805 23305 19808
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 27154 19796 27160 19848
rect 27212 19836 27218 19848
rect 30116 19845 30144 19876
rect 30852 19845 30880 19876
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 27212 19808 30113 19836
rect 27212 19796 27218 19808
rect 30101 19805 30113 19808
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 30377 19839 30435 19845
rect 30377 19805 30389 19839
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 30837 19839 30895 19845
rect 30837 19805 30849 19839
rect 30883 19805 30895 19839
rect 30944 19836 30972 19944
rect 31021 19839 31079 19845
rect 31021 19836 31033 19839
rect 30944 19808 31033 19836
rect 30837 19799 30895 19805
rect 31021 19805 31033 19808
rect 31067 19836 31079 19839
rect 31481 19839 31539 19845
rect 31481 19836 31493 19839
rect 31067 19808 31493 19836
rect 31067 19805 31079 19808
rect 31021 19799 31079 19805
rect 31481 19805 31493 19808
rect 31527 19836 31539 19839
rect 33410 19836 33416 19848
rect 31527 19808 33416 19836
rect 31527 19805 31539 19808
rect 31481 19799 31539 19805
rect 7024 19768 7052 19796
rect 7558 19768 7564 19780
rect 7024 19740 7564 19768
rect 7558 19728 7564 19740
rect 7616 19728 7622 19780
rect 16200 19771 16258 19777
rect 16200 19737 16212 19771
rect 16246 19768 16258 19771
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 16246 19740 17785 19768
rect 16246 19737 16258 19740
rect 16200 19731 16258 19737
rect 17773 19737 17785 19740
rect 17819 19737 17831 19771
rect 22557 19771 22615 19777
rect 22557 19768 22569 19771
rect 17773 19731 17831 19737
rect 22066 19740 22569 19768
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 12802 19700 12808 19712
rect 12763 19672 12808 19700
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 12952 19672 12997 19700
rect 12952 19660 12958 19672
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 22066 19700 22094 19740
rect 22557 19737 22569 19740
rect 22603 19768 22615 19771
rect 23017 19771 23075 19777
rect 23017 19768 23029 19771
rect 22603 19740 23029 19768
rect 22603 19737 22615 19740
rect 22557 19731 22615 19737
rect 23017 19737 23029 19740
rect 23063 19737 23075 19771
rect 23017 19731 23075 19737
rect 26881 19771 26939 19777
rect 26881 19737 26893 19771
rect 26927 19768 26939 19771
rect 30190 19768 30196 19780
rect 26927 19740 30196 19768
rect 26927 19737 26939 19740
rect 26881 19731 26939 19737
rect 30190 19728 30196 19740
rect 30248 19768 30254 19780
rect 30392 19768 30420 19799
rect 33410 19796 33416 19808
rect 33468 19796 33474 19848
rect 30248 19740 30420 19768
rect 30248 19728 30254 19740
rect 17736 19672 22094 19700
rect 17736 19660 17742 19672
rect 22830 19660 22836 19712
rect 22888 19700 22894 19712
rect 23201 19703 23259 19709
rect 23201 19700 23213 19703
rect 22888 19672 23213 19700
rect 22888 19660 22894 19672
rect 23201 19669 23213 19672
rect 23247 19669 23259 19703
rect 23201 19663 23259 19669
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 26973 19703 27031 19709
rect 26973 19700 26985 19703
rect 26292 19672 26985 19700
rect 26292 19660 26298 19672
rect 26973 19669 26985 19672
rect 27019 19669 27031 19703
rect 26973 19663 27031 19669
rect 27065 19703 27123 19709
rect 27065 19669 27077 19703
rect 27111 19700 27123 19703
rect 27246 19700 27252 19712
rect 27111 19672 27252 19700
rect 27111 19669 27123 19672
rect 27065 19663 27123 19669
rect 27246 19660 27252 19672
rect 27304 19660 27310 19712
rect 30926 19700 30932 19712
rect 30887 19672 30932 19700
rect 30926 19660 30932 19672
rect 30984 19660 30990 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 12250 19496 12256 19508
rect 12211 19468 12256 19496
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 19978 19496 19984 19508
rect 19939 19468 19984 19496
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 26418 19456 26424 19508
rect 26476 19496 26482 19508
rect 26973 19499 27031 19505
rect 26973 19496 26985 19499
rect 26476 19468 26985 19496
rect 26476 19456 26482 19468
rect 26973 19465 26985 19468
rect 27019 19465 27031 19499
rect 30190 19496 30196 19508
rect 30151 19468 30196 19496
rect 26973 19459 27031 19465
rect 30190 19456 30196 19468
rect 30248 19456 30254 19508
rect 33410 19496 33416 19508
rect 33371 19468 33416 19496
rect 33410 19456 33416 19468
rect 33468 19456 33474 19508
rect 34333 19499 34391 19505
rect 34333 19465 34345 19499
rect 34379 19496 34391 19499
rect 35986 19496 35992 19508
rect 34379 19468 35992 19496
rect 34379 19465 34391 19468
rect 34333 19459 34391 19465
rect 35986 19456 35992 19468
rect 36044 19496 36050 19508
rect 36265 19499 36323 19505
rect 36265 19496 36277 19499
rect 36044 19468 36277 19496
rect 36044 19456 36050 19468
rect 36265 19465 36277 19468
rect 36311 19465 36323 19499
rect 36265 19459 36323 19465
rect 12526 19428 12532 19440
rect 12452 19400 12532 19428
rect 12452 19369 12480 19400
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 12802 19428 12808 19440
rect 12636 19400 12808 19428
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12636 19360 12664 19400
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 19886 19428 19892 19440
rect 19799 19400 19892 19428
rect 19886 19388 19892 19400
rect 19944 19428 19950 19440
rect 23658 19428 23664 19440
rect 19944 19400 23664 19428
rect 19944 19388 19950 19400
rect 23658 19388 23664 19400
rect 23716 19388 23722 19440
rect 27154 19437 27160 19440
rect 27125 19431 27160 19437
rect 27125 19428 27137 19431
rect 26160 19400 27137 19428
rect 12437 19323 12495 19329
rect 12544 19332 12664 19360
rect 12713 19363 12771 19369
rect 12544 19301 12572 19332
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13078 19360 13084 19372
rect 12759 19332 13084 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 17828 19332 19625 19360
rect 17828 19320 17834 19332
rect 19613 19329 19625 19332
rect 19659 19329 19671 19363
rect 19794 19360 19800 19372
rect 19755 19332 19800 19360
rect 19613 19323 19671 19329
rect 19794 19320 19800 19332
rect 19852 19360 19858 19372
rect 20622 19360 20628 19372
rect 19852 19332 20628 19360
rect 19852 19320 19858 19332
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 23106 19320 23112 19372
rect 23164 19360 23170 19372
rect 26160 19369 26188 19400
rect 27125 19397 27137 19400
rect 27125 19391 27160 19397
rect 27154 19388 27160 19391
rect 27212 19388 27218 19440
rect 27246 19388 27252 19440
rect 27304 19428 27310 19440
rect 27341 19431 27399 19437
rect 27341 19428 27353 19431
rect 27304 19400 27353 19428
rect 27304 19388 27310 19400
rect 27341 19397 27353 19400
rect 27387 19397 27399 19431
rect 34698 19428 34704 19440
rect 27341 19391 27399 19397
rect 29656 19400 34704 19428
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 23164 19332 26157 19360
rect 23164 19320 23170 19332
rect 26145 19329 26157 19332
rect 26191 19329 26203 19363
rect 26145 19323 26203 19329
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26421 19363 26479 19369
rect 26292 19332 26385 19360
rect 26292 19320 26298 19332
rect 26421 19329 26433 19363
rect 26467 19360 26479 19363
rect 27264 19360 27292 19388
rect 26467 19332 27292 19360
rect 26467 19329 26479 19332
rect 26421 19323 26479 19329
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12621 19295 12679 19301
rect 12621 19261 12633 19295
rect 12667 19292 12679 19295
rect 12894 19292 12900 19304
rect 12667 19264 12900 19292
rect 12667 19261 12679 19264
rect 12621 19255 12679 19261
rect 12636 19224 12664 19255
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 26252 19292 26280 19320
rect 22888 19264 26280 19292
rect 22888 19252 22894 19264
rect 20162 19224 20168 19236
rect 12544 19196 12664 19224
rect 20123 19196 20168 19224
rect 12544 19168 12572 19196
rect 20162 19184 20168 19196
rect 20220 19184 20226 19236
rect 26252 19224 26280 19264
rect 26252 19196 27200 19224
rect 12526 19116 12532 19168
rect 12584 19116 12590 19168
rect 26234 19116 26240 19168
rect 26292 19156 26298 19168
rect 27172 19165 27200 19196
rect 26421 19159 26479 19165
rect 26421 19156 26433 19159
rect 26292 19128 26433 19156
rect 26292 19116 26298 19128
rect 26421 19125 26433 19128
rect 26467 19125 26479 19159
rect 26421 19119 26479 19125
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19125 27215 19159
rect 27157 19119 27215 19125
rect 28258 19116 28264 19168
rect 28316 19156 28322 19168
rect 29656 19165 29684 19400
rect 30926 19320 30932 19372
rect 30984 19360 30990 19372
rect 31588 19369 31616 19400
rect 34698 19388 34704 19400
rect 34756 19428 34762 19440
rect 36280 19428 36308 19459
rect 37461 19431 37519 19437
rect 37461 19428 37473 19431
rect 34756 19400 34928 19428
rect 36280 19400 37473 19428
rect 34756 19388 34762 19400
rect 31306 19363 31364 19369
rect 31306 19360 31318 19363
rect 30984 19332 31318 19360
rect 30984 19320 30990 19332
rect 31306 19329 31318 19332
rect 31352 19329 31364 19363
rect 31306 19323 31364 19329
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19329 31631 19363
rect 31573 19323 31631 19329
rect 33410 19320 33416 19372
rect 33468 19360 33474 19372
rect 34149 19363 34207 19369
rect 34149 19360 34161 19363
rect 33468 19332 34161 19360
rect 33468 19320 33474 19332
rect 34149 19329 34161 19332
rect 34195 19329 34207 19363
rect 34149 19323 34207 19329
rect 34425 19363 34483 19369
rect 34425 19329 34437 19363
rect 34471 19360 34483 19363
rect 34790 19360 34796 19372
rect 34471 19332 34796 19360
rect 34471 19329 34483 19332
rect 34425 19323 34483 19329
rect 34790 19320 34796 19332
rect 34848 19320 34854 19372
rect 34900 19369 34928 19400
rect 37461 19397 37473 19400
rect 37507 19397 37519 19431
rect 37461 19391 37519 19397
rect 34885 19363 34943 19369
rect 34885 19329 34897 19363
rect 34931 19329 34943 19363
rect 35141 19363 35199 19369
rect 35141 19360 35153 19363
rect 34885 19323 34943 19329
rect 34992 19332 35153 19360
rect 33965 19295 34023 19301
rect 33965 19261 33977 19295
rect 34011 19292 34023 19295
rect 34992 19292 35020 19332
rect 35141 19329 35153 19332
rect 35187 19329 35199 19363
rect 35141 19323 35199 19329
rect 37550 19320 37556 19372
rect 37608 19360 37614 19372
rect 37645 19363 37703 19369
rect 37645 19360 37657 19363
rect 37608 19332 37657 19360
rect 37608 19320 37614 19332
rect 37645 19329 37657 19332
rect 37691 19329 37703 19363
rect 37645 19323 37703 19329
rect 34011 19264 35020 19292
rect 37277 19295 37335 19301
rect 34011 19261 34023 19264
rect 33965 19255 34023 19261
rect 37277 19261 37289 19295
rect 37323 19292 37335 19295
rect 38470 19292 38476 19304
rect 37323 19264 38476 19292
rect 37323 19261 37335 19264
rect 37277 19255 37335 19261
rect 38470 19252 38476 19264
rect 38528 19252 38534 19304
rect 29641 19159 29699 19165
rect 29641 19156 29653 19159
rect 28316 19128 29653 19156
rect 28316 19116 28322 19128
rect 29641 19125 29653 19128
rect 29687 19125 29699 19159
rect 29641 19119 29699 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 19797 18955 19855 18961
rect 19797 18921 19809 18955
rect 19843 18952 19855 18955
rect 19886 18952 19892 18964
rect 19843 18924 19892 18952
rect 19843 18921 19855 18924
rect 19797 18915 19855 18921
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 23106 18952 23112 18964
rect 23067 18924 23112 18952
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 25590 18912 25596 18964
rect 25648 18952 25654 18964
rect 25685 18955 25743 18961
rect 25685 18952 25697 18955
rect 25648 18924 25697 18952
rect 25648 18912 25654 18924
rect 25685 18921 25697 18924
rect 25731 18952 25743 18955
rect 34698 18952 34704 18964
rect 25731 18924 26556 18952
rect 34659 18924 34704 18952
rect 25731 18921 25743 18924
rect 25685 18915 25743 18921
rect 26329 18887 26387 18893
rect 26329 18853 26341 18887
rect 26375 18884 26387 18887
rect 26418 18884 26424 18896
rect 26375 18856 26424 18884
rect 26375 18853 26387 18856
rect 26329 18847 26387 18853
rect 26418 18844 26424 18856
rect 26476 18844 26482 18896
rect 26528 18825 26556 18924
rect 34698 18912 34704 18924
rect 34756 18912 34762 18964
rect 26513 18819 26571 18825
rect 26513 18785 26525 18819
rect 26559 18785 26571 18819
rect 26513 18779 26571 18785
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 22830 18748 22836 18760
rect 22428 18720 22836 18748
rect 22428 18708 22434 18720
rect 22830 18708 22836 18720
rect 22888 18748 22894 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22888 18720 23029 18748
rect 22888 18708 22894 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23290 18748 23296 18760
rect 23251 18720 23296 18748
rect 23017 18711 23075 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 26234 18748 26240 18760
rect 26195 18720 26240 18748
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 37461 18751 37519 18757
rect 37461 18717 37473 18751
rect 37507 18748 37519 18751
rect 38102 18748 38108 18760
rect 37507 18720 38108 18748
rect 37507 18717 37519 18720
rect 37461 18711 37519 18717
rect 38102 18708 38108 18720
rect 38160 18708 38166 18760
rect 19794 18689 19800 18692
rect 19781 18683 19800 18689
rect 19781 18649 19793 18683
rect 19781 18643 19800 18649
rect 19794 18640 19800 18643
rect 19852 18640 19858 18692
rect 19978 18680 19984 18692
rect 19939 18652 19984 18680
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 34422 18640 34428 18692
rect 34480 18680 34486 18692
rect 34480 18652 37964 18680
rect 34480 18640 34486 18652
rect 18046 18572 18052 18624
rect 18104 18612 18110 18624
rect 18874 18612 18880 18624
rect 18104 18584 18880 18612
rect 18104 18572 18110 18584
rect 18874 18572 18880 18584
rect 18932 18612 18938 18624
rect 19613 18615 19671 18621
rect 19613 18612 19625 18615
rect 18932 18584 19625 18612
rect 18932 18572 18938 18584
rect 19613 18581 19625 18584
rect 19659 18581 19671 18615
rect 23474 18612 23480 18624
rect 23435 18584 23480 18612
rect 19613 18575 19671 18581
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 26050 18572 26056 18624
rect 26108 18612 26114 18624
rect 37936 18621 37964 18652
rect 26237 18615 26295 18621
rect 26237 18612 26249 18615
rect 26108 18584 26249 18612
rect 26108 18572 26114 18584
rect 26237 18581 26249 18584
rect 26283 18581 26295 18615
rect 26237 18575 26295 18581
rect 37921 18615 37979 18621
rect 37921 18581 37933 18615
rect 37967 18581 37979 18615
rect 37921 18575 37979 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 2961 18411 3019 18417
rect 2961 18408 2973 18411
rect 2832 18380 2973 18408
rect 2832 18368 2838 18380
rect 2961 18377 2973 18380
rect 3007 18377 3019 18411
rect 2961 18371 3019 18377
rect 17773 18411 17831 18417
rect 17773 18377 17785 18411
rect 17819 18408 17831 18411
rect 17954 18408 17960 18420
rect 17819 18380 17960 18408
rect 17819 18377 17831 18380
rect 17773 18371 17831 18377
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 3142 18272 3148 18284
rect 3103 18244 3148 18272
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 17678 18272 17684 18284
rect 17639 18244 17684 18272
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 18046 18272 18052 18284
rect 17911 18244 18052 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 4798 18204 4804 18216
rect 3467 18176 4804 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 3329 18071 3387 18077
rect 3329 18037 3341 18071
rect 3375 18068 3387 18071
rect 3970 18068 3976 18080
rect 3375 18040 3976 18068
rect 3375 18037 3387 18040
rect 3329 18031 3387 18037
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 3142 17824 3148 17876
rect 3200 17864 3206 17876
rect 3237 17867 3295 17873
rect 3237 17864 3249 17867
rect 3200 17836 3249 17864
rect 3200 17824 3206 17836
rect 3237 17833 3249 17836
rect 3283 17833 3295 17867
rect 3237 17827 3295 17833
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 8297 17867 8355 17873
rect 8297 17864 8309 17867
rect 7432 17836 8309 17864
rect 7432 17824 7438 17836
rect 8297 17833 8309 17836
rect 8343 17833 8355 17867
rect 8297 17827 8355 17833
rect 9769 17867 9827 17873
rect 9769 17833 9781 17867
rect 9815 17864 9827 17867
rect 15194 17864 15200 17876
rect 9815 17836 15200 17864
rect 9815 17833 9827 17836
rect 9769 17827 9827 17833
rect 4157 17731 4215 17737
rect 3068 17700 3924 17728
rect 3068 17669 3096 17700
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 3283 17632 3832 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 3804 17533 3832 17632
rect 3896 17592 3924 17700
rect 4157 17697 4169 17731
rect 4203 17728 4215 17731
rect 4798 17728 4804 17740
rect 4203 17700 4804 17728
rect 4203 17697 4215 17700
rect 4157 17691 4215 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 7374 17660 7380 17672
rect 4028 17632 7380 17660
rect 4028 17620 4034 17632
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 8202 17660 8208 17672
rect 8163 17632 8208 17660
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 8536 17632 8953 17660
rect 8536 17620 8542 17632
rect 8941 17629 8953 17632
rect 8987 17660 8999 17663
rect 9784 17660 9812 17827
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 22370 17864 22376 17876
rect 22331 17836 22376 17864
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 8987 17632 9812 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 23474 17620 23480 17672
rect 23532 17669 23538 17672
rect 23532 17660 23544 17669
rect 23753 17663 23811 17669
rect 23532 17632 23577 17660
rect 23532 17623 23544 17632
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 38102 17660 38108 17672
rect 23799 17632 24532 17660
rect 38063 17632 38108 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 23532 17620 23538 17623
rect 3896 17564 4752 17592
rect 3789 17527 3847 17533
rect 3789 17493 3801 17527
rect 3835 17524 3847 17527
rect 4614 17524 4620 17536
rect 3835 17496 4620 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 4724 17524 4752 17564
rect 4890 17524 4896 17536
rect 4724 17496 4896 17524
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 4948 17496 9137 17524
rect 4948 17484 4954 17496
rect 9125 17493 9137 17496
rect 9171 17524 9183 17527
rect 12434 17524 12440 17536
rect 9171 17496 12440 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 24504 17533 24532 17632
rect 38102 17620 38108 17632
rect 38160 17620 38166 17672
rect 24489 17527 24547 17533
rect 24489 17493 24501 17527
rect 24535 17524 24547 17527
rect 25774 17524 25780 17536
rect 24535 17496 25780 17524
rect 24535 17493 24547 17496
rect 24489 17487 24547 17493
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8478 17320 8484 17332
rect 8439 17292 8484 17320
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 26602 17280 26608 17332
rect 26660 17320 26666 17332
rect 34330 17320 34336 17332
rect 26660 17292 34336 17320
rect 26660 17280 26666 17292
rect 34330 17280 34336 17292
rect 34388 17280 34394 17332
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7653 17187 7711 17193
rect 7653 17184 7665 17187
rect 7432 17156 7665 17184
rect 7432 17144 7438 17156
rect 7653 17153 7665 17156
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 8496 17184 8524 17280
rect 17678 17252 17684 17264
rect 12728 17224 17684 17252
rect 7883 17156 8524 17184
rect 12253 17187 12311 17193
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 7558 17116 7564 17128
rect 7519 17088 7564 17116
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 7745 17119 7803 17125
rect 7745 17085 7757 17119
rect 7791 17085 7803 17119
rect 12268 17116 12296 17147
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12728 17184 12756 17224
rect 17678 17212 17684 17224
rect 17736 17212 17742 17264
rect 12492 17156 12756 17184
rect 12492 17144 12498 17156
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12860 17156 13185 17184
rect 12860 17144 12866 17156
rect 13173 17153 13185 17156
rect 13219 17184 13231 17187
rect 17770 17184 17776 17196
rect 13219 17156 17776 17184
rect 13219 17153 13231 17156
rect 13173 17147 13231 17153
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 33873 17187 33931 17193
rect 33873 17153 33885 17187
rect 33919 17184 33931 17187
rect 33962 17184 33968 17196
rect 33919 17156 33968 17184
rect 33919 17153 33931 17156
rect 33873 17147 33931 17153
rect 33962 17144 33968 17156
rect 34020 17144 34026 17196
rect 12342 17116 12348 17128
rect 12268 17088 12348 17116
rect 7745 17079 7803 17085
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 7760 17048 7788 17079
rect 12342 17076 12348 17088
rect 12400 17116 12406 17128
rect 12989 17119 13047 17125
rect 12989 17116 13001 17119
rect 12400 17088 13001 17116
rect 12400 17076 12406 17088
rect 12989 17085 13001 17088
rect 13035 17085 13047 17119
rect 12989 17079 13047 17085
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17085 13415 17119
rect 34146 17116 34152 17128
rect 34107 17088 34152 17116
rect 13357 17079 13415 17085
rect 7064 17020 7788 17048
rect 7064 17008 7070 17020
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 13372 17048 13400 17079
rect 34146 17076 34152 17088
rect 34204 17076 34210 17128
rect 12584 17020 13400 17048
rect 12584 17008 12590 17020
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 7377 16983 7435 16989
rect 7377 16980 7389 16983
rect 7340 16952 7389 16980
rect 7340 16940 7346 16952
rect 7377 16949 7389 16952
rect 7423 16949 7435 16983
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 7377 16943 7435 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 7006 16776 7012 16788
rect 4856 16748 7012 16776
rect 4856 16736 4862 16748
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 12802 16776 12808 16788
rect 12483 16748 12808 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 17865 16711 17923 16717
rect 17865 16677 17877 16711
rect 17911 16708 17923 16711
rect 18690 16708 18696 16720
rect 17911 16680 18696 16708
rect 17911 16677 17923 16680
rect 17865 16671 17923 16677
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 31665 16643 31723 16649
rect 17828 16612 17908 16640
rect 17828 16600 17834 16612
rect 12250 16572 12256 16584
rect 12211 16544 12256 16572
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 17678 16572 17684 16584
rect 12584 16544 12629 16572
rect 17639 16544 17684 16572
rect 12584 16532 12590 16544
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 17880 16581 17908 16612
rect 31665 16609 31677 16643
rect 31711 16640 31723 16643
rect 31938 16640 31944 16652
rect 31711 16612 31944 16640
rect 31711 16609 31723 16612
rect 31665 16603 31723 16609
rect 31938 16600 31944 16612
rect 31996 16600 32002 16652
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 31386 16572 31392 16584
rect 31347 16544 31392 16572
rect 17865 16535 17923 16541
rect 31386 16532 31392 16544
rect 31444 16532 31450 16584
rect 7190 16504 7196 16516
rect 7151 16476 7196 16504
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6993 16439 7051 16445
rect 6993 16405 7005 16439
rect 7039 16436 7051 16439
rect 8202 16436 8208 16448
rect 7039 16408 8208 16436
rect 7039 16405 7051 16408
rect 6993 16399 7051 16405
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 37553 16439 37611 16445
rect 37553 16405 37565 16439
rect 37599 16436 37611 16439
rect 37734 16436 37740 16448
rect 37599 16408 37740 16436
rect 37599 16405 37611 16408
rect 37553 16399 37611 16405
rect 37734 16396 37740 16408
rect 37792 16396 37798 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 30558 16192 30564 16244
rect 30616 16232 30622 16244
rect 30653 16235 30711 16241
rect 30653 16232 30665 16235
rect 30616 16204 30665 16232
rect 30616 16192 30622 16204
rect 30653 16201 30665 16204
rect 30699 16201 30711 16235
rect 30653 16195 30711 16201
rect 33965 16235 34023 16241
rect 33965 16201 33977 16235
rect 34011 16232 34023 16235
rect 34146 16232 34152 16244
rect 34011 16204 34152 16232
rect 34011 16201 34023 16204
rect 33965 16195 34023 16201
rect 34146 16192 34152 16204
rect 34204 16192 34210 16244
rect 34422 16232 34428 16244
rect 34383 16204 34428 16232
rect 34422 16192 34428 16204
rect 34480 16192 34486 16244
rect 37826 16232 37832 16244
rect 37787 16204 37832 16232
rect 37826 16192 37832 16204
rect 37884 16192 37890 16244
rect 4890 16164 4896 16176
rect 4264 16136 4896 16164
rect 4264 16105 4292 16136
rect 4890 16124 4896 16136
rect 4948 16124 4954 16176
rect 30009 16167 30067 16173
rect 30009 16133 30021 16167
rect 30055 16164 30067 16167
rect 30374 16164 30380 16176
rect 30055 16136 30380 16164
rect 30055 16133 30067 16136
rect 30009 16127 30067 16133
rect 30374 16124 30380 16136
rect 30432 16124 30438 16176
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 4249 16059 4307 16065
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 6822 16096 6828 16108
rect 4479 16068 6828 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 18874 16096 18880 16108
rect 18835 16068 18880 16096
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 20162 16096 20168 16108
rect 19015 16068 20168 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 28994 16056 29000 16108
rect 29052 16096 29058 16108
rect 29825 16099 29883 16105
rect 29825 16096 29837 16099
rect 29052 16068 29837 16096
rect 29052 16056 29058 16068
rect 29825 16065 29837 16068
rect 29871 16065 29883 16099
rect 30558 16096 30564 16108
rect 30519 16068 30564 16096
rect 29825 16059 29883 16065
rect 30558 16056 30564 16068
rect 30616 16056 30622 16108
rect 33410 16056 33416 16108
rect 33468 16096 33474 16108
rect 34333 16099 34391 16105
rect 34333 16096 34345 16099
rect 33468 16068 34345 16096
rect 33468 16056 33474 16068
rect 34333 16065 34345 16068
rect 34379 16065 34391 16099
rect 37734 16096 37740 16108
rect 37647 16068 37740 16096
rect 34333 16059 34391 16065
rect 37734 16056 37740 16068
rect 37792 16096 37798 16108
rect 38930 16096 38936 16108
rect 37792 16068 38936 16096
rect 37792 16056 37798 16068
rect 38930 16056 38936 16068
rect 38988 16056 38994 16108
rect 31938 15988 31944 16040
rect 31996 16028 32002 16040
rect 34609 16031 34667 16037
rect 34609 16028 34621 16031
rect 31996 16000 34621 16028
rect 31996 15988 32002 16000
rect 34609 15997 34621 16000
rect 34655 16028 34667 16031
rect 37918 16028 37924 16040
rect 34655 16000 37924 16028
rect 34655 15997 34667 16000
rect 34609 15991 34667 15997
rect 37918 15988 37924 16000
rect 37976 15988 37982 16040
rect 3970 15852 3976 15904
rect 4028 15892 4034 15904
rect 4433 15895 4491 15901
rect 4433 15892 4445 15895
rect 4028 15864 4445 15892
rect 4028 15852 4034 15864
rect 4433 15861 4445 15864
rect 4479 15861 4491 15895
rect 18506 15892 18512 15904
rect 18467 15864 18512 15892
rect 4433 15855 4491 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 33410 15892 33416 15904
rect 33371 15864 33416 15892
rect 33410 15852 33416 15864
rect 33468 15852 33474 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 4157 15691 4215 15697
rect 4157 15657 4169 15691
rect 4203 15688 4215 15691
rect 4614 15688 4620 15700
rect 4203 15660 4620 15688
rect 4203 15657 4215 15660
rect 4157 15651 4215 15657
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 12437 15691 12495 15697
rect 12437 15657 12449 15691
rect 12483 15688 12495 15691
rect 12526 15688 12532 15700
rect 12483 15660 12532 15688
rect 12483 15657 12495 15660
rect 12437 15651 12495 15657
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 20162 15648 20168 15700
rect 20220 15688 20226 15700
rect 20625 15691 20683 15697
rect 20625 15688 20637 15691
rect 20220 15660 20637 15688
rect 20220 15648 20226 15660
rect 20625 15657 20637 15660
rect 20671 15657 20683 15691
rect 20625 15651 20683 15657
rect 27157 15691 27215 15697
rect 27157 15657 27169 15691
rect 27203 15688 27215 15691
rect 27246 15688 27252 15700
rect 27203 15660 27252 15688
rect 27203 15657 27215 15660
rect 27157 15651 27215 15657
rect 27246 15648 27252 15660
rect 27304 15648 27310 15700
rect 30653 15691 30711 15697
rect 30653 15657 30665 15691
rect 30699 15688 30711 15691
rect 31386 15688 31392 15700
rect 30699 15660 31392 15688
rect 30699 15657 30711 15660
rect 30653 15651 30711 15657
rect 31386 15648 31392 15660
rect 31444 15648 31450 15700
rect 32214 15688 32220 15700
rect 31680 15660 32220 15688
rect 31680 15629 31708 15660
rect 32214 15648 32220 15660
rect 32272 15688 32278 15700
rect 32401 15691 32459 15697
rect 32401 15688 32413 15691
rect 32272 15660 32413 15688
rect 32272 15648 32278 15660
rect 32401 15657 32413 15660
rect 32447 15657 32459 15691
rect 34790 15688 34796 15700
rect 34751 15660 34796 15688
rect 32401 15651 32459 15657
rect 34790 15648 34796 15660
rect 34848 15648 34854 15700
rect 37918 15688 37924 15700
rect 37879 15660 37924 15688
rect 37918 15648 37924 15660
rect 37976 15648 37982 15700
rect 31665 15623 31723 15629
rect 31665 15589 31677 15623
rect 31711 15589 31723 15623
rect 31665 15583 31723 15589
rect 18506 15512 18512 15564
rect 18564 15552 18570 15564
rect 31938 15552 31944 15564
rect 18564 15524 19380 15552
rect 31899 15524 31944 15552
rect 18564 15512 18570 15524
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 4249 15447 4307 15453
rect 10520 15456 11069 15484
rect 3786 15348 3792 15360
rect 3747 15320 3792 15348
rect 3786 15308 3792 15320
rect 3844 15308 3850 15360
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 10042 15348 10048 15360
rect 6972 15320 10048 15348
rect 6972 15308 6978 15320
rect 10042 15308 10048 15320
rect 10100 15348 10106 15360
rect 10520 15357 10548 15456
rect 11057 15453 11069 15456
rect 11103 15484 11115 15487
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 11103 15456 18613 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 18601 15453 18613 15456
rect 18647 15484 18659 15487
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18647 15456 19257 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19352 15484 19380 15524
rect 31938 15512 31944 15524
rect 31996 15512 32002 15564
rect 19501 15487 19559 15493
rect 19501 15484 19513 15487
rect 19352 15456 19513 15484
rect 19245 15447 19303 15453
rect 19501 15453 19513 15456
rect 19547 15453 19559 15487
rect 25774 15484 25780 15496
rect 25687 15456 25780 15484
rect 19501 15447 19559 15453
rect 25774 15444 25780 15456
rect 25832 15484 25838 15496
rect 27617 15487 27675 15493
rect 27617 15484 27629 15487
rect 25832 15456 27629 15484
rect 25832 15444 25838 15456
rect 27617 15453 27629 15456
rect 27663 15484 27675 15487
rect 28258 15484 28264 15496
rect 27663 15456 28264 15484
rect 27663 15453 27675 15456
rect 27617 15447 27675 15453
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 29178 15444 29184 15496
rect 29236 15484 29242 15496
rect 30469 15487 30527 15493
rect 30469 15484 30481 15487
rect 29236 15456 30481 15484
rect 29236 15444 29242 15456
rect 30469 15453 30481 15456
rect 30515 15484 30527 15487
rect 31956 15484 31984 15512
rect 30515 15456 31984 15484
rect 30515 15453 30527 15456
rect 30469 15447 30527 15453
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34756 15456 34897 15484
rect 34756 15444 34762 15456
rect 34885 15453 34897 15456
rect 34931 15484 34943 15487
rect 35345 15487 35403 15493
rect 35345 15484 35357 15487
rect 34931 15456 35357 15484
rect 34931 15453 34943 15456
rect 34885 15447 34943 15453
rect 35345 15453 35357 15456
rect 35391 15453 35403 15487
rect 38010 15484 38016 15496
rect 37971 15456 38016 15484
rect 35345 15447 35403 15453
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 11324 15419 11382 15425
rect 11324 15385 11336 15419
rect 11370 15416 11382 15419
rect 12066 15416 12072 15428
rect 11370 15388 12072 15416
rect 11370 15385 11382 15388
rect 11324 15379 11382 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 18782 15376 18788 15428
rect 18840 15416 18846 15428
rect 26050 15425 26056 15428
rect 26044 15416 26056 15425
rect 18840 15388 22094 15416
rect 26011 15388 26056 15416
rect 18840 15376 18846 15388
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10100 15320 10517 15348
rect 10100 15308 10106 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 22066 15348 22094 15388
rect 26044 15379 26056 15388
rect 26050 15376 26056 15379
rect 26108 15376 26114 15428
rect 29733 15419 29791 15425
rect 29733 15416 29745 15419
rect 27080 15388 29745 15416
rect 27080 15348 27108 15388
rect 29733 15385 29745 15388
rect 29779 15416 29791 15419
rect 30285 15419 30343 15425
rect 30285 15416 30297 15419
rect 29779 15388 30297 15416
rect 29779 15385 29791 15388
rect 29733 15379 29791 15385
rect 30285 15385 30297 15388
rect 30331 15385 30343 15419
rect 36446 15416 36452 15428
rect 36407 15388 36452 15416
rect 30285 15379 30343 15385
rect 36446 15376 36452 15388
rect 36504 15416 36510 15428
rect 37185 15419 37243 15425
rect 37185 15416 37197 15419
rect 36504 15388 37197 15416
rect 36504 15376 36510 15388
rect 37185 15385 37197 15388
rect 37231 15385 37243 15419
rect 37185 15379 37243 15385
rect 31478 15348 31484 15360
rect 22066 15320 27108 15348
rect 31439 15320 31484 15348
rect 10505 15311 10563 15317
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 36630 15308 36636 15360
rect 36688 15348 36694 15360
rect 37093 15351 37151 15357
rect 37093 15348 37105 15351
rect 36688 15320 37105 15348
rect 36688 15308 36694 15320
rect 37093 15317 37105 15320
rect 37139 15317 37151 15351
rect 37093 15311 37151 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 7285 15147 7343 15153
rect 7285 15113 7297 15147
rect 7331 15144 7343 15147
rect 7558 15144 7564 15156
rect 7331 15116 7564 15144
rect 7331 15113 7343 15116
rect 7285 15107 7343 15113
rect 7558 15104 7564 15116
rect 7616 15104 7622 15156
rect 17126 15144 17132 15156
rect 17087 15116 17132 15144
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 23198 15144 23204 15156
rect 23159 15116 23204 15144
rect 23198 15104 23204 15116
rect 23256 15104 23262 15156
rect 28261 15147 28319 15153
rect 28261 15113 28273 15147
rect 28307 15144 28319 15147
rect 28994 15144 29000 15156
rect 28307 15116 29000 15144
rect 28307 15113 28319 15116
rect 28261 15107 28319 15113
rect 28994 15104 29000 15116
rect 29052 15104 29058 15156
rect 29641 15147 29699 15153
rect 29641 15113 29653 15147
rect 29687 15144 29699 15147
rect 30558 15144 30564 15156
rect 29687 15116 30564 15144
rect 29687 15113 29699 15116
rect 29641 15107 29699 15113
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 36538 15104 36544 15156
rect 36596 15144 36602 15156
rect 36633 15147 36691 15153
rect 36633 15144 36645 15147
rect 36596 15116 36645 15144
rect 36596 15104 36602 15116
rect 36633 15113 36645 15116
rect 36679 15113 36691 15147
rect 38010 15144 38016 15156
rect 37971 15116 38016 15144
rect 36633 15107 36691 15113
rect 38010 15104 38016 15116
rect 38068 15104 38074 15156
rect 21910 15036 21916 15088
rect 21968 15076 21974 15088
rect 22373 15079 22431 15085
rect 22373 15076 22385 15079
rect 21968 15048 22385 15076
rect 21968 15036 21974 15048
rect 22373 15045 22385 15048
rect 22419 15045 22431 15079
rect 22373 15039 22431 15045
rect 28721 15079 28779 15085
rect 28721 15045 28733 15079
rect 28767 15076 28779 15079
rect 29178 15076 29184 15088
rect 28767 15048 29184 15076
rect 28767 15045 28779 15048
rect 28721 15039 28779 15045
rect 29178 15036 29184 15048
rect 29236 15036 29242 15088
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 7190 15008 7196 15020
rect 4120 14980 7196 15008
rect 4120 14968 4126 14980
rect 7190 14968 7196 14980
rect 7248 15008 7254 15020
rect 7469 15011 7527 15017
rect 7469 15008 7481 15011
rect 7248 14980 7481 15008
rect 7248 14968 7254 14980
rect 7469 14977 7481 14980
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 16942 14968 16948 15020
rect 17000 15008 17006 15020
rect 17221 15011 17279 15017
rect 17221 15008 17233 15011
rect 17000 14980 17233 15008
rect 17000 14968 17006 14980
rect 17221 14977 17233 14980
rect 17267 14977 17279 15011
rect 22554 15008 22560 15020
rect 22515 14980 22560 15008
rect 17221 14971 17279 14977
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 31726 14980 35894 15008
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 8294 14940 8300 14952
rect 7699 14912 8300 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 23658 14832 23664 14884
rect 23716 14872 23722 14884
rect 23753 14875 23811 14881
rect 23753 14872 23765 14875
rect 23716 14844 23765 14872
rect 23716 14832 23722 14844
rect 23753 14841 23765 14844
rect 23799 14841 23811 14875
rect 23753 14835 23811 14841
rect 27801 14875 27859 14881
rect 27801 14841 27813 14875
rect 27847 14872 27859 14875
rect 28445 14875 28503 14881
rect 28445 14872 28457 14875
rect 27847 14844 28457 14872
rect 27847 14841 27859 14844
rect 27801 14835 27859 14841
rect 28445 14841 28457 14844
rect 28491 14872 28503 14875
rect 28534 14872 28540 14884
rect 28491 14844 28540 14872
rect 28491 14841 28503 14844
rect 28445 14835 28503 14841
rect 28534 14832 28540 14844
rect 28592 14832 28598 14884
rect 29454 14872 29460 14884
rect 29415 14844 29460 14872
rect 29454 14832 29460 14844
rect 29512 14832 29518 14884
rect 14642 14804 14648 14816
rect 14603 14776 14648 14804
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 31726 14804 31754 14980
rect 35866 14872 35894 14980
rect 35986 14968 35992 15020
rect 36044 15008 36050 15020
rect 36541 15011 36599 15017
rect 36541 15008 36553 15011
rect 36044 14980 36553 15008
rect 36044 14968 36050 14980
rect 36541 14977 36553 14980
rect 36587 14977 36599 15011
rect 36541 14971 36599 14977
rect 37277 15011 37335 15017
rect 37277 14977 37289 15011
rect 37323 15008 37335 15011
rect 37366 15008 37372 15020
rect 37323 14980 37372 15008
rect 37323 14977 37335 14980
rect 37277 14971 37335 14977
rect 37366 14968 37372 14980
rect 37424 14968 37430 15020
rect 37461 14875 37519 14881
rect 37461 14872 37473 14875
rect 35866 14844 37473 14872
rect 37461 14841 37473 14844
rect 37507 14841 37519 14875
rect 37461 14835 37519 14841
rect 35986 14804 35992 14816
rect 20312 14776 31754 14804
rect 35947 14776 35992 14804
rect 20312 14764 20318 14776
rect 35986 14764 35992 14776
rect 36044 14764 36050 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 13780 14572 14289 14600
rect 13780 14560 13786 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14792 14572 15117 14600
rect 14792 14560 14798 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 34698 14600 34704 14612
rect 15795 14572 34704 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 6880 14436 7604 14464
rect 6880 14424 6886 14436
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7576 14405 7604 14436
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 8294 14396 8300 14408
rect 7791 14368 8300 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15764 14396 15792 14563
rect 34698 14560 34704 14572
rect 34756 14560 34762 14612
rect 23845 14535 23903 14541
rect 22066 14504 23336 14532
rect 15838 14424 15844 14476
rect 15896 14464 15902 14476
rect 22066 14464 22094 14504
rect 15896 14436 22094 14464
rect 23109 14467 23167 14473
rect 15896 14424 15902 14436
rect 23109 14433 23121 14467
rect 23155 14464 23167 14467
rect 23198 14464 23204 14476
rect 23155 14436 23204 14464
rect 23155 14433 23167 14436
rect 23109 14427 23167 14433
rect 23198 14424 23204 14436
rect 23256 14424 23262 14476
rect 23308 14464 23336 14504
rect 23845 14501 23857 14535
rect 23891 14532 23903 14535
rect 24854 14532 24860 14544
rect 23891 14504 24860 14532
rect 23891 14501 23903 14504
rect 23845 14495 23903 14501
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 28994 14464 29000 14476
rect 23308 14436 29000 14464
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 36722 14424 36728 14476
rect 36780 14464 36786 14476
rect 37553 14467 37611 14473
rect 37553 14464 37565 14467
rect 36780 14436 37565 14464
rect 36780 14424 36786 14436
rect 37553 14433 37565 14436
rect 37599 14433 37611 14467
rect 37553 14427 37611 14433
rect 15059 14368 15792 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 22462 14356 22468 14408
rect 22520 14396 22526 14408
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22520 14368 22845 14396
rect 22520 14356 22526 14368
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 23658 14396 23664 14408
rect 23619 14368 23664 14396
rect 22833 14359 22891 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 24118 14356 24124 14408
rect 24176 14396 24182 14408
rect 29454 14396 29460 14408
rect 24176 14368 29460 14396
rect 24176 14356 24182 14368
rect 29454 14356 29460 14368
rect 29512 14396 29518 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 29512 14368 29561 14396
rect 29512 14356 29518 14368
rect 29549 14365 29561 14368
rect 29595 14365 29607 14399
rect 29549 14359 29607 14365
rect 36817 14399 36875 14405
rect 36817 14365 36829 14399
rect 36863 14396 36875 14399
rect 37274 14396 37280 14408
rect 36863 14368 37280 14396
rect 36863 14365 36875 14368
rect 36817 14359 36875 14365
rect 37274 14356 37280 14368
rect 37332 14356 37338 14408
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 14829 14331 14887 14337
rect 14829 14328 14841 14331
rect 14700 14300 14841 14328
rect 14700 14288 14706 14300
rect 14829 14297 14841 14300
rect 14875 14297 14887 14331
rect 14829 14291 14887 14297
rect 18414 14288 18420 14340
rect 18472 14328 18478 14340
rect 31386 14328 31392 14340
rect 18472 14300 31392 14328
rect 18472 14288 18478 14300
rect 31386 14288 31392 14300
rect 31444 14288 31450 14340
rect 7101 14263 7159 14269
rect 7101 14229 7113 14263
rect 7147 14260 7159 14263
rect 7190 14260 7196 14272
rect 7147 14232 7196 14260
rect 7147 14229 7159 14232
rect 7101 14223 7159 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 24397 14263 24455 14269
rect 24397 14260 24409 14263
rect 24360 14232 24409 14260
rect 24360 14220 24366 14232
rect 24397 14229 24409 14232
rect 24443 14229 24455 14263
rect 24397 14223 24455 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15838 14056 15844 14068
rect 15151 14028 15844 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 25593 14059 25651 14065
rect 25593 14056 25605 14059
rect 16172 14028 25605 14056
rect 16172 14016 16178 14028
rect 25593 14025 25605 14028
rect 25639 14025 25651 14059
rect 26326 14056 26332 14068
rect 25593 14019 25651 14025
rect 25700 14028 26332 14056
rect 4525 13991 4583 13997
rect 4525 13988 4537 13991
rect 2700 13960 4537 13988
rect 2700 13929 2728 13960
rect 4525 13957 4537 13960
rect 4571 13988 4583 13991
rect 6914 13988 6920 14000
rect 4571 13960 6920 13988
rect 4571 13957 4583 13960
rect 4525 13951 4583 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 14185 13991 14243 13997
rect 14185 13957 14197 13991
rect 14231 13988 14243 13991
rect 14274 13988 14280 14000
rect 14231 13960 14280 13988
rect 14231 13957 14243 13960
rect 14185 13951 14243 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 15930 13948 15936 14000
rect 15988 13988 15994 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 15988 13960 17049 13988
rect 15988 13948 15994 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 17954 13948 17960 14000
rect 18012 13988 18018 14000
rect 24118 13988 24124 14000
rect 18012 13960 24124 13988
rect 18012 13948 18018 13960
rect 24118 13948 24124 13960
rect 24176 13948 24182 14000
rect 24302 13988 24308 14000
rect 24263 13960 24308 13988
rect 24302 13948 24308 13960
rect 24360 13948 24366 14000
rect 24489 13991 24547 13997
rect 24489 13957 24501 13991
rect 24535 13988 24547 13991
rect 25406 13988 25412 14000
rect 24535 13960 25412 13988
rect 24535 13957 24547 13960
rect 24489 13951 24547 13957
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 25700 13997 25728 14028
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 31386 14056 31392 14068
rect 31347 14028 31392 14056
rect 31386 14016 31392 14028
rect 31444 14016 31450 14068
rect 25685 13991 25743 13997
rect 25685 13957 25697 13991
rect 25731 13957 25743 13991
rect 31478 13988 31484 14000
rect 31439 13960 31484 13988
rect 25685 13951 25743 13957
rect 31478 13948 31484 13960
rect 31536 13948 31542 14000
rect 37921 13991 37979 13997
rect 37921 13957 37933 13991
rect 37967 13988 37979 13991
rect 38286 13988 38292 14000
rect 37967 13960 38292 13988
rect 37967 13957 37979 13960
rect 37921 13951 37979 13957
rect 38286 13948 38292 13960
rect 38344 13948 38350 14000
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2952 13923 3010 13929
rect 2952 13889 2964 13923
rect 2998 13920 3010 13923
rect 3786 13920 3792 13932
rect 2998 13892 3792 13920
rect 2998 13889 3010 13892
rect 2952 13883 3010 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 13998 13920 14004 13932
rect 13959 13892 14004 13920
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 17184 13892 17233 13920
rect 17184 13880 17190 13892
rect 17221 13889 17233 13892
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 23566 13880 23572 13932
rect 23624 13920 23630 13932
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 23624 13892 23765 13920
rect 23624 13880 23630 13892
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 37734 13920 37740 13932
rect 37695 13892 37740 13920
rect 23753 13883 23811 13889
rect 37734 13880 37740 13892
rect 37792 13880 37798 13932
rect 14642 13852 14648 13864
rect 14603 13824 14648 13852
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15562 13812 15568 13864
rect 15620 13852 15626 13864
rect 23477 13855 23535 13861
rect 23477 13852 23489 13855
rect 15620 13824 23489 13852
rect 15620 13812 15626 13824
rect 23477 13821 23489 13824
rect 23523 13821 23535 13855
rect 23477 13815 23535 13821
rect 13722 13744 13728 13796
rect 13780 13784 13786 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 13780 13756 14933 13784
rect 13780 13744 13786 13756
rect 14921 13753 14933 13756
rect 14967 13753 14979 13787
rect 14921 13747 14979 13753
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22612 13484 22845 13512
rect 22612 13472 22618 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 23566 13472 23572 13524
rect 23624 13512 23630 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 23624 13484 24409 13512
rect 23624 13472 23630 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 36722 13512 36728 13524
rect 24397 13475 24455 13481
rect 31726 13484 36728 13512
rect 31726 13444 31754 13484
rect 36722 13472 36728 13484
rect 36780 13472 36786 13524
rect 23308 13416 31754 13444
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 23308 13385 23336 13416
rect 23293 13379 23351 13385
rect 11204 13348 19334 13376
rect 11204 13336 11210 13348
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 19306 13308 19334 13348
rect 23293 13345 23305 13379
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 23658 13376 23664 13388
rect 23523 13348 23664 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 10744 13280 17172 13308
rect 19306 13280 23520 13308
rect 10744 13268 10750 13280
rect 13262 13132 13268 13184
rect 13320 13172 13326 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 13320 13144 14473 13172
rect 13320 13132 13326 13144
rect 14461 13141 14473 13144
rect 14507 13172 14519 13175
rect 14642 13172 14648 13184
rect 14507 13144 14648 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 17144 13172 17172 13280
rect 22278 13240 22284 13252
rect 22239 13212 22284 13240
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 23198 13240 23204 13252
rect 23159 13212 23204 13240
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 23492 13240 23520 13280
rect 23566 13268 23572 13320
rect 23624 13308 23630 13320
rect 33686 13308 33692 13320
rect 23624 13280 33692 13308
rect 23624 13268 23630 13280
rect 33686 13268 33692 13280
rect 33744 13268 33750 13320
rect 31846 13240 31852 13252
rect 23492 13212 31852 13240
rect 31846 13200 31852 13212
rect 31904 13200 31910 13252
rect 23106 13172 23112 13184
rect 17144 13144 23112 13172
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 37553 13175 37611 13181
rect 37553 13141 37565 13175
rect 37599 13172 37611 13175
rect 37734 13172 37740 13184
rect 37599 13144 37740 13172
rect 37599 13141 37611 13144
rect 37553 13135 37611 13141
rect 37734 13132 37740 13144
rect 37792 13172 37798 13184
rect 38470 13172 38476 13184
rect 37792 13144 38476 13172
rect 37792 13132 37798 13144
rect 38470 13132 38476 13144
rect 38528 13132 38534 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 23474 12968 23480 12980
rect 20588 12940 23480 12968
rect 20588 12928 20594 12940
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 23658 12968 23664 12980
rect 23619 12940 23664 12968
rect 23658 12928 23664 12940
rect 23716 12968 23722 12980
rect 23842 12968 23848 12980
rect 23716 12940 23848 12968
rect 23716 12928 23722 12940
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 8757 12903 8815 12909
rect 8757 12900 8769 12903
rect 6932 12872 8769 12900
rect 6932 12844 6960 12872
rect 8757 12869 8769 12872
rect 8803 12869 8815 12903
rect 8757 12863 8815 12869
rect 13265 12903 13323 12909
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 13906 12900 13912 12912
rect 13311 12872 13912 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 28994 12860 29000 12912
rect 29052 12900 29058 12912
rect 34057 12903 34115 12909
rect 34057 12900 34069 12903
rect 29052 12872 34069 12900
rect 29052 12860 29058 12872
rect 6914 12832 6920 12844
rect 6875 12804 6920 12832
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7190 12841 7196 12844
rect 7184 12832 7196 12841
rect 7151 12804 7196 12832
rect 7184 12795 7196 12804
rect 7190 12792 7196 12795
rect 7248 12792 7254 12844
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13170 12832 13176 12844
rect 13127 12804 13176 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 25961 12835 26019 12841
rect 25961 12801 25973 12835
rect 26007 12832 26019 12835
rect 27522 12832 27528 12844
rect 26007 12804 27528 12832
rect 26007 12801 26019 12804
rect 25961 12795 26019 12801
rect 27522 12792 27528 12804
rect 27580 12792 27586 12844
rect 32122 12832 32128 12844
rect 32083 12804 32128 12832
rect 32122 12792 32128 12804
rect 32180 12792 32186 12844
rect 33428 12841 33456 12872
rect 34057 12869 34069 12872
rect 34103 12869 34115 12903
rect 34057 12863 34115 12869
rect 33413 12835 33471 12841
rect 33413 12801 33425 12835
rect 33459 12801 33471 12835
rect 33413 12795 33471 12801
rect 32398 12764 32404 12776
rect 32359 12736 32404 12764
rect 32398 12724 32404 12736
rect 32456 12724 32462 12776
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 25777 12699 25835 12705
rect 25777 12696 25789 12699
rect 9824 12668 25789 12696
rect 9824 12656 9830 12668
rect 25777 12665 25789 12668
rect 25823 12665 25835 12699
rect 25777 12659 25835 12665
rect 19794 12628 19800 12640
rect 19755 12600 19800 12628
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 33597 12631 33655 12637
rect 33597 12597 33609 12631
rect 33643 12628 33655 12631
rect 33686 12628 33692 12640
rect 33643 12600 33692 12628
rect 33643 12597 33655 12600
rect 33597 12591 33655 12597
rect 33686 12588 33692 12600
rect 33744 12588 33750 12640
rect 38102 12628 38108 12640
rect 38063 12600 38108 12628
rect 38102 12588 38108 12600
rect 38160 12588 38166 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 20714 12424 20720 12436
rect 19567 12396 20720 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 22646 12424 22652 12436
rect 22066 12396 22652 12424
rect 4433 12359 4491 12365
rect 4433 12325 4445 12359
rect 4479 12356 4491 12359
rect 4614 12356 4620 12368
rect 4479 12328 4620 12356
rect 4479 12325 4491 12328
rect 4433 12319 4491 12325
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 9677 12359 9735 12365
rect 9677 12325 9689 12359
rect 9723 12356 9735 12359
rect 11698 12356 11704 12368
rect 9723 12328 11704 12356
rect 9723 12325 9735 12328
rect 9677 12319 9735 12325
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 20625 12359 20683 12365
rect 20625 12325 20637 12359
rect 20671 12356 20683 12359
rect 21913 12359 21971 12365
rect 21913 12356 21925 12359
rect 20671 12328 21925 12356
rect 20671 12325 20683 12328
rect 20625 12319 20683 12325
rect 21913 12325 21925 12328
rect 21959 12356 21971 12359
rect 22066 12356 22094 12396
rect 22646 12384 22652 12396
rect 22704 12384 22710 12436
rect 21959 12328 22094 12356
rect 21959 12325 21971 12328
rect 21913 12319 21971 12325
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 16298 12288 16304 12300
rect 7800 12260 16304 12288
rect 7800 12248 7806 12260
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 9539 12192 9674 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 4249 12155 4307 12161
rect 4249 12121 4261 12155
rect 4295 12152 4307 12155
rect 4706 12152 4712 12164
rect 4295 12124 4712 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 9646 12084 9674 12192
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 31021 12223 31079 12229
rect 31021 12220 31033 12223
rect 11480 12192 31033 12220
rect 11480 12180 11486 12192
rect 31021 12189 31033 12192
rect 31067 12189 31079 12223
rect 31021 12183 31079 12189
rect 19245 12155 19303 12161
rect 19245 12121 19257 12155
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 10229 12087 10287 12093
rect 10229 12084 10241 12087
rect 9646 12056 10241 12084
rect 10229 12053 10241 12056
rect 10275 12084 10287 12087
rect 14550 12084 14556 12096
rect 10275 12056 14556 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18288 12056 18613 12084
rect 18288 12044 18294 12056
rect 18601 12053 18613 12056
rect 18647 12084 18659 12087
rect 19260 12084 19288 12115
rect 19334 12112 19340 12164
rect 19392 12152 19398 12164
rect 19429 12155 19487 12161
rect 19429 12152 19441 12155
rect 19392 12124 19441 12152
rect 19392 12112 19398 12124
rect 19429 12121 19441 12124
rect 19475 12152 19487 12155
rect 19794 12152 19800 12164
rect 19475 12124 19800 12152
rect 19475 12121 19487 12124
rect 19429 12115 19487 12121
rect 19794 12112 19800 12124
rect 19852 12152 19858 12164
rect 20901 12155 20959 12161
rect 20901 12152 20913 12155
rect 19852 12124 20913 12152
rect 19852 12112 19858 12124
rect 20901 12121 20913 12124
rect 20947 12152 20959 12155
rect 21453 12155 21511 12161
rect 21453 12152 21465 12155
rect 20947 12124 21465 12152
rect 20947 12121 20959 12124
rect 20901 12115 20959 12121
rect 21453 12121 21465 12124
rect 21499 12152 21511 12155
rect 23842 12152 23848 12164
rect 21499 12124 23848 12152
rect 21499 12121 21511 12124
rect 21453 12115 21511 12121
rect 23842 12112 23848 12124
rect 23900 12152 23906 12164
rect 31386 12152 31392 12164
rect 23900 12124 31064 12152
rect 31347 12124 31392 12152
rect 23900 12112 23906 12124
rect 20438 12084 20444 12096
rect 18647 12056 19288 12084
rect 20399 12056 20444 12084
rect 18647 12053 18659 12056
rect 18601 12047 18659 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 22002 12044 22008 12096
rect 22060 12084 22066 12096
rect 27893 12087 27951 12093
rect 27893 12084 27905 12087
rect 22060 12056 27905 12084
rect 22060 12044 22066 12056
rect 27893 12053 27905 12056
rect 27939 12084 27951 12087
rect 28350 12084 28356 12096
rect 27939 12056 28356 12084
rect 27939 12053 27951 12056
rect 27893 12047 27951 12053
rect 28350 12044 28356 12056
rect 28408 12044 28414 12096
rect 31036 12084 31064 12124
rect 31386 12112 31392 12124
rect 31444 12112 31450 12164
rect 37918 12084 37924 12096
rect 31036 12056 37924 12084
rect 37918 12044 37924 12056
rect 37976 12044 37982 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 16724 11852 17693 11880
rect 16724 11840 16730 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 19058 11880 19064 11892
rect 19019 11852 19064 11880
rect 17681 11843 17739 11849
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 19208 11852 22140 11880
rect 19208 11840 19214 11852
rect 2961 11815 3019 11821
rect 2961 11781 2973 11815
rect 3007 11812 3019 11815
rect 3050 11812 3056 11824
rect 3007 11784 3056 11812
rect 3007 11781 3019 11784
rect 2961 11775 3019 11781
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3697 11815 3755 11821
rect 3697 11781 3709 11815
rect 3743 11812 3755 11815
rect 5074 11812 5080 11824
rect 3743 11784 5080 11812
rect 3743 11781 3755 11784
rect 3697 11775 3755 11781
rect 5074 11772 5080 11784
rect 5132 11772 5138 11824
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 22002 11812 22008 11824
rect 7892 11784 22008 11812
rect 7892 11772 7898 11784
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 22112 11812 22140 11852
rect 22186 11840 22192 11892
rect 22244 11880 22250 11892
rect 22373 11883 22431 11889
rect 22373 11880 22385 11883
rect 22244 11852 22385 11880
rect 22244 11840 22250 11852
rect 22373 11849 22385 11852
rect 22419 11849 22431 11883
rect 22373 11843 22431 11849
rect 27522 11840 27528 11892
rect 27580 11880 27586 11892
rect 30193 11883 30251 11889
rect 30193 11880 30205 11883
rect 27580 11852 30205 11880
rect 27580 11840 27586 11852
rect 30193 11849 30205 11852
rect 30239 11849 30251 11883
rect 30193 11843 30251 11849
rect 31113 11883 31171 11889
rect 31113 11849 31125 11883
rect 31159 11880 31171 11883
rect 31386 11880 31392 11892
rect 31159 11852 31392 11880
rect 31159 11849 31171 11852
rect 31113 11843 31171 11849
rect 31386 11840 31392 11852
rect 31444 11840 31450 11892
rect 24578 11812 24584 11824
rect 22112 11784 24584 11812
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 27617 11815 27675 11821
rect 27617 11781 27629 11815
rect 27663 11812 27675 11815
rect 27982 11812 27988 11824
rect 27663 11784 27988 11812
rect 27663 11781 27675 11784
rect 27617 11775 27675 11781
rect 27982 11772 27988 11784
rect 28040 11812 28046 11824
rect 28077 11815 28135 11821
rect 28077 11812 28089 11815
rect 28040 11784 28089 11812
rect 28040 11772 28046 11784
rect 28077 11781 28089 11784
rect 28123 11812 28135 11815
rect 30653 11815 30711 11821
rect 30653 11812 30665 11815
rect 28123 11784 30665 11812
rect 28123 11781 28135 11784
rect 28077 11775 28135 11781
rect 30653 11781 30665 11784
rect 30699 11812 30711 11815
rect 31573 11815 31631 11821
rect 31573 11812 31585 11815
rect 30699 11784 31585 11812
rect 30699 11781 30711 11784
rect 30653 11775 30711 11781
rect 31573 11781 31585 11784
rect 31619 11812 31631 11815
rect 32398 11812 32404 11824
rect 31619 11784 32404 11812
rect 31619 11781 31631 11784
rect 31573 11775 31631 11781
rect 32398 11772 32404 11784
rect 32456 11772 32462 11824
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2464 11716 2789 11744
rect 2464 11704 2470 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3384 11716 3525 11744
rect 3384 11704 3390 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11744 10195 11747
rect 20438 11744 20444 11756
rect 10183 11716 20444 11744
rect 10183 11713 10195 11716
rect 10137 11707 10195 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 22278 11744 22284 11756
rect 22239 11716 22284 11744
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 10928 11648 12081 11676
rect 10928 11636 10934 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 18141 11679 18199 11685
rect 12069 11639 12127 11645
rect 12176 11648 17908 11676
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 12176 11608 12204 11648
rect 9916 11580 12204 11608
rect 12437 11611 12495 11617
rect 9916 11568 9922 11580
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 12483 11580 13124 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 10318 11540 10324 11552
rect 10279 11512 10324 11540
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 12526 11540 12532 11552
rect 12487 11512 12532 11540
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13096 11549 13124 11580
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 17773 11611 17831 11617
rect 17773 11608 17785 11611
rect 15068 11580 17785 11608
rect 15068 11568 15074 11580
rect 17773 11577 17785 11580
rect 17819 11577 17831 11611
rect 17880 11608 17908 11648
rect 18141 11645 18153 11679
rect 18187 11676 18199 11679
rect 18601 11679 18659 11685
rect 18601 11676 18613 11679
rect 18187 11648 18613 11676
rect 18187 11645 18199 11648
rect 18141 11639 18199 11645
rect 18601 11645 18613 11648
rect 18647 11676 18659 11679
rect 19334 11676 19340 11688
rect 18647 11648 19340 11676
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 19334 11636 19340 11648
rect 19392 11676 19398 11688
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 19392 11648 19533 11676
rect 19392 11636 19398 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 18877 11611 18935 11617
rect 18877 11608 18889 11611
rect 17880 11580 18889 11608
rect 17773 11571 17831 11577
rect 18877 11577 18889 11580
rect 18923 11577 18935 11611
rect 18877 11571 18935 11577
rect 27062 11568 27068 11620
rect 27120 11608 27126 11620
rect 27249 11611 27307 11617
rect 27249 11608 27261 11611
rect 27120 11580 27261 11608
rect 27120 11568 27126 11580
rect 27249 11577 27261 11580
rect 27295 11577 27307 11611
rect 28350 11608 28356 11620
rect 28311 11580 28356 11608
rect 27249 11571 27307 11577
rect 28350 11568 28356 11580
rect 28408 11568 28414 11620
rect 30377 11611 30435 11617
rect 30377 11577 30389 11611
rect 30423 11577 30435 11611
rect 30377 11571 30435 11577
rect 13081 11543 13139 11549
rect 13081 11509 13093 11543
rect 13127 11540 13139 11543
rect 19150 11540 19156 11552
rect 13127 11512 19156 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 27157 11543 27215 11549
rect 27157 11509 27169 11543
rect 27203 11540 27215 11543
rect 28442 11540 28448 11552
rect 27203 11512 28448 11540
rect 27203 11509 27215 11512
rect 27157 11503 27215 11509
rect 28442 11500 28448 11512
rect 28500 11500 28506 11552
rect 28537 11543 28595 11549
rect 28537 11509 28549 11543
rect 28583 11540 28595 11543
rect 28994 11540 29000 11552
rect 28583 11512 29000 11540
rect 28583 11509 28595 11512
rect 28537 11503 28595 11509
rect 28994 11500 29000 11512
rect 29052 11500 29058 11552
rect 30392 11540 30420 11571
rect 30558 11568 30564 11620
rect 30616 11608 30622 11620
rect 31205 11611 31263 11617
rect 31205 11608 31217 11611
rect 30616 11580 31217 11608
rect 30616 11568 30622 11580
rect 31205 11577 31217 11580
rect 31251 11577 31263 11611
rect 31205 11571 31263 11577
rect 31938 11540 31944 11552
rect 30392 11512 31944 11540
rect 31938 11500 31944 11512
rect 31996 11500 32002 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 12713 11339 12771 11345
rect 12713 11305 12725 11339
rect 12759 11336 12771 11339
rect 15102 11336 15108 11348
rect 12759 11308 15108 11336
rect 12759 11305 12771 11308
rect 12713 11299 12771 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 27062 11336 27068 11348
rect 16356 11308 27068 11336
rect 16356 11296 16362 11308
rect 27062 11296 27068 11308
rect 27120 11296 27126 11348
rect 33226 11336 33232 11348
rect 33187 11308 33232 11336
rect 33226 11296 33232 11308
rect 33284 11296 33290 11348
rect 37918 11336 37924 11348
rect 37879 11308 37924 11336
rect 37918 11296 37924 11308
rect 37976 11296 37982 11348
rect 18325 11271 18383 11277
rect 18325 11237 18337 11271
rect 18371 11268 18383 11271
rect 19334 11268 19340 11280
rect 18371 11240 19340 11268
rect 18371 11237 18383 11240
rect 18325 11231 18383 11237
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 23106 11228 23112 11280
rect 23164 11268 23170 11280
rect 27798 11268 27804 11280
rect 23164 11240 27804 11268
rect 23164 11228 23170 11240
rect 27798 11228 27804 11240
rect 27856 11268 27862 11280
rect 28261 11271 28319 11277
rect 28261 11268 28273 11271
rect 27856 11240 28273 11268
rect 27856 11228 27862 11240
rect 28261 11237 28273 11240
rect 28307 11237 28319 11271
rect 28261 11231 28319 11237
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 2915 11172 14504 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2096 11104 2697 11132
rect 2096 11092 2102 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 10928 11104 12817 11132
rect 10928 11092 10934 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13630 11064 13636 11076
rect 13035 11036 13636 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 14476 11064 14504 11172
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 25590 11200 25596 11212
rect 16724 11172 25596 11200
rect 16724 11160 16730 11172
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 27982 11200 27988 11212
rect 27943 11172 27988 11200
rect 27982 11160 27988 11172
rect 28040 11160 28046 11212
rect 28445 11203 28503 11209
rect 28445 11169 28457 11203
rect 28491 11200 28503 11203
rect 30006 11200 30012 11212
rect 28491 11172 30012 11200
rect 28491 11169 28503 11172
rect 28445 11163 28503 11169
rect 30006 11160 30012 11172
rect 30064 11160 30070 11212
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 20346 11132 20352 11144
rect 14608 11104 20352 11132
rect 14608 11092 14614 11104
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 37369 11135 37427 11141
rect 37369 11101 37381 11135
rect 37415 11132 37427 11135
rect 38102 11132 38108 11144
rect 37415 11104 38108 11132
rect 37415 11101 37427 11104
rect 37369 11095 37427 11101
rect 38102 11092 38108 11104
rect 38160 11092 38166 11144
rect 16666 11064 16672 11076
rect 14476 11036 16672 11064
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 18156 11036 18368 11064
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 18156 10996 18184 11036
rect 3476 10968 18184 10996
rect 18340 10996 18368 11036
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 22097 11067 22155 11073
rect 22097 11064 22109 11067
rect 19392 11036 22109 11064
rect 19392 11024 19398 11036
rect 22097 11033 22109 11036
rect 22143 11064 22155 11067
rect 22278 11064 22284 11076
rect 22143 11036 22284 11064
rect 22143 11033 22155 11036
rect 22097 11027 22155 11033
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 30374 11024 30380 11076
rect 30432 11064 30438 11076
rect 33137 11067 33195 11073
rect 33137 11064 33149 11067
rect 30432 11036 33149 11064
rect 30432 11024 30438 11036
rect 33137 11033 33149 11036
rect 33183 11033 33195 11067
rect 33137 11027 33195 11033
rect 19426 10996 19432 11008
rect 18340 10968 19432 10996
rect 3476 10956 3482 10968
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 3234 10752 3240 10804
rect 3292 10792 3298 10804
rect 27798 10792 27804 10804
rect 3292 10764 6914 10792
rect 27759 10764 27804 10792
rect 3292 10752 3298 10764
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 5534 10724 5540 10736
rect 5123 10696 5540 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 6886 10724 6914 10764
rect 27798 10752 27804 10764
rect 27856 10752 27862 10804
rect 24394 10724 24400 10736
rect 6886 10696 24400 10724
rect 24394 10684 24400 10696
rect 24452 10684 24458 10736
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10656 4951 10659
rect 4982 10656 4988 10668
rect 4939 10628 4988 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12526 10656 12532 10668
rect 12207 10628 12532 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 35989 10659 36047 10665
rect 35989 10656 36001 10659
rect 19024 10628 36001 10656
rect 19024 10616 19030 10628
rect 35989 10625 36001 10628
rect 36035 10656 36047 10659
rect 36541 10659 36599 10665
rect 36541 10656 36553 10659
rect 36035 10628 36553 10656
rect 36035 10625 36047 10628
rect 35989 10619 36047 10625
rect 36541 10625 36553 10628
rect 36587 10625 36599 10659
rect 36541 10619 36599 10625
rect 37277 10659 37335 10665
rect 37277 10625 37289 10659
rect 37323 10625 37335 10659
rect 37277 10619 37335 10625
rect 3694 10548 3700 10600
rect 3752 10588 3758 10600
rect 25958 10588 25964 10600
rect 3752 10560 25964 10588
rect 3752 10548 3758 10560
rect 25958 10548 25964 10560
rect 26016 10548 26022 10600
rect 35894 10548 35900 10600
rect 35952 10588 35958 10600
rect 37292 10588 37320 10619
rect 35952 10560 37320 10588
rect 35952 10548 35958 10560
rect 21082 10480 21088 10532
rect 21140 10520 21146 10532
rect 37461 10523 37519 10529
rect 37461 10520 37473 10523
rect 21140 10492 37473 10520
rect 21140 10480 21146 10492
rect 37461 10489 37473 10492
rect 37507 10489 37519 10523
rect 37461 10483 37519 10489
rect 12345 10455 12403 10461
rect 12345 10421 12357 10455
rect 12391 10452 12403 10455
rect 12986 10452 12992 10464
rect 12391 10424 12992 10452
rect 12391 10421 12403 10424
rect 12345 10415 12403 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 36725 10455 36783 10461
rect 36725 10421 36737 10455
rect 36771 10452 36783 10455
rect 37274 10452 37280 10464
rect 36771 10424 37280 10452
rect 36771 10421 36783 10424
rect 36725 10415 36783 10421
rect 37274 10412 37280 10424
rect 37332 10412 37338 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2866 10248 2872 10260
rect 2827 10220 2872 10248
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 17681 10251 17739 10257
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 17862 10248 17868 10260
rect 17727 10220 17868 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 7098 10180 7104 10192
rect 6227 10152 7104 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 14829 10183 14887 10189
rect 14829 10149 14841 10183
rect 14875 10180 14887 10183
rect 17037 10183 17095 10189
rect 14875 10152 15516 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 15488 10053 15516 10152
rect 17037 10149 17049 10183
rect 17083 10180 17095 10183
rect 17402 10180 17408 10192
rect 17083 10152 17408 10180
rect 17083 10149 17095 10152
rect 17037 10143 17095 10149
rect 17402 10140 17408 10152
rect 17460 10140 17466 10192
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 35802 10112 35808 10124
rect 17175 10084 35808 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 35802 10072 35808 10084
rect 35860 10072 35866 10124
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10044 15531 10047
rect 25682 10044 25688 10056
rect 15519 10016 25688 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 25682 10004 25688 10016
rect 25740 10004 25746 10056
rect 28442 10044 28448 10056
rect 28403 10016 28448 10044
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 2774 9976 2780 9988
rect 2735 9948 2780 9976
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 5997 9979 6055 9985
rect 5997 9945 6009 9979
rect 6043 9976 6055 9979
rect 6178 9976 6184 9988
rect 6043 9948 6184 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 6178 9936 6184 9948
rect 6236 9936 6242 9988
rect 14274 9936 14280 9988
rect 14332 9976 14338 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 14332 9948 14473 9976
rect 14332 9936 14338 9948
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 14461 9939 14519 9945
rect 16669 9979 16727 9985
rect 16669 9945 16681 9979
rect 16715 9976 16727 9979
rect 17773 9979 17831 9985
rect 17773 9976 17785 9979
rect 16715 9948 16749 9976
rect 17512 9948 17785 9976
rect 16715 9945 16727 9948
rect 16669 9939 16727 9945
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 13504 9880 14933 9908
rect 13504 9868 13510 9880
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 14921 9871 14979 9877
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9908 16267 9911
rect 16684 9908 16712 9939
rect 17512 9920 17540 9948
rect 17773 9945 17785 9948
rect 17819 9945 17831 9979
rect 17773 9939 17831 9945
rect 17957 9979 18015 9985
rect 17957 9945 17969 9979
rect 18003 9945 18015 9979
rect 17957 9939 18015 9945
rect 17494 9908 17500 9920
rect 16255 9880 17500 9908
rect 16255 9877 16267 9880
rect 16209 9871 16267 9877
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 17972 9908 18000 9939
rect 18506 9908 18512 9920
rect 17972 9880 18512 9908
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 28629 9911 28687 9917
rect 28629 9877 28641 9911
rect 28675 9908 28687 9911
rect 29730 9908 29736 9920
rect 28675 9880 29736 9908
rect 28675 9877 28687 9880
rect 28629 9871 28687 9877
rect 29730 9868 29736 9880
rect 29788 9868 29794 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 17313 9707 17371 9713
rect 17313 9673 17325 9707
rect 17359 9704 17371 9707
rect 17402 9704 17408 9716
rect 17359 9676 17408 9704
rect 17359 9673 17371 9676
rect 17313 9667 17371 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 4614 9596 4620 9648
rect 4672 9636 4678 9648
rect 26878 9636 26884 9648
rect 4672 9608 26884 9636
rect 4672 9596 4678 9608
rect 26878 9596 26884 9608
rect 26936 9596 26942 9648
rect 13446 9568 13452 9580
rect 13407 9540 13452 9568
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 14274 9568 14280 9580
rect 13872 9540 14280 9568
rect 13872 9528 13878 9540
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 15930 9568 15936 9580
rect 14507 9540 15936 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 24765 9571 24823 9577
rect 24351 9540 24716 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9640 9472 9873 9500
rect 9640 9460 9646 9472
rect 9861 9469 9873 9472
rect 9907 9500 9919 9503
rect 22922 9500 22928 9512
rect 9907 9472 22928 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 24394 9500 24400 9512
rect 24355 9472 24400 9500
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 24688 9500 24716 9540
rect 24765 9537 24777 9571
rect 24811 9568 24823 9571
rect 25130 9568 25136 9580
rect 24811 9540 25136 9568
rect 24811 9537 24823 9540
rect 24765 9531 24823 9537
rect 25130 9528 25136 9540
rect 25188 9528 25194 9580
rect 28994 9568 29000 9580
rect 28955 9540 29000 9568
rect 28994 9528 29000 9540
rect 29052 9528 29058 9580
rect 30006 9568 30012 9580
rect 29967 9540 30012 9568
rect 30006 9528 30012 9540
rect 30064 9528 30070 9580
rect 37734 9568 37740 9580
rect 37695 9540 37740 9568
rect 37734 9528 37740 9540
rect 37792 9528 37798 9580
rect 25038 9500 25044 9512
rect 24688 9472 25044 9500
rect 25038 9460 25044 9472
rect 25096 9500 25102 9512
rect 25317 9503 25375 9509
rect 25317 9500 25329 9503
rect 25096 9472 25329 9500
rect 25096 9460 25102 9472
rect 25317 9469 25329 9472
rect 25363 9469 25375 9503
rect 38013 9503 38071 9509
rect 38013 9500 38025 9503
rect 25317 9463 25375 9469
rect 26206 9472 38025 9500
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 24670 9432 24676 9444
rect 3936 9404 24676 9432
rect 3936 9392 3942 9404
rect 24670 9392 24676 9404
rect 24728 9392 24734 9444
rect 25406 9392 25412 9444
rect 25464 9432 25470 9444
rect 26206 9432 26234 9472
rect 38013 9469 38025 9472
rect 38059 9469 38071 9503
rect 38013 9463 38071 9469
rect 25464 9404 26234 9432
rect 29181 9435 29239 9441
rect 25464 9392 25470 9404
rect 29181 9401 29193 9435
rect 29227 9432 29239 9435
rect 31018 9432 31024 9444
rect 29227 9404 31024 9432
rect 29227 9401 29239 9404
rect 29181 9395 29239 9401
rect 31018 9392 31024 9404
rect 31076 9392 31082 9444
rect 13633 9367 13691 9373
rect 13633 9333 13645 9367
rect 13679 9364 13691 9367
rect 13722 9364 13728 9376
rect 13679 9336 13728 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 15746 9364 15752 9376
rect 14231 9336 15752 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 30193 9367 30251 9373
rect 30193 9333 30205 9367
rect 30239 9364 30251 9367
rect 32214 9364 32220 9376
rect 30239 9336 32220 9364
rect 30239 9333 30251 9336
rect 30193 9327 30251 9333
rect 32214 9324 32220 9336
rect 32272 9324 32278 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3510 9160 3516 9172
rect 2884 9132 3516 9160
rect 2884 9101 2912 9132
rect 3510 9120 3516 9132
rect 3568 9160 3574 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 3568 9132 3801 9160
rect 3568 9120 3574 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 3789 9123 3847 9129
rect 4985 9163 5043 9169
rect 4985 9129 4997 9163
rect 5031 9160 5043 9163
rect 5258 9160 5264 9172
rect 5031 9132 5264 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 5258 9120 5264 9132
rect 5316 9160 5322 9172
rect 5316 9132 5764 9160
rect 5316 9120 5322 9132
rect 5736 9101 5764 9132
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 25777 9163 25835 9169
rect 25777 9160 25789 9163
rect 5868 9132 25789 9160
rect 5868 9120 5874 9132
rect 25777 9129 25789 9132
rect 25823 9129 25835 9163
rect 25777 9123 25835 9129
rect 34054 9120 34060 9172
rect 34112 9160 34118 9172
rect 34793 9163 34851 9169
rect 34793 9160 34805 9163
rect 34112 9132 34805 9160
rect 34112 9120 34118 9132
rect 34793 9129 34805 9132
rect 34839 9129 34851 9163
rect 34793 9123 34851 9129
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9061 2927 9095
rect 2869 9055 2927 9061
rect 5721 9095 5779 9101
rect 5721 9061 5733 9095
rect 5767 9061 5779 9095
rect 9582 9092 9588 9104
rect 9543 9064 9588 9092
rect 5721 9055 5779 9061
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 10505 9095 10563 9101
rect 10505 9061 10517 9095
rect 10551 9092 10563 9095
rect 11606 9092 11612 9104
rect 10551 9064 11612 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 20990 9092 20996 9104
rect 20951 9064 20996 9092
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 32306 9024 32312 9036
rect 12676 8996 32312 9024
rect 12676 8984 12682 8996
rect 32306 8984 32312 8996
rect 32364 8984 32370 9036
rect 35345 9027 35403 9033
rect 35345 8993 35357 9027
rect 35391 9024 35403 9027
rect 36078 9024 36084 9036
rect 35391 8996 36084 9024
rect 35391 8993 35403 8996
rect 35345 8987 35403 8993
rect 36078 8984 36084 8996
rect 36136 8984 36142 9036
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 9232 8928 10333 8956
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 3050 8888 3056 8900
rect 2547 8860 3056 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 5408 8860 5457 8888
rect 5408 8848 5414 8860
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 5445 8851 5503 8857
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9232 8897 9260 8928
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8956 20223 8959
rect 20346 8956 20352 8968
rect 20211 8928 20352 8956
rect 20211 8925 20223 8928
rect 20165 8919 20223 8925
rect 20346 8916 20352 8928
rect 20404 8956 20410 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20404 8928 20637 8956
rect 20404 8916 20410 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 24489 8959 24547 8965
rect 24489 8956 24501 8959
rect 23900 8928 24501 8956
rect 23900 8916 23906 8928
rect 24489 8925 24501 8928
rect 24535 8925 24547 8959
rect 24489 8919 24547 8925
rect 24949 8959 25007 8965
rect 24949 8925 24961 8959
rect 24995 8956 25007 8959
rect 25038 8956 25044 8968
rect 24995 8928 25044 8956
rect 24995 8925 25007 8928
rect 24949 8919 25007 8925
rect 25038 8916 25044 8928
rect 25096 8956 25102 8968
rect 25869 8959 25927 8965
rect 25869 8956 25881 8959
rect 25096 8928 25881 8956
rect 25096 8916 25102 8928
rect 25869 8925 25881 8928
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 9088 8860 9229 8888
rect 9088 8848 9094 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 9217 8851 9275 8857
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 9548 8860 10149 8888
rect 9548 8848 9554 8860
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 21637 8891 21695 8897
rect 21637 8888 21649 8891
rect 21048 8860 21649 8888
rect 21048 8848 21054 8860
rect 21637 8857 21649 8860
rect 21683 8888 21695 8891
rect 25222 8888 25228 8900
rect 21683 8860 25228 8888
rect 21683 8857 21695 8860
rect 21637 8851 21695 8857
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 2958 8820 2964 8832
rect 2919 8792 2964 8820
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 5902 8820 5908 8832
rect 5863 8792 5908 8820
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9766 8820 9772 8832
rect 9723 8792 9772 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 21085 8823 21143 8829
rect 21085 8820 21097 8823
rect 20220 8792 21097 8820
rect 20220 8780 20226 8792
rect 21085 8789 21097 8792
rect 21131 8789 21143 8823
rect 21085 8783 21143 8789
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 23382 8820 23388 8832
rect 21232 8792 23388 8820
rect 21232 8780 21238 8792
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 24670 8820 24676 8832
rect 24631 8792 24676 8820
rect 24670 8780 24676 8792
rect 24728 8780 24734 8832
rect 25884 8820 25912 8919
rect 35802 8916 35808 8968
rect 35860 8956 35866 8968
rect 35897 8959 35955 8965
rect 35897 8956 35909 8959
rect 35860 8928 35909 8956
rect 35860 8916 35866 8928
rect 35897 8925 35909 8928
rect 35943 8956 35955 8959
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 35943 8928 36553 8956
rect 35943 8925 35955 8928
rect 35897 8919 35955 8925
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 36541 8919 36599 8925
rect 37461 8959 37519 8965
rect 37461 8925 37473 8959
rect 37507 8956 37519 8959
rect 38102 8956 38108 8968
rect 37507 8928 38108 8956
rect 37507 8925 37519 8928
rect 37461 8919 37519 8925
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 26053 8891 26111 8897
rect 26053 8857 26065 8891
rect 26099 8888 26111 8891
rect 26970 8888 26976 8900
rect 26099 8860 26976 8888
rect 26099 8857 26111 8860
rect 26053 8851 26111 8857
rect 26970 8848 26976 8860
rect 27028 8848 27034 8900
rect 34790 8848 34796 8900
rect 34848 8888 34854 8900
rect 35069 8891 35127 8897
rect 35069 8888 35081 8891
rect 34848 8860 35081 8888
rect 34848 8848 34854 8860
rect 35069 8857 35081 8860
rect 35115 8857 35127 8891
rect 35069 8851 35127 8857
rect 36004 8860 37964 8888
rect 26326 8820 26332 8832
rect 25884 8792 26332 8820
rect 26326 8780 26332 8792
rect 26384 8820 26390 8832
rect 26513 8823 26571 8829
rect 26513 8820 26525 8823
rect 26384 8792 26525 8820
rect 26384 8780 26390 8792
rect 26513 8789 26525 8792
rect 26559 8789 26571 8823
rect 26513 8783 26571 8789
rect 35253 8823 35311 8829
rect 35253 8789 35265 8823
rect 35299 8820 35311 8823
rect 36004 8820 36032 8860
rect 35299 8792 36032 8820
rect 36081 8823 36139 8829
rect 35299 8789 35311 8792
rect 35253 8783 35311 8789
rect 36081 8789 36093 8823
rect 36127 8820 36139 8823
rect 36446 8820 36452 8832
rect 36127 8792 36452 8820
rect 36127 8789 36139 8792
rect 36081 8783 36139 8789
rect 36446 8780 36452 8792
rect 36504 8780 36510 8832
rect 37936 8829 37964 8860
rect 37921 8823 37979 8829
rect 37921 8789 37933 8823
rect 37967 8789 37979 8823
rect 37921 8783 37979 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8616 2743 8619
rect 2774 8616 2780 8628
rect 2731 8588 2780 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4614 8616 4620 8628
rect 4203 8588 4620 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 21174 8616 21180 8628
rect 5960 8588 12572 8616
rect 5960 8576 5966 8588
rect 2958 8508 2964 8560
rect 3016 8548 3022 8560
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 3016 8520 4077 8548
rect 3016 8508 3022 8520
rect 4065 8517 4077 8520
rect 4111 8517 4123 8551
rect 4065 8511 4123 8517
rect 6365 8551 6423 8557
rect 6365 8517 6377 8551
rect 6411 8548 6423 8551
rect 6454 8548 6460 8560
rect 6411 8520 6460 8548
rect 6411 8517 6423 8520
rect 6365 8511 6423 8517
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 7285 8551 7343 8557
rect 7285 8548 7297 8551
rect 6886 8520 7297 8548
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3418 8480 3424 8492
rect 3099 8452 3424 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 2884 8412 2912 8443
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5408 8452 6561 8480
rect 5408 8440 5414 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6886 8480 6914 8520
rect 7285 8517 7297 8520
rect 7331 8548 7343 8551
rect 9950 8548 9956 8560
rect 7331 8520 9956 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 12544 8548 12572 8588
rect 19306 8588 21180 8616
rect 16482 8548 16488 8560
rect 12544 8520 16488 8548
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 9766 8480 9772 8492
rect 6779 8452 6914 8480
rect 9727 8452 9772 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 19306 8480 19334 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 23937 8619 23995 8625
rect 23937 8585 23949 8619
rect 23983 8616 23995 8619
rect 24854 8616 24860 8628
rect 23983 8588 24860 8616
rect 23983 8585 23995 8588
rect 23937 8579 23995 8585
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 34606 8616 34612 8628
rect 25280 8588 34612 8616
rect 25280 8576 25286 8588
rect 34606 8576 34612 8588
rect 34664 8576 34670 8628
rect 37826 8576 37832 8628
rect 37884 8616 37890 8628
rect 38105 8619 38163 8625
rect 38105 8616 38117 8619
rect 37884 8588 38117 8616
rect 37884 8576 37890 8588
rect 38105 8585 38117 8588
rect 38151 8616 38163 8619
rect 38562 8616 38568 8628
rect 38151 8588 38568 8616
rect 38151 8585 38163 8588
rect 38105 8579 38163 8585
rect 38562 8576 38568 8588
rect 38620 8576 38626 8628
rect 20346 8508 20352 8560
rect 20404 8548 20410 8560
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 20404 8520 20729 8548
rect 20404 8508 20410 8520
rect 20717 8517 20729 8520
rect 20763 8517 20775 8551
rect 20717 8511 20775 8517
rect 20901 8551 20959 8557
rect 20901 8517 20913 8551
rect 20947 8548 20959 8551
rect 30374 8548 30380 8560
rect 20947 8520 30380 8548
rect 20947 8517 20959 8520
rect 20901 8511 20959 8517
rect 30374 8508 30380 8520
rect 30432 8508 30438 8560
rect 32306 8548 32312 8560
rect 32267 8520 32312 8548
rect 32306 8508 32312 8520
rect 32364 8508 32370 8560
rect 32766 8508 32772 8560
rect 32824 8548 32830 8560
rect 33229 8551 33287 8557
rect 33229 8548 33241 8551
rect 32824 8520 33241 8548
rect 32824 8508 32830 8520
rect 33229 8517 33241 8520
rect 33275 8517 33287 8551
rect 33229 8511 33287 8517
rect 33413 8551 33471 8557
rect 33413 8517 33425 8551
rect 33459 8548 33471 8551
rect 36078 8548 36084 8560
rect 33459 8520 36084 8548
rect 33459 8517 33471 8520
rect 33413 8511 33471 8517
rect 12575 8452 19334 8480
rect 19889 8483 19947 8489
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20162 8480 20168 8492
rect 19935 8452 20168 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 11517 8415 11575 8421
rect 2884 8384 3096 8412
rect 3068 8356 3096 8384
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 11606 8412 11612 8424
rect 11563 8384 11612 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 3050 8304 3056 8356
rect 3108 8304 3114 8356
rect 9953 8347 10011 8353
rect 9953 8313 9965 8347
rect 9999 8344 10011 8347
rect 11790 8344 11796 8356
rect 9999 8316 11796 8344
rect 9999 8313 10011 8316
rect 9953 8307 10011 8313
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 11885 8347 11943 8353
rect 11885 8313 11897 8347
rect 11931 8344 11943 8347
rect 12544 8344 12572 8443
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 11931 8316 12572 8344
rect 20073 8347 20131 8353
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 20073 8313 20085 8347
rect 20119 8344 20131 8347
rect 20254 8344 20260 8356
rect 20119 8316 20260 8344
rect 20119 8313 20131 8316
rect 20073 8307 20131 8313
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 20548 8344 20576 8443
rect 25222 8440 25228 8492
rect 25280 8480 25286 8492
rect 25590 8480 25596 8492
rect 25280 8452 25596 8480
rect 25280 8440 25286 8452
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 32674 8480 32680 8492
rect 32635 8452 32680 8480
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8381 24455 8415
rect 24397 8375 24455 8381
rect 32217 8415 32275 8421
rect 32217 8381 32229 8415
rect 32263 8412 32275 8415
rect 32306 8412 32312 8424
rect 32263 8384 32312 8412
rect 32263 8381 32275 8384
rect 32217 8375 32275 8381
rect 20714 8344 20720 8356
rect 20548 8316 20720 8344
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 23474 8344 23480 8356
rect 23435 8316 23480 8344
rect 23474 8304 23480 8316
rect 23532 8344 23538 8356
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23532 8316 24041 8344
rect 23532 8304 23538 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 24412 8344 24440 8375
rect 32306 8372 32312 8384
rect 32364 8412 32370 8424
rect 33428 8412 33456 8511
rect 36078 8508 36084 8520
rect 36136 8508 36142 8560
rect 33594 8480 33600 8492
rect 33555 8452 33600 8480
rect 33594 8440 33600 8452
rect 33652 8440 33658 8492
rect 32364 8384 33456 8412
rect 35713 8415 35771 8421
rect 32364 8372 32370 8384
rect 35713 8381 35725 8415
rect 35759 8412 35771 8415
rect 37918 8412 37924 8424
rect 35759 8384 37924 8412
rect 35759 8381 35771 8384
rect 35713 8375 35771 8381
rect 37918 8372 37924 8384
rect 37976 8372 37982 8424
rect 24949 8347 25007 8353
rect 24949 8344 24961 8347
rect 24412 8316 24961 8344
rect 24029 8307 24087 8313
rect 24949 8313 24961 8316
rect 24995 8344 25007 8347
rect 25501 8347 25559 8353
rect 25501 8344 25513 8347
rect 24995 8316 25513 8344
rect 24995 8313 25007 8316
rect 24949 8307 25007 8313
rect 25501 8313 25513 8316
rect 25547 8344 25559 8347
rect 26326 8344 26332 8356
rect 25547 8316 26332 8344
rect 25547 8313 25559 8316
rect 25501 8307 25559 8313
rect 26326 8304 26332 8316
rect 26384 8304 26390 8356
rect 36262 8344 36268 8356
rect 36223 8316 36268 8344
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 37458 8344 37464 8356
rect 37419 8316 37464 8344
rect 37458 8304 37464 8316
rect 37516 8304 37522 8356
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 11977 8279 12035 8285
rect 11977 8276 11989 8279
rect 11572 8248 11989 8276
rect 11572 8236 11578 8248
rect 11977 8245 11989 8248
rect 12023 8245 12035 8279
rect 11977 8239 12035 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 36906 8032 36912 8084
rect 36964 8072 36970 8084
rect 37185 8075 37243 8081
rect 37185 8072 37197 8075
rect 36964 8044 37197 8072
rect 36964 8032 36970 8044
rect 37185 8041 37197 8044
rect 37231 8041 37243 8075
rect 37185 8035 37243 8041
rect 11793 8007 11851 8013
rect 11793 7973 11805 8007
rect 11839 8004 11851 8007
rect 13354 8004 13360 8016
rect 11839 7976 13360 8004
rect 11839 7973 11851 7976
rect 11793 7967 11851 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 30193 8007 30251 8013
rect 30193 7973 30205 8007
rect 30239 8004 30251 8007
rect 32950 8004 32956 8016
rect 30239 7976 32956 8004
rect 30239 7973 30251 7976
rect 30193 7967 30251 7973
rect 32950 7964 32956 7976
rect 33008 7964 33014 8016
rect 31846 7896 31852 7948
rect 31904 7936 31910 7948
rect 32033 7939 32091 7945
rect 32033 7936 32045 7939
rect 31904 7908 32045 7936
rect 31904 7896 31910 7908
rect 32033 7905 32045 7908
rect 32079 7905 32091 7939
rect 32033 7899 32091 7905
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 11606 7868 11612 7880
rect 9732 7840 11612 7868
rect 9732 7828 9738 7840
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 24854 7868 24860 7880
rect 24815 7840 24860 7868
rect 24854 7828 24860 7840
rect 24912 7828 24918 7880
rect 32398 7868 32404 7880
rect 32359 7840 32404 7868
rect 32398 7828 32404 7840
rect 32456 7828 32462 7880
rect 38102 7868 38108 7880
rect 38063 7840 38108 7868
rect 38102 7828 38108 7840
rect 38160 7828 38166 7880
rect 11422 7800 11428 7812
rect 11383 7772 11428 7800
rect 11422 7760 11428 7772
rect 11480 7760 11486 7812
rect 30006 7800 30012 7812
rect 29967 7772 30012 7800
rect 30006 7760 30012 7772
rect 30064 7760 30070 7812
rect 31941 7803 31999 7809
rect 31941 7769 31953 7803
rect 31987 7800 31999 7803
rect 32306 7800 32312 7812
rect 31987 7772 32312 7800
rect 31987 7769 31999 7772
rect 31941 7763 31999 7769
rect 32306 7760 32312 7772
rect 32364 7760 32370 7812
rect 35069 7803 35127 7809
rect 35069 7769 35081 7803
rect 35115 7800 35127 7803
rect 35710 7800 35716 7812
rect 35115 7772 35716 7800
rect 35115 7769 35127 7772
rect 35069 7763 35127 7769
rect 35710 7760 35716 7772
rect 35768 7760 35774 7812
rect 36722 7760 36728 7812
rect 36780 7800 36786 7812
rect 37093 7803 37151 7809
rect 37093 7800 37105 7803
rect 36780 7772 37105 7800
rect 36780 7760 36786 7772
rect 37093 7769 37105 7772
rect 37139 7769 37151 7803
rect 37093 7763 37151 7769
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3418 7732 3424 7744
rect 3283 7704 3424 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 20346 7732 20352 7744
rect 20307 7704 20352 7732
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 25041 7735 25099 7741
rect 25041 7701 25053 7735
rect 25087 7732 25099 7735
rect 25866 7732 25872 7744
rect 25087 7704 25872 7732
rect 25087 7701 25099 7704
rect 25041 7695 25099 7701
rect 25866 7692 25872 7704
rect 25924 7692 25930 7744
rect 35342 7692 35348 7744
rect 35400 7732 35406 7744
rect 35529 7735 35587 7741
rect 35529 7732 35541 7735
rect 35400 7704 35541 7732
rect 35400 7692 35406 7704
rect 35529 7701 35541 7704
rect 35575 7701 35587 7735
rect 35529 7695 35587 7701
rect 36541 7735 36599 7741
rect 36541 7701 36553 7735
rect 36587 7732 36599 7735
rect 38194 7732 38200 7744
rect 36587 7704 38200 7732
rect 36587 7701 36599 7704
rect 36541 7695 36599 7701
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 25038 7528 25044 7540
rect 7055 7500 25044 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 28626 7528 28632 7540
rect 28092 7500 28632 7528
rect 7469 7463 7527 7469
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 8110 7460 8116 7472
rect 7515 7432 8116 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 14182 7420 14188 7472
rect 14240 7460 14246 7472
rect 28092 7469 28120 7500
rect 28626 7488 28632 7500
rect 28684 7488 28690 7540
rect 15197 7463 15255 7469
rect 15197 7460 15209 7463
rect 14240 7432 15209 7460
rect 14240 7420 14246 7432
rect 15197 7429 15209 7432
rect 15243 7429 15255 7463
rect 28077 7463 28135 7469
rect 15197 7423 15255 7429
rect 18432 7432 28028 7460
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 6886 7364 7665 7392
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 6730 7324 6736 7336
rect 6595 7296 6736 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 6730 7284 6736 7296
rect 6788 7324 6794 7336
rect 6886 7324 6914 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 11514 7392 11520 7404
rect 7883 7364 8432 7392
rect 11475 7364 11520 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 6788 7296 6914 7324
rect 6788 7284 6794 7296
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 8404 7265 8432 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 15381 7395 15439 7401
rect 15381 7392 15393 7395
rect 14292 7364 15393 7392
rect 14292 7336 14320 7364
rect 15381 7361 15393 7364
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16206 7392 16212 7404
rect 15611 7364 16212 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 14274 7324 14280 7336
rect 14235 7296 14280 7324
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 17218 7324 17224 7336
rect 14568 7296 17224 7324
rect 6825 7259 6883 7265
rect 6825 7256 6837 7259
rect 6696 7228 6837 7256
rect 6696 7216 6702 7228
rect 6825 7225 6837 7228
rect 6871 7225 6883 7259
rect 6825 7219 6883 7225
rect 8389 7259 8447 7265
rect 8389 7225 8401 7259
rect 8435 7256 8447 7259
rect 14568 7256 14596 7296
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 8435 7228 14596 7256
rect 14645 7259 14703 7265
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 14645 7225 14657 7259
rect 14691 7256 14703 7259
rect 14918 7256 14924 7268
rect 14691 7228 14924 7256
rect 14691 7225 14703 7228
rect 14645 7219 14703 7225
rect 14918 7216 14924 7228
rect 14976 7216 14982 7268
rect 18432 7256 18460 7432
rect 26421 7395 26479 7401
rect 26421 7392 26433 7395
rect 15212 7228 18460 7256
rect 18524 7364 26433 7392
rect 11701 7191 11759 7197
rect 11701 7157 11713 7191
rect 11747 7188 11759 7191
rect 12618 7188 12624 7200
rect 11747 7160 12624 7188
rect 11747 7157 11759 7160
rect 11701 7151 11759 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15212 7188 15240 7228
rect 14783 7160 15240 7188
rect 16117 7191 16175 7197
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 16117 7157 16129 7191
rect 16163 7188 16175 7191
rect 16206 7188 16212 7200
rect 16163 7160 16212 7188
rect 16163 7157 16175 7160
rect 16117 7151 16175 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 18524 7188 18552 7364
rect 26421 7361 26433 7364
rect 26467 7392 26479 7395
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26467 7364 26985 7392
rect 26467 7361 26479 7364
rect 26421 7355 26479 7361
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 28000 7392 28028 7432
rect 28077 7429 28089 7463
rect 28123 7429 28135 7463
rect 37826 7460 37832 7472
rect 37787 7432 37832 7460
rect 28077 7423 28135 7429
rect 37826 7420 37832 7432
rect 37884 7420 37890 7472
rect 33962 7392 33968 7404
rect 28000 7364 33968 7392
rect 26973 7355 27031 7361
rect 33962 7352 33968 7364
rect 34020 7352 34026 7404
rect 35986 7352 35992 7404
rect 36044 7392 36050 7404
rect 36538 7392 36544 7404
rect 36044 7364 36544 7392
rect 36044 7352 36050 7364
rect 36538 7352 36544 7364
rect 36596 7352 36602 7404
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7324 20407 7327
rect 20438 7324 20444 7336
rect 20395 7296 20444 7324
rect 20395 7293 20407 7296
rect 20349 7287 20407 7293
rect 20438 7284 20444 7296
rect 20496 7284 20502 7336
rect 34057 7327 34115 7333
rect 34057 7293 34069 7327
rect 34103 7324 34115 7327
rect 37826 7324 37832 7336
rect 34103 7296 37832 7324
rect 34103 7293 34115 7296
rect 34057 7287 34115 7293
rect 37826 7284 37832 7296
rect 37884 7284 37890 7336
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 20588 7228 20637 7256
rect 20588 7216 20594 7228
rect 20625 7225 20637 7228
rect 20671 7225 20683 7259
rect 20625 7219 20683 7225
rect 27614 7216 27620 7268
rect 27672 7256 27678 7268
rect 27893 7259 27951 7265
rect 27893 7256 27905 7259
rect 27672 7228 27905 7256
rect 27672 7216 27678 7228
rect 27893 7225 27905 7228
rect 27939 7225 27951 7259
rect 27893 7219 27951 7225
rect 30926 7216 30932 7268
rect 30984 7256 30990 7268
rect 37645 7259 37703 7265
rect 37645 7256 37657 7259
rect 30984 7228 37657 7256
rect 30984 7216 30990 7228
rect 37645 7225 37657 7228
rect 37691 7225 37703 7259
rect 37645 7219 37703 7225
rect 20806 7188 20812 7200
rect 16540 7160 18552 7188
rect 20767 7160 20812 7188
rect 16540 7148 16546 7160
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 27157 7191 27215 7197
rect 27157 7157 27169 7191
rect 27203 7188 27215 7191
rect 27798 7188 27804 7200
rect 27203 7160 27804 7188
rect 27203 7157 27215 7160
rect 27157 7151 27215 7157
rect 27798 7148 27804 7160
rect 27856 7148 27862 7200
rect 34606 7188 34612 7200
rect 34567 7160 34612 7188
rect 34606 7148 34612 7160
rect 34664 7148 34670 7200
rect 35621 7191 35679 7197
rect 35621 7157 35633 7191
rect 35667 7188 35679 7191
rect 35986 7188 35992 7200
rect 35667 7160 35992 7188
rect 35667 7157 35679 7160
rect 35621 7151 35679 7157
rect 35986 7148 35992 7160
rect 36044 7148 36050 7200
rect 36170 7188 36176 7200
rect 36131 7160 36176 7188
rect 36170 7148 36176 7160
rect 36228 7148 36234 7200
rect 36725 7191 36783 7197
rect 36725 7157 36737 7191
rect 36771 7188 36783 7191
rect 38102 7188 38108 7200
rect 36771 7160 38108 7188
rect 36771 7157 36783 7160
rect 36725 7151 36783 7157
rect 38102 7148 38108 7160
rect 38160 7148 38166 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 14918 6984 14924 6996
rect 14879 6956 14924 6984
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 28902 6984 28908 6996
rect 17276 6956 28908 6984
rect 17276 6944 17282 6956
rect 28902 6944 28908 6956
rect 28960 6944 28966 6996
rect 16853 6919 16911 6925
rect 16853 6885 16865 6919
rect 16899 6885 16911 6919
rect 16853 6879 16911 6885
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6696 6820 7113 6848
rect 6696 6808 6702 6820
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 16022 6848 16028 6860
rect 15983 6820 16028 6848
rect 7101 6811 7159 6817
rect 16022 6808 16028 6820
rect 16080 6848 16086 6860
rect 16868 6848 16896 6879
rect 20530 6876 20536 6928
rect 20588 6916 20594 6928
rect 20901 6919 20959 6925
rect 20901 6916 20913 6919
rect 20588 6888 20913 6916
rect 20588 6876 20594 6888
rect 20901 6885 20913 6888
rect 20947 6885 20959 6919
rect 20901 6879 20959 6885
rect 23198 6876 23204 6928
rect 23256 6916 23262 6928
rect 30926 6916 30932 6928
rect 23256 6888 30932 6916
rect 23256 6876 23262 6888
rect 30926 6876 30932 6888
rect 30984 6876 30990 6928
rect 31757 6919 31815 6925
rect 31757 6885 31769 6919
rect 31803 6885 31815 6919
rect 31757 6879 31815 6885
rect 16080 6820 16896 6848
rect 17037 6851 17095 6857
rect 16080 6808 16086 6820
rect 17037 6817 17049 6851
rect 17083 6848 17095 6851
rect 17083 6820 22094 6848
rect 17083 6817 17095 6820
rect 17037 6811 17095 6817
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 20806 6780 20812 6792
rect 19567 6752 20812 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 22066 6780 22094 6820
rect 24946 6808 24952 6860
rect 25004 6848 25010 6860
rect 25041 6851 25099 6857
rect 25041 6848 25053 6851
rect 25004 6820 25053 6848
rect 25004 6808 25010 6820
rect 25041 6817 25053 6820
rect 25087 6817 25099 6851
rect 25041 6811 25099 6817
rect 25148 6820 28672 6848
rect 25148 6780 25176 6820
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 22066 6752 25176 6780
rect 25240 6752 27629 6780
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 16577 6715 16635 6721
rect 16577 6712 16589 6715
rect 16540 6684 16589 6712
rect 16540 6672 16546 6684
rect 16577 6681 16589 6684
rect 16623 6681 16635 6715
rect 19978 6712 19984 6724
rect 19939 6684 19984 6712
rect 16577 6675 16635 6681
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 20165 6715 20223 6721
rect 20165 6681 20177 6715
rect 20211 6681 20223 6715
rect 20165 6675 20223 6681
rect 20349 6715 20407 6721
rect 20349 6681 20361 6715
rect 20395 6712 20407 6715
rect 24854 6712 24860 6724
rect 20395 6684 22094 6712
rect 24815 6684 24860 6712
rect 20395 6681 20407 6684
rect 20349 6675 20407 6681
rect 5258 6644 5264 6656
rect 5219 6616 5264 6644
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 19426 6644 19432 6656
rect 19383 6616 19432 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 20180 6644 20208 6675
rect 20438 6644 20444 6656
rect 20180 6616 20444 6644
rect 20438 6604 20444 6616
rect 20496 6644 20502 6656
rect 20622 6644 20628 6656
rect 20496 6616 20628 6644
rect 20496 6604 20502 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 22066 6644 22094 6684
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 25038 6672 25044 6724
rect 25096 6712 25102 6724
rect 25240 6712 25268 6752
rect 27617 6749 27629 6752
rect 27663 6780 27675 6783
rect 28261 6783 28319 6789
rect 28261 6780 28273 6783
rect 27663 6752 28273 6780
rect 27663 6749 27675 6752
rect 27617 6743 27675 6749
rect 28261 6749 28273 6752
rect 28307 6749 28319 6783
rect 28644 6780 28672 6820
rect 28718 6808 28724 6860
rect 28776 6848 28782 6860
rect 31113 6851 31171 6857
rect 31113 6848 31125 6851
rect 28776 6820 31125 6848
rect 28776 6808 28782 6820
rect 31113 6817 31125 6820
rect 31159 6848 31171 6851
rect 31772 6848 31800 6879
rect 31159 6820 31800 6848
rect 32125 6851 32183 6857
rect 31159 6817 31171 6820
rect 31113 6811 31171 6817
rect 32125 6817 32137 6851
rect 32171 6848 32183 6851
rect 32306 6848 32312 6860
rect 32171 6820 32312 6848
rect 32171 6817 32183 6820
rect 32125 6811 32183 6817
rect 32306 6808 32312 6820
rect 32364 6808 32370 6860
rect 35253 6783 35311 6789
rect 35253 6780 35265 6783
rect 28644 6752 35265 6780
rect 28261 6743 28319 6749
rect 35253 6749 35265 6752
rect 35299 6780 35311 6783
rect 35618 6780 35624 6792
rect 35299 6752 35624 6780
rect 35299 6749 35311 6752
rect 35253 6743 35311 6749
rect 35618 6740 35624 6752
rect 35676 6740 35682 6792
rect 37185 6783 37243 6789
rect 37185 6749 37197 6783
rect 37231 6749 37243 6783
rect 37185 6743 37243 6749
rect 30006 6712 30012 6724
rect 25096 6684 25268 6712
rect 26206 6684 30012 6712
rect 25096 6672 25102 6684
rect 26206 6644 26234 6684
rect 30006 6672 30012 6684
rect 30064 6672 30070 6724
rect 33229 6715 33287 6721
rect 33229 6681 33241 6715
rect 33275 6712 33287 6715
rect 34514 6712 34520 6724
rect 33275 6684 34520 6712
rect 33275 6681 33287 6684
rect 33229 6675 33287 6681
rect 34514 6672 34520 6684
rect 34572 6672 34578 6724
rect 34793 6715 34851 6721
rect 34793 6681 34805 6715
rect 34839 6712 34851 6715
rect 35342 6712 35348 6724
rect 34839 6684 35348 6712
rect 34839 6681 34851 6684
rect 34793 6675 34851 6681
rect 35342 6672 35348 6684
rect 35400 6672 35406 6724
rect 36725 6715 36783 6721
rect 36725 6681 36737 6715
rect 36771 6712 36783 6715
rect 37200 6712 37228 6743
rect 37274 6740 37280 6792
rect 37332 6780 37338 6792
rect 37829 6783 37887 6789
rect 37829 6780 37841 6783
rect 37332 6752 37841 6780
rect 37332 6740 37338 6752
rect 37829 6749 37841 6752
rect 37875 6749 37887 6783
rect 37829 6743 37887 6749
rect 39574 6712 39580 6724
rect 36771 6684 39580 6712
rect 36771 6681 36783 6684
rect 36725 6675 36783 6681
rect 39574 6672 39580 6684
rect 39632 6672 39638 6724
rect 22066 6616 26234 6644
rect 27801 6647 27859 6653
rect 27801 6613 27813 6647
rect 27847 6644 27859 6647
rect 28626 6644 28632 6656
rect 27847 6616 28632 6644
rect 27847 6613 27859 6616
rect 27801 6607 27859 6613
rect 28626 6604 28632 6616
rect 28684 6604 28690 6656
rect 29914 6644 29920 6656
rect 29875 6616 29920 6644
rect 29914 6604 29920 6616
rect 29972 6604 29978 6656
rect 30374 6604 30380 6656
rect 30432 6644 30438 6656
rect 30561 6647 30619 6653
rect 30561 6644 30573 6647
rect 30432 6616 30573 6644
rect 30432 6604 30438 6616
rect 30561 6613 30573 6616
rect 30607 6613 30619 6647
rect 30561 6607 30619 6613
rect 31665 6647 31723 6653
rect 31665 6613 31677 6647
rect 31711 6644 31723 6647
rect 32306 6644 32312 6656
rect 31711 6616 32312 6644
rect 31711 6613 31723 6616
rect 31665 6607 31723 6613
rect 32306 6604 32312 6616
rect 32364 6604 32370 6656
rect 32582 6644 32588 6656
rect 32543 6616 32588 6644
rect 32582 6604 32588 6616
rect 32640 6604 32646 6656
rect 33781 6647 33839 6653
rect 33781 6613 33793 6647
rect 33827 6644 33839 6647
rect 33870 6644 33876 6656
rect 33827 6616 33876 6644
rect 33827 6613 33839 6616
rect 33781 6607 33839 6613
rect 33870 6604 33876 6616
rect 33928 6604 33934 6656
rect 35802 6604 35808 6656
rect 35860 6644 35866 6656
rect 36081 6647 36139 6653
rect 36081 6644 36093 6647
rect 35860 6616 36093 6644
rect 35860 6604 35866 6616
rect 36081 6613 36093 6616
rect 36127 6613 36139 6647
rect 37366 6644 37372 6656
rect 37327 6616 37372 6644
rect 36081 6607 36139 6613
rect 37366 6604 37372 6616
rect 37424 6604 37430 6656
rect 38013 6647 38071 6653
rect 38013 6613 38025 6647
rect 38059 6644 38071 6647
rect 38470 6644 38476 6656
rect 38059 6616 38476 6644
rect 38059 6613 38071 6616
rect 38013 6607 38071 6613
rect 38470 6604 38476 6616
rect 38528 6604 38534 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 5166 6440 5172 6452
rect 4387 6412 5172 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4356 6304 4384 6403
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 15562 6440 15568 6452
rect 15523 6412 15568 6440
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 35437 6443 35495 6449
rect 35437 6409 35449 6443
rect 35483 6440 35495 6443
rect 35894 6440 35900 6452
rect 35483 6412 35900 6440
rect 35483 6409 35495 6412
rect 35437 6403 35495 6409
rect 35894 6400 35900 6412
rect 35952 6400 35958 6452
rect 36725 6443 36783 6449
rect 36725 6409 36737 6443
rect 36771 6440 36783 6443
rect 37734 6440 37740 6452
rect 36771 6412 37740 6440
rect 36771 6409 36783 6412
rect 36725 6403 36783 6409
rect 37734 6400 37740 6412
rect 37792 6400 37798 6452
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 16669 6375 16727 6381
rect 16669 6372 16681 6375
rect 16632 6344 16681 6372
rect 16632 6332 16638 6344
rect 16669 6341 16681 6344
rect 16715 6341 16727 6375
rect 16669 6335 16727 6341
rect 34793 6375 34851 6381
rect 34793 6341 34805 6375
rect 34839 6372 34851 6375
rect 34839 6344 35940 6372
rect 34839 6341 34851 6344
rect 34793 6335 34851 6341
rect 35912 6316 35940 6344
rect 35986 6332 35992 6384
rect 36044 6372 36050 6384
rect 36044 6344 36584 6372
rect 36044 6332 36050 6344
rect 3712 6276 4384 6304
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 2832 6208 3341 6236
rect 2832 6196 2838 6208
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 3329 6199 3387 6205
rect 3712 6177 3740 6276
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 16482 6304 16488 6316
rect 15896 6276 16488 6304
rect 15896 6264 15902 6276
rect 16482 6264 16488 6276
rect 16540 6304 16546 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16540 6276 16865 6304
rect 16540 6264 16546 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17678 6304 17684 6316
rect 17083 6276 17684 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 35250 6304 35256 6316
rect 35211 6276 35256 6304
rect 35250 6264 35256 6276
rect 35308 6264 35314 6316
rect 35894 6264 35900 6316
rect 35952 6304 35958 6316
rect 36556 6313 36584 6344
rect 37366 6332 37372 6384
rect 37424 6372 37430 6384
rect 37829 6375 37887 6381
rect 37829 6372 37841 6375
rect 37424 6344 37841 6372
rect 37424 6332 37430 6344
rect 37829 6341 37841 6344
rect 37875 6372 37887 6375
rect 38746 6372 38752 6384
rect 37875 6344 38752 6372
rect 37875 6341 37887 6344
rect 37829 6335 37887 6341
rect 38746 6332 38752 6344
rect 38804 6332 38810 6384
rect 36081 6307 36139 6313
rect 36081 6304 36093 6307
rect 35952 6276 36093 6304
rect 35952 6264 35958 6276
rect 36081 6273 36093 6276
rect 36127 6273 36139 6307
rect 36081 6267 36139 6273
rect 36541 6307 36599 6313
rect 36541 6273 36553 6307
rect 36587 6304 36599 6307
rect 39022 6304 39028 6316
rect 36587 6276 39028 6304
rect 36587 6273 36599 6276
rect 36541 6267 36599 6273
rect 39022 6264 39028 6276
rect 39080 6264 39086 6316
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6236 3847 6239
rect 25682 6236 25688 6248
rect 3835 6208 25688 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 31846 6196 31852 6248
rect 31904 6236 31910 6248
rect 31904 6208 35940 6236
rect 31904 6196 31910 6208
rect 3697 6171 3755 6177
rect 3697 6137 3709 6171
rect 3743 6137 3755 6171
rect 3697 6131 3755 6137
rect 30006 6128 30012 6180
rect 30064 6168 30070 6180
rect 31481 6171 31539 6177
rect 31481 6168 31493 6171
rect 30064 6140 31493 6168
rect 30064 6128 30070 6140
rect 31481 6137 31493 6140
rect 31527 6137 31539 6171
rect 31481 6131 31539 6137
rect 33689 6171 33747 6177
rect 33689 6137 33701 6171
rect 33735 6168 33747 6171
rect 34514 6168 34520 6180
rect 33735 6140 34520 6168
rect 33735 6137 33747 6140
rect 33689 6131 33747 6137
rect 34514 6128 34520 6140
rect 34572 6128 34578 6180
rect 35912 6177 35940 6208
rect 35897 6171 35955 6177
rect 35897 6137 35909 6171
rect 35943 6137 35955 6171
rect 35897 6131 35955 6137
rect 1489 6103 1547 6109
rect 1489 6069 1501 6103
rect 1535 6100 1547 6103
rect 1578 6100 1584 6112
rect 1535 6072 1584 6100
rect 1535 6069 1547 6072
rect 1489 6063 1547 6069
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2498 6100 2504 6112
rect 2459 6072 2504 6100
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5442 6100 5448 6112
rect 5403 6072 5448 6100
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 15102 6100 15108 6112
rect 15063 6072 15108 6100
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 17589 6103 17647 6109
rect 17589 6069 17601 6103
rect 17635 6100 17647 6103
rect 17678 6100 17684 6112
rect 17635 6072 17684 6100
rect 17635 6069 17647 6072
rect 17589 6063 17647 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 29638 6100 29644 6112
rect 29599 6072 29644 6100
rect 29638 6060 29644 6072
rect 29696 6060 29702 6112
rect 30466 6100 30472 6112
rect 30427 6072 30472 6100
rect 30466 6060 30472 6072
rect 30524 6060 30530 6112
rect 30926 6100 30932 6112
rect 30887 6072 30932 6100
rect 30926 6060 30932 6072
rect 30984 6060 30990 6112
rect 31754 6060 31760 6112
rect 31812 6100 31818 6112
rect 32125 6103 32183 6109
rect 32125 6100 32137 6103
rect 31812 6072 32137 6100
rect 31812 6060 31818 6072
rect 32125 6069 32137 6072
rect 32171 6069 32183 6103
rect 32950 6100 32956 6112
rect 32911 6072 32956 6100
rect 32125 6063 32183 6069
rect 32950 6060 32956 6072
rect 33008 6060 33014 6112
rect 34054 6060 34060 6112
rect 34112 6100 34118 6112
rect 34149 6103 34207 6109
rect 34149 6100 34161 6103
rect 34112 6072 34161 6100
rect 34112 6060 34118 6072
rect 34149 6069 34161 6072
rect 34195 6069 34207 6103
rect 37734 6100 37740 6112
rect 37695 6072 37740 6100
rect 34149 6063 34207 6069
rect 37734 6060 37740 6072
rect 37792 6060 37798 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 4706 5896 4712 5908
rect 3835 5868 4712 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 16114 5896 16120 5908
rect 16075 5868 16120 5896
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 18472 5868 18521 5896
rect 18472 5856 18478 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 30650 5896 30656 5908
rect 30611 5868 30656 5896
rect 18509 5859 18567 5865
rect 30650 5856 30656 5868
rect 30708 5856 30714 5908
rect 31202 5896 31208 5908
rect 31163 5868 31208 5896
rect 31202 5856 31208 5868
rect 31260 5856 31266 5908
rect 32674 5856 32680 5908
rect 32732 5896 32738 5908
rect 33321 5899 33379 5905
rect 33321 5896 33333 5899
rect 32732 5868 33333 5896
rect 32732 5856 32738 5868
rect 33321 5865 33333 5868
rect 33367 5865 33379 5899
rect 33962 5896 33968 5908
rect 33923 5868 33968 5896
rect 33321 5859 33379 5865
rect 33962 5856 33968 5868
rect 34020 5856 34026 5908
rect 34790 5856 34796 5908
rect 34848 5896 34854 5908
rect 34885 5899 34943 5905
rect 34885 5896 34897 5899
rect 34848 5868 34897 5896
rect 34848 5856 34854 5868
rect 34885 5865 34897 5868
rect 34931 5865 34943 5899
rect 34885 5859 34943 5865
rect 36449 5899 36507 5905
rect 36449 5865 36461 5899
rect 36495 5896 36507 5899
rect 39298 5896 39304 5908
rect 36495 5868 39304 5896
rect 36495 5865 36507 5868
rect 36449 5859 36507 5865
rect 39298 5856 39304 5868
rect 39356 5856 39362 5908
rect 24026 5788 24032 5840
rect 24084 5828 24090 5840
rect 37734 5828 37740 5840
rect 24084 5800 37740 5828
rect 24084 5788 24090 5800
rect 37734 5788 37740 5800
rect 37792 5788 37798 5840
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 13814 5760 13820 5772
rect 12575 5732 13820 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 29917 5763 29975 5769
rect 29917 5760 29929 5763
rect 22336 5732 29929 5760
rect 22336 5720 22342 5732
rect 29917 5729 29929 5732
rect 29963 5729 29975 5763
rect 29917 5723 29975 5729
rect 36078 5720 36084 5772
rect 36136 5760 36142 5772
rect 37829 5763 37887 5769
rect 37829 5760 37841 5763
rect 36136 5732 37841 5760
rect 36136 5720 36142 5732
rect 37829 5729 37841 5732
rect 37875 5729 37887 5763
rect 37829 5723 37887 5729
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 6696 5664 12633 5692
rect 6696 5652 6702 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 25682 5692 25688 5704
rect 25643 5664 25688 5692
rect 12621 5655 12679 5661
rect 25682 5652 25688 5664
rect 25740 5692 25746 5704
rect 26329 5695 26387 5701
rect 26329 5692 26341 5695
rect 25740 5664 26341 5692
rect 25740 5652 25746 5664
rect 26329 5661 26341 5664
rect 26375 5661 26387 5695
rect 26329 5655 26387 5661
rect 30101 5695 30159 5701
rect 30101 5661 30113 5695
rect 30147 5692 30159 5695
rect 30650 5692 30656 5704
rect 30147 5664 30656 5692
rect 30147 5661 30159 5664
rect 30101 5655 30159 5661
rect 30650 5652 30656 5664
rect 30708 5652 30714 5704
rect 33505 5695 33563 5701
rect 33505 5692 33517 5695
rect 33244 5664 33517 5692
rect 1762 5584 1768 5636
rect 1820 5624 1826 5636
rect 2501 5627 2559 5633
rect 2501 5624 2513 5627
rect 1820 5596 2513 5624
rect 1820 5584 1826 5596
rect 2501 5593 2513 5596
rect 2547 5593 2559 5627
rect 2501 5587 2559 5593
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3973 5627 4031 5633
rect 3973 5624 3985 5627
rect 2832 5596 3985 5624
rect 2832 5584 2838 5596
rect 3973 5593 3985 5596
rect 4019 5593 4031 5627
rect 3973 5587 4031 5593
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4706 5624 4712 5636
rect 4203 5596 4712 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 24854 5624 24860 5636
rect 13096 5596 24860 5624
rect 1394 5556 1400 5568
rect 1355 5528 1400 5556
rect 1394 5516 1400 5528
rect 1452 5516 1458 5568
rect 1670 5516 1676 5568
rect 1728 5556 1734 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1728 5528 1961 5556
rect 1728 5516 1734 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 3142 5556 3148 5568
rect 3103 5528 3148 5556
rect 1949 5519 2007 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 5132 5528 5181 5556
rect 5132 5516 5138 5528
rect 5169 5525 5181 5528
rect 5215 5525 5227 5559
rect 5169 5519 5227 5525
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5684 5528 5733 5556
rect 5684 5516 5690 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 6362 5556 6368 5568
rect 6323 5528 6368 5556
rect 5721 5519 5779 5525
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 8018 5556 8024 5568
rect 6972 5528 7017 5556
rect 7979 5528 8024 5556
rect 6972 5516 6978 5528
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11146 5556 11152 5568
rect 11103 5528 11152 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13096 5565 13124 5596
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 33244 5568 33272 5664
rect 33505 5661 33517 5664
rect 33551 5661 33563 5695
rect 33505 5655 33563 5661
rect 34054 5652 34060 5704
rect 34112 5692 34118 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 34112 5664 34713 5692
rect 34112 5652 34118 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 35437 5695 35495 5701
rect 35437 5661 35449 5695
rect 35483 5692 35495 5695
rect 35618 5692 35624 5704
rect 35483 5664 35624 5692
rect 35483 5661 35495 5664
rect 35437 5655 35495 5661
rect 35618 5652 35624 5664
rect 35676 5652 35682 5704
rect 36630 5692 36636 5704
rect 36591 5664 36636 5692
rect 36630 5652 36636 5664
rect 36688 5652 36694 5704
rect 37090 5692 37096 5704
rect 37051 5664 37096 5692
rect 37090 5652 37096 5664
rect 37148 5652 37154 5704
rect 35802 5584 35808 5636
rect 35860 5624 35866 5636
rect 38010 5624 38016 5636
rect 35860 5596 38016 5624
rect 35860 5584 35866 5596
rect 38010 5584 38016 5596
rect 38068 5584 38074 5636
rect 13081 5559 13139 5565
rect 13081 5525 13093 5559
rect 13127 5525 13139 5559
rect 14182 5556 14188 5568
rect 14143 5528 14188 5556
rect 13081 5519 13139 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15654 5556 15660 5568
rect 15615 5528 15660 5556
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 20349 5559 20407 5565
rect 20349 5556 20361 5559
rect 20128 5528 20361 5556
rect 20128 5516 20134 5528
rect 20349 5525 20361 5528
rect 20395 5525 20407 5559
rect 20349 5519 20407 5525
rect 20898 5516 20904 5568
rect 20956 5556 20962 5568
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 20956 5528 21189 5556
rect 20956 5516 20962 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 22094 5556 22100 5568
rect 22055 5528 22100 5556
rect 21177 5519 21235 5525
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 24486 5556 24492 5568
rect 24447 5528 24492 5556
rect 24486 5516 24492 5528
rect 24544 5516 24550 5568
rect 25222 5556 25228 5568
rect 25135 5528 25228 5556
rect 25222 5516 25228 5528
rect 25280 5556 25286 5568
rect 25406 5556 25412 5568
rect 25280 5528 25412 5556
rect 25280 5516 25286 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 25869 5559 25927 5565
rect 25869 5525 25881 5559
rect 25915 5556 25927 5559
rect 26418 5556 26424 5568
rect 25915 5528 26424 5556
rect 25915 5525 25927 5528
rect 25869 5519 25927 5525
rect 26418 5516 26424 5528
rect 26476 5516 26482 5568
rect 26510 5516 26516 5568
rect 26568 5556 26574 5568
rect 26878 5556 26884 5568
rect 26568 5528 26884 5556
rect 26568 5516 26574 5528
rect 26878 5516 26884 5528
rect 26936 5516 26942 5568
rect 28997 5559 29055 5565
rect 28997 5525 29009 5559
rect 29043 5556 29055 5559
rect 29086 5556 29092 5568
rect 29043 5528 29092 5556
rect 29043 5525 29055 5528
rect 28997 5519 29055 5525
rect 29086 5516 29092 5528
rect 29144 5516 29150 5568
rect 31294 5516 31300 5568
rect 31352 5556 31358 5568
rect 31941 5559 31999 5565
rect 31941 5556 31953 5559
rect 31352 5528 31953 5556
rect 31352 5516 31358 5528
rect 31941 5525 31953 5528
rect 31987 5525 31999 5559
rect 31941 5519 31999 5525
rect 32861 5559 32919 5565
rect 32861 5525 32873 5559
rect 32907 5556 32919 5559
rect 33226 5556 33232 5568
rect 32907 5528 33232 5556
rect 32907 5525 32919 5528
rect 32861 5519 32919 5525
rect 33226 5516 33232 5528
rect 33284 5516 33290 5568
rect 35621 5559 35679 5565
rect 35621 5525 35633 5559
rect 35667 5556 35679 5559
rect 36078 5556 36084 5568
rect 35667 5528 36084 5556
rect 35667 5525 35679 5528
rect 35621 5519 35679 5525
rect 36078 5516 36084 5528
rect 36136 5516 36142 5568
rect 37277 5559 37335 5565
rect 37277 5525 37289 5559
rect 37323 5556 37335 5559
rect 37734 5556 37740 5568
rect 37323 5528 37740 5556
rect 37323 5525 37335 5528
rect 37277 5519 37335 5525
rect 37734 5516 37740 5528
rect 37792 5516 37798 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 26050 5312 26056 5364
rect 26108 5352 26114 5364
rect 26329 5355 26387 5361
rect 26329 5352 26341 5355
rect 26108 5324 26341 5352
rect 26108 5312 26114 5324
rect 26329 5321 26341 5324
rect 26375 5352 26387 5355
rect 26602 5352 26608 5364
rect 26375 5324 26608 5352
rect 26375 5321 26387 5324
rect 26329 5315 26387 5321
rect 26602 5312 26608 5324
rect 26660 5312 26666 5364
rect 29270 5352 29276 5364
rect 29231 5324 29276 5352
rect 29270 5312 29276 5324
rect 29328 5312 29334 5364
rect 31938 5312 31944 5364
rect 31996 5352 32002 5364
rect 32125 5355 32183 5361
rect 32125 5352 32137 5355
rect 31996 5324 32137 5352
rect 31996 5312 32002 5324
rect 32125 5321 32137 5324
rect 32171 5321 32183 5355
rect 32125 5315 32183 5321
rect 32398 5312 32404 5364
rect 32456 5352 32462 5364
rect 33045 5355 33103 5361
rect 33045 5352 33057 5355
rect 32456 5324 33057 5352
rect 32456 5312 32462 5324
rect 33045 5321 33057 5324
rect 33091 5321 33103 5355
rect 33045 5315 33103 5321
rect 33594 5312 33600 5364
rect 33652 5352 33658 5364
rect 33873 5355 33931 5361
rect 33873 5352 33885 5355
rect 33652 5324 33885 5352
rect 33652 5312 33658 5324
rect 33873 5321 33885 5324
rect 33919 5321 33931 5355
rect 34882 5352 34888 5364
rect 34843 5324 34888 5352
rect 33873 5315 33931 5321
rect 34882 5312 34888 5324
rect 34940 5312 34946 5364
rect 35526 5352 35532 5364
rect 35487 5324 35532 5352
rect 35526 5312 35532 5324
rect 35584 5312 35590 5364
rect 37366 5352 37372 5364
rect 37327 5324 37372 5352
rect 37366 5312 37372 5324
rect 37424 5312 37430 5364
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 13262 5284 13268 5296
rect 12308 5256 13268 5284
rect 12308 5244 12314 5256
rect 13262 5244 13268 5256
rect 13320 5244 13326 5296
rect 29288 5216 29316 5312
rect 31294 5244 31300 5296
rect 31352 5284 31358 5296
rect 31352 5256 31754 5284
rect 31352 5244 31358 5256
rect 29825 5219 29883 5225
rect 29825 5216 29837 5219
rect 29288 5188 29837 5216
rect 29825 5185 29837 5188
rect 29871 5185 29883 5219
rect 29825 5179 29883 5185
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5216 30619 5219
rect 30650 5216 30656 5228
rect 30607 5188 30656 5216
rect 30607 5185 30619 5188
rect 30561 5179 30619 5185
rect 30650 5176 30656 5188
rect 30708 5176 30714 5228
rect 31202 5176 31208 5228
rect 31260 5216 31266 5228
rect 31389 5219 31447 5225
rect 31389 5216 31401 5219
rect 31260 5188 31401 5216
rect 31260 5176 31266 5188
rect 31389 5185 31401 5188
rect 31435 5185 31447 5219
rect 31726 5216 31754 5256
rect 32858 5244 32864 5296
rect 32916 5284 32922 5296
rect 35621 5287 35679 5293
rect 35621 5284 35633 5287
rect 32916 5256 35633 5284
rect 32916 5244 32922 5256
rect 35621 5253 35633 5256
rect 35667 5253 35679 5287
rect 35621 5247 35679 5253
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31726 5188 32321 5216
rect 31389 5179 31447 5185
rect 32309 5185 32321 5188
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 32950 5176 32956 5228
rect 33008 5216 33014 5228
rect 33229 5219 33287 5225
rect 33229 5216 33241 5219
rect 33008 5188 33241 5216
rect 33008 5176 33014 5188
rect 33229 5185 33241 5188
rect 33275 5185 33287 5219
rect 33229 5179 33287 5185
rect 33870 5176 33876 5228
rect 33928 5216 33934 5228
rect 34057 5219 34115 5225
rect 34057 5216 34069 5219
rect 33928 5188 34069 5216
rect 33928 5176 33934 5188
rect 34057 5185 34069 5188
rect 34103 5185 34115 5219
rect 34057 5179 34115 5185
rect 34238 5176 34244 5228
rect 34296 5216 34302 5228
rect 34793 5219 34851 5225
rect 34793 5216 34805 5219
rect 34296 5188 34805 5216
rect 34296 5176 34302 5188
rect 34793 5185 34805 5188
rect 34839 5185 34851 5219
rect 36446 5216 36452 5228
rect 36407 5188 36452 5216
rect 34793 5179 34851 5185
rect 36446 5176 36452 5188
rect 36504 5176 36510 5228
rect 38102 5216 38108 5228
rect 38063 5188 38108 5216
rect 38102 5176 38108 5188
rect 38160 5176 38166 5228
rect 11698 5108 11704 5160
rect 11756 5148 11762 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 11756 5120 12265 5148
rect 11756 5108 11762 5120
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 27430 5108 27436 5160
rect 27488 5148 27494 5160
rect 27488 5120 32996 5148
rect 27488 5108 27494 5120
rect 4525 5083 4583 5089
rect 4525 5049 4537 5083
rect 4571 5080 4583 5083
rect 4706 5080 4712 5092
rect 4571 5052 4712 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 16390 5040 16396 5092
rect 16448 5080 16454 5092
rect 27614 5080 27620 5092
rect 16448 5052 27620 5080
rect 16448 5040 16454 5052
rect 27614 5040 27620 5052
rect 27672 5040 27678 5092
rect 30009 5083 30067 5089
rect 30009 5049 30021 5083
rect 30055 5080 30067 5083
rect 32030 5080 32036 5092
rect 30055 5052 32036 5080
rect 30055 5049 30067 5052
rect 30009 5043 30067 5049
rect 32030 5040 32036 5052
rect 32088 5040 32094 5092
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 2590 5012 2596 5024
rect 2551 4984 2596 5012
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 3016 4984 3065 5012
rect 3016 4972 3022 4984
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 3694 5012 3700 5024
rect 3655 4984 3700 5012
rect 3053 4975 3111 4981
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4672 4984 4997 5012
rect 4672 4972 4678 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 4985 4975 5043 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6454 5012 6460 5024
rect 6415 4984 6460 5012
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 7190 5012 7196 5024
rect 7151 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 7929 5015 7987 5021
rect 7929 5012 7941 5015
rect 7800 4984 7941 5012
rect 7800 4972 7806 4984
rect 7929 4981 7941 4984
rect 7975 4981 7987 5015
rect 7929 4975 7987 4981
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 8260 4984 8493 5012
rect 8260 4972 8266 4984
rect 8481 4981 8493 4984
rect 8527 4981 8539 5015
rect 8481 4975 8539 4981
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 8628 4984 9045 5012
rect 8628 4972 8634 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 9582 5012 9588 5024
rect 9543 4984 9588 5012
rect 9033 4975 9091 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 10134 5012 10140 5024
rect 10095 4984 10140 5012
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11296 4984 11713 5012
rect 11296 4972 11302 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12584 4984 12817 5012
rect 12584 4972 12590 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 13354 5012 13360 5024
rect 13315 4984 13360 5012
rect 12805 4975 12863 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14090 5012 14096 5024
rect 14047 4984 14096 5012
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14826 5012 14832 5024
rect 14787 4984 14832 5012
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 15746 5012 15752 5024
rect 15707 4984 15752 5012
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 16482 4972 16488 5024
rect 16540 5012 16546 5024
rect 16669 5015 16727 5021
rect 16669 5012 16681 5015
rect 16540 4984 16681 5012
rect 16540 4972 16546 4984
rect 16669 4981 16681 4984
rect 16715 4981 16727 5015
rect 17218 5012 17224 5024
rect 17179 4984 17224 5012
rect 16669 4975 16727 4981
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 18322 5012 18328 5024
rect 18283 4984 18328 5012
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 18966 5012 18972 5024
rect 18927 4984 18972 5012
rect 18966 4972 18972 4984
rect 19024 4972 19030 5024
rect 19150 4972 19156 5024
rect 19208 5012 19214 5024
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 19208 4984 19441 5012
rect 19208 4972 19214 4984
rect 19429 4981 19441 4984
rect 19475 4981 19487 5015
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 19429 4975 19487 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 21085 5015 21143 5021
rect 21085 4981 21097 5015
rect 21131 5012 21143 5015
rect 21174 5012 21180 5024
rect 21131 4984 21180 5012
rect 21131 4981 21143 4984
rect 21085 4975 21143 4981
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 21450 4972 21456 5024
rect 21508 5012 21514 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21508 4984 21833 5012
rect 21508 4972 21514 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 22370 5012 22376 5024
rect 22331 4984 22376 5012
rect 21821 4975 21879 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 22925 5015 22983 5021
rect 22925 5012 22937 5015
rect 22612 4984 22937 5012
rect 22612 4972 22618 4984
rect 22925 4981 22937 4984
rect 22971 4981 22983 5015
rect 22925 4975 22983 4981
rect 23753 5015 23811 5021
rect 23753 4981 23765 5015
rect 23799 5012 23811 5015
rect 24210 5012 24216 5024
rect 23799 4984 24216 5012
rect 23799 4981 23811 4984
rect 23753 4975 23811 4981
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 24305 5015 24363 5021
rect 24305 4981 24317 5015
rect 24351 5012 24363 5015
rect 24394 5012 24400 5024
rect 24351 4984 24400 5012
rect 24351 4981 24363 4984
rect 24305 4975 24363 4981
rect 24394 4972 24400 4984
rect 24452 4972 24458 5024
rect 25038 5012 25044 5024
rect 24999 4984 25044 5012
rect 25038 4972 25044 4984
rect 25096 4972 25102 5024
rect 25777 5015 25835 5021
rect 25777 4981 25789 5015
rect 25823 5012 25835 5015
rect 26694 5012 26700 5024
rect 25823 4984 26700 5012
rect 25823 4981 25835 4984
rect 25777 4975 25835 4981
rect 26694 4972 26700 4984
rect 26752 4972 26758 5024
rect 27522 5012 27528 5024
rect 27483 4984 27528 5012
rect 27522 4972 27528 4984
rect 27580 4972 27586 5024
rect 27982 5012 27988 5024
rect 27943 4984 27988 5012
rect 27982 4972 27988 4984
rect 28040 4972 28046 5024
rect 28074 4972 28080 5024
rect 28132 5012 28138 5024
rect 28629 5015 28687 5021
rect 28629 5012 28641 5015
rect 28132 4984 28641 5012
rect 28132 4972 28138 4984
rect 28629 4981 28641 4984
rect 28675 4981 28687 5015
rect 28629 4975 28687 4981
rect 31573 5015 31631 5021
rect 31573 4981 31585 5015
rect 31619 5012 31631 5015
rect 31938 5012 31944 5024
rect 31619 4984 31944 5012
rect 31619 4981 31631 4984
rect 31573 4975 31631 4981
rect 31938 4972 31944 4984
rect 31996 4972 32002 5024
rect 32968 5012 32996 5120
rect 37921 5083 37979 5089
rect 37921 5080 37933 5083
rect 34900 5052 37933 5080
rect 34900 5012 34928 5052
rect 37921 5049 37933 5052
rect 37967 5049 37979 5083
rect 37921 5043 37979 5049
rect 32968 4984 34928 5012
rect 36633 5015 36691 5021
rect 36633 4981 36645 5015
rect 36679 5012 36691 5015
rect 36814 5012 36820 5024
rect 36679 4984 36820 5012
rect 36679 4981 36691 4984
rect 36633 4975 36691 4981
rect 36814 4972 36820 4984
rect 36872 4972 36878 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 5166 4808 5172 4820
rect 2271 4780 5172 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 9585 4811 9643 4817
rect 9585 4777 9597 4811
rect 9631 4808 9643 4811
rect 9631 4780 12434 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 2866 4740 2872 4752
rect 1627 4712 2872 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 5537 4743 5595 4749
rect 5537 4709 5549 4743
rect 5583 4740 5595 4743
rect 8478 4740 8484 4752
rect 5583 4712 8484 4740
rect 5583 4709 5595 4712
rect 5537 4703 5595 4709
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 12250 4740 12256 4752
rect 12211 4712 12256 4740
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 12406 4740 12434 4780
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 12768 4780 14105 4808
rect 12768 4768 12774 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 25130 4808 25136 4820
rect 25091 4780 25136 4808
rect 14093 4771 14151 4777
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 30558 4808 30564 4820
rect 26620 4780 30420 4808
rect 30519 4780 30564 4808
rect 19334 4740 19340 4752
rect 12406 4712 19340 4740
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 21085 4743 21143 4749
rect 21085 4709 21097 4743
rect 21131 4740 21143 4743
rect 22186 4740 22192 4752
rect 21131 4712 22192 4740
rect 21131 4709 21143 4712
rect 21085 4703 21143 4709
rect 22186 4700 22192 4712
rect 22244 4700 22250 4752
rect 8294 4672 8300 4684
rect 2884 4644 8300 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1578 4604 1584 4616
rect 1443 4576 1584 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 1820 4576 2053 4604
rect 1820 4564 1826 4576
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2685 4607 2743 4613
rect 2685 4604 2697 4607
rect 2556 4576 2697 4604
rect 2556 4564 2562 4576
rect 2685 4573 2697 4576
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2884 4477 2912 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 22462 4672 22468 4684
rect 8435 4644 12572 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 5316 4576 5365 4604
rect 5316 4564 5322 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6972 4576 7113 4604
rect 6972 4564 6978 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 7984 4576 9168 4604
rect 7984 4564 7990 4576
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8205 4539 8263 4545
rect 8205 4536 8217 4539
rect 7800 4508 8217 4536
rect 7800 4496 7806 4508
rect 8205 4505 8217 4508
rect 8251 4505 8263 4539
rect 9030 4536 9036 4548
rect 8991 4508 9036 4536
rect 8205 4499 8263 4505
rect 9030 4496 9036 4508
rect 9088 4496 9094 4548
rect 9140 4545 9168 4576
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11204 4576 11345 4604
rect 11204 4564 11210 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 9125 4539 9183 4545
rect 9125 4505 9137 4539
rect 9171 4505 9183 4539
rect 9125 4499 9183 4505
rect 9309 4539 9367 4545
rect 9309 4505 9321 4539
rect 9355 4536 9367 4539
rect 12544 4536 12572 4644
rect 16592 4644 22468 4672
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 12768 4576 13001 4604
rect 12768 4564 12774 4576
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 13354 4604 13360 4616
rect 13035 4576 13360 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13446 4564 13452 4616
rect 13504 4604 13510 4616
rect 14182 4604 14188 4616
rect 13504 4576 14188 4604
rect 13504 4564 13510 4576
rect 14182 4564 14188 4576
rect 14240 4604 14246 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 14240 4576 14289 4604
rect 14240 4564 14246 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 16390 4604 16396 4616
rect 15795 4576 16396 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16592 4613 16620 4644
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 25958 4672 25964 4684
rect 25919 4644 25964 4672
rect 25958 4632 25964 4644
rect 26016 4632 26022 4684
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 20070 4604 20076 4616
rect 16577 4567 16635 4573
rect 17052 4576 19932 4604
rect 20031 4576 20076 4604
rect 17052 4536 17080 4576
rect 9355 4508 11192 4536
rect 12544 4508 17080 4536
rect 17129 4539 17187 4545
rect 9355 4505 9367 4508
rect 9309 4499 9367 4505
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4437 2927 4471
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 2869 4431 2927 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 4212 4440 4353 4468
rect 4212 4428 4218 4440
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 6086 4468 6092 4480
rect 6047 4440 6092 4468
rect 4341 4431 4399 4437
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6546 4468 6552 4480
rect 6507 4440 6552 4468
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 8110 4468 8116 4480
rect 7331 4440 8116 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 11164 4477 11192 4508
rect 17129 4505 17141 4539
rect 17175 4536 17187 4539
rect 17494 4536 17500 4548
rect 17175 4508 17500 4536
rect 17175 4505 17187 4508
rect 17129 4499 17187 4505
rect 17494 4496 17500 4508
rect 17552 4496 17558 4548
rect 19904 4536 19932 4576
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 21508 4576 21557 4604
rect 21508 4564 21514 4576
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 21726 4564 21732 4616
rect 21784 4604 21790 4616
rect 22094 4604 22100 4616
rect 21784 4576 22100 4604
rect 21784 4564 21790 4576
rect 22094 4564 22100 4576
rect 22152 4604 22158 4616
rect 22189 4607 22247 4613
rect 22189 4604 22201 4607
rect 22152 4576 22201 4604
rect 22152 4564 22158 4576
rect 22189 4573 22201 4576
rect 22235 4573 22247 4607
rect 22189 4567 22247 4573
rect 25038 4564 25044 4616
rect 25096 4604 25102 4616
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 25096 4576 25329 4604
rect 25096 4564 25102 4576
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 26620 4613 26648 4780
rect 27246 4700 27252 4752
rect 27304 4740 27310 4752
rect 27985 4743 28043 4749
rect 27985 4740 27997 4743
rect 27304 4712 27997 4740
rect 27304 4700 27310 4712
rect 27985 4709 27997 4712
rect 28031 4709 28043 4743
rect 30392 4740 30420 4780
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 33413 4811 33471 4817
rect 33413 4777 33425 4811
rect 33459 4808 33471 4811
rect 33502 4808 33508 4820
rect 33459 4780 33508 4808
rect 33459 4777 33471 4780
rect 33413 4771 33471 4777
rect 33502 4768 33508 4780
rect 33560 4768 33566 4820
rect 31846 4740 31852 4752
rect 30392 4712 31852 4740
rect 27985 4703 28043 4709
rect 31846 4700 31852 4712
rect 31904 4700 31910 4752
rect 32309 4743 32367 4749
rect 32309 4709 32321 4743
rect 32355 4740 32367 4743
rect 33594 4740 33600 4752
rect 32355 4712 33600 4740
rect 32355 4709 32367 4712
rect 32309 4703 32367 4709
rect 33594 4700 33600 4712
rect 33652 4700 33658 4752
rect 35345 4743 35403 4749
rect 35345 4709 35357 4743
rect 35391 4740 35403 4743
rect 35434 4740 35440 4752
rect 35391 4712 35440 4740
rect 35391 4709 35403 4712
rect 35345 4703 35403 4709
rect 35434 4700 35440 4712
rect 35492 4700 35498 4752
rect 27062 4632 27068 4684
rect 27120 4672 27126 4684
rect 27120 4644 33272 4672
rect 27120 4632 27126 4644
rect 26421 4607 26479 4613
rect 26421 4604 26433 4607
rect 26384 4576 26433 4604
rect 26384 4564 26390 4576
rect 26421 4573 26433 4576
rect 26467 4573 26479 4607
rect 26421 4567 26479 4573
rect 26605 4607 26663 4613
rect 26605 4573 26617 4607
rect 26651 4573 26663 4607
rect 26605 4567 26663 4573
rect 26697 4607 26755 4613
rect 26697 4573 26709 4607
rect 26743 4604 26755 4607
rect 27614 4604 27620 4616
rect 26743 4576 27620 4604
rect 26743 4573 26755 4576
rect 26697 4567 26755 4573
rect 27614 4564 27620 4576
rect 27672 4564 27678 4616
rect 30374 4604 30380 4616
rect 30335 4576 30380 4604
rect 30374 4564 30380 4576
rect 30432 4564 30438 4616
rect 31018 4604 31024 4616
rect 30979 4576 31024 4604
rect 31018 4564 31024 4576
rect 31076 4564 31082 4616
rect 33244 4613 33272 4644
rect 32125 4607 32183 4613
rect 32125 4604 32137 4607
rect 31726 4576 32137 4604
rect 20990 4536 20996 4548
rect 19904 4508 20996 4536
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 26786 4536 26792 4548
rect 22066 4508 26792 4536
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 10008 4440 10149 4468
rect 10008 4428 10014 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 12805 4471 12863 4477
rect 12805 4468 12817 4471
rect 12400 4440 12817 4468
rect 12400 4428 12406 4440
rect 12805 4437 12817 4440
rect 12851 4437 12863 4471
rect 12805 4431 12863 4437
rect 13541 4471 13599 4477
rect 13541 4437 13553 4471
rect 13587 4468 13599 4471
rect 13906 4468 13912 4480
rect 13587 4440 13912 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 14921 4471 14979 4477
rect 14921 4468 14933 4471
rect 14516 4440 14933 4468
rect 14516 4428 14522 4440
rect 14921 4437 14933 4440
rect 14967 4437 14979 4471
rect 14921 4431 14979 4437
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 15528 4440 15577 4468
rect 15528 4428 15534 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 15565 4431 15623 4437
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16264 4440 16405 4468
rect 16264 4428 16270 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 17586 4468 17592 4480
rect 17547 4440 17592 4468
rect 16393 4431 16451 4437
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 18141 4471 18199 4477
rect 18141 4468 18153 4471
rect 18104 4440 18153 4468
rect 18104 4428 18110 4440
rect 18141 4437 18153 4440
rect 18187 4437 18199 4471
rect 18141 4431 18199 4437
rect 19613 4471 19671 4477
rect 19613 4437 19625 4471
rect 19659 4468 19671 4471
rect 20162 4468 20168 4480
rect 19659 4440 20168 4468
rect 19659 4437 19671 4440
rect 19613 4431 19671 4437
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 20530 4468 20536 4480
rect 20303 4440 20536 4468
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 21729 4471 21787 4477
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 22066 4468 22094 4508
rect 26786 4496 26792 4508
rect 26844 4496 26850 4548
rect 27154 4496 27160 4548
rect 27212 4536 27218 4548
rect 28537 4539 28595 4545
rect 28537 4536 28549 4539
rect 27212 4508 28549 4536
rect 27212 4496 27218 4508
rect 28537 4505 28549 4508
rect 28583 4505 28595 4539
rect 28537 4499 28595 4505
rect 28718 4496 28724 4548
rect 28776 4536 28782 4548
rect 31726 4536 31754 4576
rect 32125 4573 32137 4576
rect 32171 4573 32183 4607
rect 32125 4567 32183 4573
rect 33229 4607 33287 4613
rect 33229 4573 33241 4607
rect 33275 4573 33287 4607
rect 33962 4604 33968 4616
rect 33923 4576 33968 4604
rect 33229 4567 33287 4573
rect 33962 4564 33968 4576
rect 34020 4564 34026 4616
rect 36078 4604 36084 4616
rect 36039 4576 36084 4604
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 37090 4564 37096 4616
rect 37148 4604 37154 4616
rect 38105 4607 38163 4613
rect 38105 4604 38117 4607
rect 37148 4576 38117 4604
rect 37148 4564 37154 4576
rect 38105 4573 38117 4576
rect 38151 4573 38163 4607
rect 38105 4567 38163 4573
rect 28776 4508 31754 4536
rect 28776 4496 28782 4508
rect 33502 4496 33508 4548
rect 33560 4536 33566 4548
rect 35161 4539 35219 4545
rect 35161 4536 35173 4539
rect 33560 4508 35173 4536
rect 33560 4496 33566 4508
rect 35161 4505 35173 4508
rect 35207 4505 35219 4539
rect 37182 4536 37188 4548
rect 37143 4508 37188 4536
rect 35161 4499 35219 4505
rect 37182 4496 37188 4508
rect 37240 4496 37246 4548
rect 37274 4496 37280 4548
rect 37332 4536 37338 4548
rect 37369 4539 37427 4545
rect 37369 4536 37381 4539
rect 37332 4508 37381 4536
rect 37332 4496 37338 4508
rect 37369 4505 37381 4508
rect 37415 4536 37427 4539
rect 37918 4536 37924 4548
rect 37415 4508 37924 4536
rect 37415 4505 37427 4508
rect 37369 4499 37427 4505
rect 37918 4496 37924 4508
rect 37976 4496 37982 4548
rect 21775 4440 22094 4468
rect 22373 4471 22431 4477
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 22373 4437 22385 4471
rect 22419 4468 22431 4471
rect 22738 4468 22744 4480
rect 22419 4440 22744 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 22738 4428 22744 4440
rect 22796 4428 22802 4480
rect 22922 4468 22928 4480
rect 22883 4440 22928 4468
rect 22922 4428 22928 4440
rect 22980 4428 22986 4480
rect 23750 4468 23756 4480
rect 23711 4440 23756 4468
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 24578 4468 24584 4480
rect 24539 4440 24584 4468
rect 24578 4428 24584 4440
rect 24636 4428 24642 4480
rect 26326 4428 26332 4480
rect 26384 4468 26390 4480
rect 27430 4468 27436 4480
rect 26384 4440 27436 4468
rect 26384 4428 26390 4440
rect 27430 4428 27436 4440
rect 27488 4428 27494 4480
rect 29641 4471 29699 4477
rect 29641 4437 29653 4471
rect 29687 4468 29699 4471
rect 29822 4468 29828 4480
rect 29687 4440 29828 4468
rect 29687 4437 29699 4440
rect 29641 4431 29699 4437
rect 29822 4428 29828 4440
rect 29880 4428 29886 4480
rect 30190 4428 30196 4480
rect 30248 4468 30254 4480
rect 31205 4471 31263 4477
rect 31205 4468 31217 4471
rect 30248 4440 31217 4468
rect 30248 4428 30254 4440
rect 31205 4437 31217 4440
rect 31251 4437 31263 4471
rect 34146 4468 34152 4480
rect 34107 4440 34152 4468
rect 31205 4431 31263 4437
rect 34146 4428 34152 4440
rect 34204 4428 34210 4480
rect 35986 4428 35992 4480
rect 36044 4468 36050 4480
rect 36265 4471 36323 4477
rect 36265 4468 36277 4471
rect 36044 4440 36277 4468
rect 36044 4428 36050 4440
rect 36265 4437 36277 4440
rect 36311 4437 36323 4471
rect 36265 4431 36323 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2777 4267 2835 4273
rect 2777 4233 2789 4267
rect 2823 4264 2835 4267
rect 3878 4264 3884 4276
rect 2823 4236 3884 4264
rect 2823 4233 2835 4236
rect 2777 4227 2835 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 10137 4267 10195 4273
rect 10137 4264 10149 4267
rect 8536 4236 10149 4264
rect 8536 4224 8542 4236
rect 10137 4233 10149 4236
rect 10183 4233 10195 4267
rect 10137 4227 10195 4233
rect 12250 4224 12256 4276
rect 12308 4264 12314 4276
rect 12345 4267 12403 4273
rect 12345 4264 12357 4267
rect 12308 4236 12357 4264
rect 12308 4224 12314 4236
rect 12345 4233 12357 4236
rect 12391 4233 12403 4267
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 12345 4227 12403 4233
rect 15856 4236 19257 4264
rect 5074 4196 5080 4208
rect 4172 4168 5080 4196
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 624 4100 1409 4128
rect 624 4088 630 4100
rect 1397 4097 1409 4100
rect 1443 4128 1455 4131
rect 1946 4128 1952 4140
rect 1443 4100 1952 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 2924 4100 2969 4128
rect 2924 4088 2930 4100
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 3292 4100 3617 4128
rect 3292 4088 3298 4100
rect 3605 4097 3617 4100
rect 3651 4128 3663 4131
rect 4172 4128 4200 4168
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 5626 4196 5632 4208
rect 5368 4168 5632 4196
rect 3651 4100 4200 4128
rect 4249 4131 4307 4137
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4798 4128 4804 4140
rect 4295 4100 4804 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 290 4020 296 4072
rect 348 4060 354 4072
rect 1578 4060 1584 4072
rect 348 4032 1584 4060
rect 348 4020 354 4032
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 3050 4060 3056 4072
rect 3011 4032 3056 4060
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 4264 4060 4292 4091
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5368 4128 5396 4168
rect 5626 4156 5632 4168
rect 5684 4156 5690 4208
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 7469 4199 7527 4205
rect 7469 4196 7481 4199
rect 7248 4168 7481 4196
rect 7248 4156 7254 4168
rect 7469 4165 7481 4168
rect 7515 4165 7527 4199
rect 7469 4159 7527 4165
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 15856 4196 15884 4236
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 20530 4264 20536 4276
rect 20491 4236 20536 4264
rect 19245 4227 19303 4233
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 20916 4196 20944 4227
rect 20990 4224 20996 4276
rect 21048 4264 21054 4276
rect 21910 4264 21916 4276
rect 21048 4236 21916 4264
rect 21048 4224 21054 4236
rect 21910 4224 21916 4236
rect 21968 4264 21974 4276
rect 24489 4267 24547 4273
rect 24489 4264 24501 4267
rect 21968 4236 24501 4264
rect 21968 4224 21974 4236
rect 24489 4233 24501 4236
rect 24535 4264 24547 4267
rect 24578 4264 24584 4276
rect 24535 4236 24584 4264
rect 24535 4233 24547 4236
rect 24489 4227 24547 4233
rect 24578 4224 24584 4236
rect 24636 4224 24642 4276
rect 25958 4224 25964 4276
rect 26016 4264 26022 4276
rect 27614 4264 27620 4276
rect 26016 4236 27200 4264
rect 27575 4236 27620 4264
rect 26016 4224 26022 4236
rect 27062 4196 27068 4208
rect 8168 4168 15884 4196
rect 19168 4168 19472 4196
rect 20916 4168 27068 4196
rect 8168 4156 8174 4168
rect 4948 4100 5396 4128
rect 4948 4088 4954 4100
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5500 4100 5549 4128
rect 5500 4088 5506 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 6420 4100 6469 4128
rect 6420 4088 6426 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 11330 4128 11336 4140
rect 8987 4100 11336 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11756 4100 11897 4128
rect 11756 4088 11762 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12526 4128 12532 4140
rect 12032 4100 12532 4128
rect 12032 4088 12038 4100
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13722 4128 13728 4140
rect 13683 4100 13728 4128
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 16114 4128 16120 4140
rect 15519 4100 16120 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 7558 4060 7564 4072
rect 3620 4032 4292 4060
rect 4448 4032 7564 4060
rect 3620 4004 3648 4032
rect 2406 3992 2412 4004
rect 2367 3964 2412 3992
rect 2406 3952 2412 3964
rect 2464 3952 2470 4004
rect 3602 3952 3608 4004
rect 3660 3952 3666 4004
rect 4448 4001 4476 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8478 4060 8484 4072
rect 7699 4032 8484 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8628 4032 8677 4060
rect 8628 4020 8634 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10042 4060 10048 4072
rect 9732 4032 10048 4060
rect 9732 4020 9738 4032
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 12250 4060 12256 4072
rect 10275 4032 12256 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 14752 4060 14780 4091
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4128 17463 4131
rect 19168 4128 19196 4168
rect 19334 4128 19340 4140
rect 17451 4100 19196 4128
rect 19295 4100 19340 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19444 4128 19472 4168
rect 27062 4156 27068 4168
rect 27120 4156 27126 4208
rect 27172 4196 27200 4236
rect 27614 4224 27620 4236
rect 27672 4224 27678 4276
rect 28258 4224 28264 4276
rect 28316 4264 28322 4276
rect 28316 4236 30328 4264
rect 28316 4224 28322 4236
rect 27172 4168 27568 4196
rect 27540 4140 27568 4168
rect 22278 4128 22284 4140
rect 19444 4100 22284 4128
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4128 22431 4131
rect 23014 4128 23020 4140
rect 22419 4100 23020 4128
rect 22419 4097 22431 4100
rect 22373 4091 22431 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 24026 4128 24032 4140
rect 23987 4100 24032 4128
rect 24026 4088 24032 4100
rect 24084 4088 24090 4140
rect 25225 4131 25283 4137
rect 25225 4097 25237 4131
rect 25271 4128 25283 4131
rect 27157 4131 27215 4137
rect 25271 4100 26188 4128
rect 25271 4097 25283 4100
rect 25225 4091 25283 4097
rect 15562 4060 15568 4072
rect 12406 4032 14688 4060
rect 14752 4032 15568 4060
rect 4433 3995 4491 4001
rect 4433 3961 4445 3995
rect 4479 3961 4491 3995
rect 5626 3992 5632 4004
rect 4433 3955 4491 3961
rect 4908 3964 5632 3992
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2774 3924 2780 3936
rect 1627 3896 2780 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3789 3927 3847 3933
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 4908 3924 4936 3964
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 5721 3995 5779 4001
rect 5721 3961 5733 3995
rect 5767 3992 5779 3995
rect 7926 3992 7932 4004
rect 5767 3964 7932 3992
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 7926 3952 7932 3964
rect 7984 3952 7990 4004
rect 10594 3992 10600 4004
rect 10555 3964 10600 3992
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 11701 3995 11759 4001
rect 11701 3992 11713 3995
rect 11480 3964 11713 3992
rect 11480 3952 11486 3964
rect 11701 3961 11713 3964
rect 11747 3961 11759 3995
rect 12406 3992 12434 4032
rect 11701 3955 11759 3961
rect 12084 3964 12434 3992
rect 5074 3924 5080 3936
rect 3835 3896 4936 3924
rect 5035 3896 5080 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5534 3924 5540 3936
rect 5408 3896 5540 3924
rect 5408 3884 5414 3896
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6638 3924 6644 3936
rect 6599 3896 6644 3924
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 12084 3924 12112 3964
rect 12986 3952 12992 4004
rect 13044 3992 13050 4004
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 13044 3964 13921 3992
rect 13044 3952 13050 3964
rect 13909 3961 13921 3964
rect 13955 3961 13967 3995
rect 14660 3992 14688 4032
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 19058 4060 19064 4072
rect 19019 4032 19064 4060
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19886 4020 19892 4072
rect 19944 4060 19950 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19944 4032 20269 4060
rect 19944 4020 19950 4032
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20438 4060 20444 4072
rect 20399 4032 20444 4060
rect 20257 4023 20315 4029
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 22646 4060 22652 4072
rect 20916 4032 22652 4060
rect 15838 3992 15844 4004
rect 14660 3964 15844 3992
rect 13909 3955 13967 3961
rect 15838 3952 15844 3964
rect 15896 3952 15902 4004
rect 17310 3952 17316 4004
rect 17368 3992 17374 4004
rect 17957 3995 18015 4001
rect 17957 3992 17969 3995
rect 17368 3964 17969 3992
rect 17368 3952 17374 3964
rect 17957 3961 17969 3964
rect 18003 3992 18015 3995
rect 19705 3995 19763 4001
rect 18003 3964 18644 3992
rect 18003 3961 18015 3964
rect 17957 3955 18015 3961
rect 11020 3896 12112 3924
rect 11020 3884 11026 3896
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12216 3896 13185 3924
rect 12216 3884 12222 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 13173 3887 13231 3893
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 13780 3896 14565 3924
rect 13780 3884 13786 3896
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14553 3887 14611 3893
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 14792 3896 15301 3924
rect 14792 3884 14798 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 15289 3887 15347 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 17092 3896 17233 3924
rect 17092 3884 17098 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18196 3896 18429 3924
rect 18196 3884 18202 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18616 3924 18644 3964
rect 19705 3961 19717 3995
rect 19751 3992 19763 3995
rect 20806 3992 20812 4004
rect 19751 3964 20812 3992
rect 19751 3961 19763 3964
rect 19705 3955 19763 3961
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 20916 3924 20944 4032
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 24578 4020 24584 4072
rect 24636 4060 24642 4072
rect 25314 4060 25320 4072
rect 24636 4032 25320 4060
rect 24636 4020 24642 4032
rect 25314 4020 25320 4032
rect 25372 4060 25378 4072
rect 26160 4069 26188 4100
rect 27157 4097 27169 4131
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 25685 4063 25743 4069
rect 25685 4060 25697 4063
rect 25372 4032 25697 4060
rect 25372 4020 25378 4032
rect 25685 4029 25697 4032
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 26145 4063 26203 4069
rect 26145 4029 26157 4063
rect 26191 4029 26203 4063
rect 26145 4023 26203 4029
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 25041 3995 25099 4001
rect 25041 3992 25053 3995
rect 21048 3964 25053 3992
rect 21048 3952 21054 3964
rect 25041 3961 25053 3964
rect 25087 3961 25099 3995
rect 26050 3992 26056 4004
rect 26011 3964 26056 3992
rect 25041 3955 25099 3961
rect 26050 3952 26056 3964
rect 26108 3952 26114 4004
rect 26970 3992 26976 4004
rect 26931 3964 26976 3992
rect 26970 3952 26976 3964
rect 27028 3952 27034 4004
rect 18616 3896 20944 3924
rect 18417 3887 18475 3893
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22189 3927 22247 3933
rect 22189 3924 22201 3927
rect 22060 3896 22201 3924
rect 22060 3884 22066 3896
rect 22189 3893 22201 3896
rect 22235 3893 22247 3927
rect 22189 3887 22247 3893
rect 22830 3884 22836 3936
rect 22888 3924 22894 3936
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22888 3896 23029 3924
rect 22888 3884 22894 3896
rect 23017 3893 23029 3896
rect 23063 3893 23075 3927
rect 23017 3887 23075 3893
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 23716 3896 23857 3924
rect 23716 3884 23722 3896
rect 23845 3893 23857 3896
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 25774 3884 25780 3936
rect 25832 3924 25838 3936
rect 27172 3924 27200 4091
rect 27522 4088 27528 4140
rect 27580 4128 27586 4140
rect 27801 4131 27859 4137
rect 27801 4128 27813 4131
rect 27580 4100 27813 4128
rect 27580 4088 27586 4100
rect 27801 4097 27813 4100
rect 27847 4097 27859 4131
rect 28626 4128 28632 4140
rect 28587 4100 28632 4128
rect 27801 4091 27859 4097
rect 28626 4088 28632 4100
rect 28684 4088 28690 4140
rect 29362 4088 29368 4140
rect 29420 4128 29426 4140
rect 30300 4128 30328 4236
rect 30374 4224 30380 4276
rect 30432 4264 30438 4276
rect 31478 4264 31484 4276
rect 30432 4236 31484 4264
rect 30432 4224 30438 4236
rect 31478 4224 31484 4236
rect 31536 4224 31542 4276
rect 31662 4224 31668 4276
rect 31720 4264 31726 4276
rect 34238 4264 34244 4276
rect 31720 4236 34244 4264
rect 31720 4224 31726 4236
rect 34238 4224 34244 4236
rect 34296 4224 34302 4276
rect 30926 4196 30932 4208
rect 30576 4168 30932 4196
rect 30469 4131 30527 4137
rect 30469 4128 30481 4131
rect 29420 4100 29960 4128
rect 30300 4100 30481 4128
rect 29420 4088 29426 4100
rect 29822 4060 29828 4072
rect 29783 4032 29828 4060
rect 29822 4020 29828 4032
rect 29880 4020 29886 4072
rect 29932 4060 29960 4100
rect 30469 4097 30481 4100
rect 30515 4128 30527 4131
rect 30576 4128 30604 4168
rect 30926 4156 30932 4168
rect 30984 4156 30990 4208
rect 33796 4168 34100 4196
rect 30515 4100 30604 4128
rect 30515 4097 30527 4100
rect 30469 4091 30527 4097
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 31021 4131 31079 4137
rect 31021 4128 31033 4131
rect 30800 4100 31033 4128
rect 30800 4088 30806 4100
rect 31021 4097 31033 4100
rect 31067 4097 31079 4131
rect 31021 4091 31079 4097
rect 32125 4131 32183 4137
rect 32125 4097 32137 4131
rect 32171 4128 32183 4131
rect 32214 4128 32220 4140
rect 32171 4100 32220 4128
rect 32171 4097 32183 4100
rect 32125 4091 32183 4097
rect 32214 4088 32220 4100
rect 32272 4088 32278 4140
rect 32306 4088 32312 4140
rect 32364 4128 32370 4140
rect 32861 4131 32919 4137
rect 32861 4128 32873 4131
rect 32364 4100 32873 4128
rect 32364 4088 32370 4100
rect 32861 4097 32873 4100
rect 32907 4097 32919 4131
rect 33796 4128 33824 4168
rect 33962 4128 33968 4140
rect 32861 4091 32919 4097
rect 32968 4100 33824 4128
rect 33923 4100 33968 4128
rect 29932 4032 31248 4060
rect 29457 3995 29515 4001
rect 29457 3961 29469 3995
rect 29503 3961 29515 3995
rect 29457 3955 29515 3961
rect 25832 3896 27200 3924
rect 25832 3884 25838 3896
rect 28534 3884 28540 3936
rect 28592 3924 28598 3936
rect 28813 3927 28871 3933
rect 28813 3924 28825 3927
rect 28592 3896 28825 3924
rect 28592 3884 28598 3896
rect 28813 3893 28825 3896
rect 28859 3893 28871 3927
rect 28813 3887 28871 3893
rect 28994 3884 29000 3936
rect 29052 3924 29058 3936
rect 29365 3927 29423 3933
rect 29365 3924 29377 3927
rect 29052 3896 29377 3924
rect 29052 3884 29058 3896
rect 29365 3893 29377 3896
rect 29411 3893 29423 3927
rect 29472 3924 29500 3955
rect 29546 3952 29552 4004
rect 29604 3992 29610 4004
rect 31220 4001 31248 4032
rect 30285 3995 30343 4001
rect 30285 3992 30297 3995
rect 29604 3964 30297 3992
rect 29604 3952 29610 3964
rect 30285 3961 30297 3964
rect 30331 3961 30343 3995
rect 30285 3955 30343 3961
rect 31205 3995 31263 4001
rect 31205 3961 31217 3995
rect 31251 3961 31263 3995
rect 31205 3955 31263 3961
rect 32214 3952 32220 4004
rect 32272 3992 32278 4004
rect 32968 3992 32996 4100
rect 33962 4088 33968 4100
rect 34020 4088 34026 4140
rect 33134 4020 33140 4072
rect 33192 4060 33198 4072
rect 34072 4060 34100 4168
rect 36262 4156 36268 4208
rect 36320 4196 36326 4208
rect 36541 4199 36599 4205
rect 36541 4196 36553 4199
rect 36320 4168 36553 4196
rect 36320 4156 36326 4168
rect 36541 4165 36553 4168
rect 36587 4165 36599 4199
rect 36541 4159 36599 4165
rect 34146 4088 34152 4140
rect 34204 4128 34210 4140
rect 35253 4131 35311 4137
rect 35253 4128 35265 4131
rect 34204 4100 35265 4128
rect 34204 4088 34210 4100
rect 35253 4097 35265 4100
rect 35299 4097 35311 4131
rect 37274 4128 37280 4140
rect 37235 4100 37280 4128
rect 35253 4091 35311 4097
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 38105 4131 38163 4137
rect 38105 4097 38117 4131
rect 38151 4128 38163 4131
rect 38378 4128 38384 4140
rect 38151 4100 38384 4128
rect 38151 4097 38163 4100
rect 38105 4091 38163 4097
rect 38378 4088 38384 4100
rect 38436 4088 38442 4140
rect 33192 4032 34008 4060
rect 34072 4032 34744 4060
rect 33192 4020 33198 4032
rect 32272 3964 32996 3992
rect 32272 3952 32278 3964
rect 30650 3924 30656 3936
rect 29472 3896 30656 3924
rect 29365 3887 29423 3893
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 31846 3884 31852 3936
rect 31904 3924 31910 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 31904 3896 32321 3924
rect 31904 3884 31910 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 32309 3887 32367 3893
rect 33045 3927 33103 3933
rect 33045 3893 33057 3927
rect 33091 3924 33103 3927
rect 33778 3924 33784 3936
rect 33091 3896 33784 3924
rect 33091 3893 33103 3896
rect 33045 3887 33103 3893
rect 33778 3884 33784 3896
rect 33836 3884 33842 3936
rect 33980 3924 34008 4032
rect 34716 4001 34744 4032
rect 34701 3995 34759 4001
rect 34701 3961 34713 3995
rect 34747 3961 34759 3995
rect 34701 3955 34759 3961
rect 37461 3995 37519 4001
rect 37461 3961 37473 3995
rect 37507 3992 37519 3995
rect 38654 3992 38660 4004
rect 37507 3964 38660 3992
rect 37507 3961 37519 3964
rect 37461 3955 37519 3961
rect 38654 3952 38660 3964
rect 38712 3952 38718 4004
rect 34149 3927 34207 3933
rect 34149 3924 34161 3927
rect 33980 3896 34161 3924
rect 34149 3893 34161 3896
rect 34195 3893 34207 3927
rect 34149 3887 34207 3893
rect 34422 3884 34428 3936
rect 34480 3924 34486 3936
rect 34790 3924 34796 3936
rect 34480 3896 34796 3924
rect 34480 3884 34486 3896
rect 34790 3884 34796 3896
rect 34848 3884 34854 3936
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 35437 3927 35495 3933
rect 35437 3924 35449 3927
rect 35400 3896 35449 3924
rect 35400 3884 35406 3896
rect 35437 3893 35449 3896
rect 35483 3893 35495 3927
rect 36446 3924 36452 3936
rect 36407 3896 36452 3924
rect 35437 3887 35495 3893
rect 36446 3884 36452 3896
rect 36504 3884 36510 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 4982 3720 4988 3732
rect 4943 3692 4988 3720
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 6178 3720 6184 3732
rect 6139 3692 6184 3720
rect 6178 3680 6184 3692
rect 6236 3680 6242 3732
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 11514 3720 11520 3732
rect 7616 3692 11376 3720
rect 11475 3692 11520 3720
rect 7616 3680 7622 3692
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 3142 3652 3148 3664
rect 2004 3624 3148 3652
rect 2004 3612 2010 3624
rect 3142 3612 3148 3624
rect 3200 3652 3206 3664
rect 3973 3655 4031 3661
rect 3200 3624 3832 3652
rect 3200 3612 3206 3624
rect 842 3544 848 3596
rect 900 3584 906 3596
rect 2958 3584 2964 3596
rect 900 3556 2964 3584
rect 900 3544 906 3556
rect 2958 3544 2964 3556
rect 3016 3584 3022 3596
rect 3016 3556 3280 3584
rect 3016 3544 3022 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 3252 3525 3280 3556
rect 3804 3525 3832 3624
rect 3973 3621 3985 3655
rect 4019 3652 4031 3655
rect 7745 3655 7803 3661
rect 4019 3624 6684 3652
rect 4019 3621 4031 3624
rect 3973 3615 4031 3621
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5224 3556 5457 3584
rect 5224 3544 5230 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 6656 3593 6684 3624
rect 7745 3621 7757 3655
rect 7791 3652 7803 3655
rect 8294 3652 8300 3664
rect 7791 3624 8300 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 11348 3652 11376 3692
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 13170 3720 13176 3732
rect 13131 3692 13176 3720
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13998 3680 14004 3732
rect 14056 3720 14062 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 14056 3692 14105 3720
rect 14056 3680 14062 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 16942 3720 16948 3732
rect 16903 3692 16948 3720
rect 14093 3683 14151 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 19334 3720 19340 3732
rect 19295 3692 19340 3720
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 19981 3723 20039 3729
rect 19981 3720 19993 3723
rect 19944 3692 19993 3720
rect 19944 3680 19950 3692
rect 19981 3689 19993 3692
rect 20027 3720 20039 3723
rect 20530 3720 20536 3732
rect 20027 3692 20536 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 22557 3723 22615 3729
rect 22557 3689 22569 3723
rect 22603 3720 22615 3723
rect 23382 3720 23388 3732
rect 22603 3692 23388 3720
rect 22603 3689 22615 3692
rect 22557 3683 22615 3689
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 23934 3720 23940 3732
rect 23799 3692 23940 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 23934 3680 23940 3692
rect 23992 3680 23998 3732
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 36446 3720 36452 3732
rect 24084 3692 36452 3720
rect 24084 3680 24090 3692
rect 36446 3680 36452 3692
rect 36504 3680 36510 3732
rect 16485 3655 16543 3661
rect 11348 3624 16068 3652
rect 6641 3587 6699 3593
rect 5592 3556 5685 3584
rect 5592 3544 5598 3556
rect 6641 3553 6653 3587
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6788 3556 6881 3584
rect 6788 3544 6794 3556
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 9769 3587 9827 3593
rect 8444 3556 9720 3584
rect 8444 3544 8450 3556
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1728 3488 1777 3516
rect 1728 3476 1734 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 3237 3519 3295 3525
rect 2087 3488 3188 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 3016 3352 3065 3380
rect 3016 3340 3022 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3160 3380 3188 3488
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4430 3476 4436 3528
rect 4488 3516 4494 3528
rect 5552 3516 5580 3544
rect 6748 3516 6776 3544
rect 4488 3488 5580 3516
rect 6472 3488 6776 3516
rect 4488 3476 4494 3488
rect 4522 3448 4528 3460
rect 4483 3420 4528 3448
rect 4522 3408 4528 3420
rect 4580 3408 4586 3460
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 6086 3448 6092 3460
rect 5399 3420 6092 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 6472 3380 6500 3488
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 8202 3516 8208 3528
rect 7524 3488 8208 3516
rect 7524 3476 7530 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9692 3516 9720 3556
rect 9769 3553 9781 3587
rect 9815 3584 9827 3587
rect 9858 3584 9864 3596
rect 9815 3556 9864 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 10836 3556 12480 3584
rect 10836 3544 10842 3556
rect 11241 3519 11299 3525
rect 9692 3488 11100 3516
rect 9493 3479 9551 3485
rect 6549 3451 6607 3457
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 6595 3420 6776 3448
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 3160 3352 6500 3380
rect 6748 3380 6776 3420
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 6880 3420 7573 3448
rect 6880 3408 6886 3420
rect 7561 3417 7573 3420
rect 7607 3448 7619 3451
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 7607 3420 8953 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 8941 3417 8953 3420
rect 8987 3417 8999 3451
rect 8941 3411 8999 3417
rect 9858 3408 9864 3460
rect 9916 3448 9922 3460
rect 10870 3448 10876 3460
rect 9916 3420 10876 3448
rect 9916 3408 9922 3420
rect 10870 3408 10876 3420
rect 10928 3448 10934 3460
rect 10965 3451 11023 3457
rect 10965 3448 10977 3451
rect 10928 3420 10977 3448
rect 10928 3408 10934 3420
rect 10965 3417 10977 3420
rect 11011 3417 11023 3451
rect 11072 3448 11100 3488
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 12342 3516 12348 3528
rect 11287 3488 12348 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12452 3516 12480 3556
rect 12526 3544 12532 3596
rect 12584 3584 12590 3596
rect 12584 3556 12629 3584
rect 12584 3544 12590 3556
rect 14182 3544 14188 3596
rect 14240 3584 14246 3596
rect 14645 3587 14703 3593
rect 14645 3584 14657 3587
rect 14240 3556 14657 3584
rect 14240 3544 14246 3556
rect 14645 3553 14657 3556
rect 14691 3553 14703 3587
rect 15838 3584 15844 3596
rect 15799 3556 15844 3584
rect 14645 3547 14703 3553
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16040 3593 16068 3624
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 17126 3652 17132 3664
rect 16531 3624 17132 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 26234 3652 26240 3664
rect 17420 3624 26240 3652
rect 16025 3587 16083 3593
rect 16025 3553 16037 3587
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 17420 3584 17448 3624
rect 26234 3612 26240 3624
rect 26292 3612 26298 3664
rect 28350 3652 28356 3664
rect 26344 3624 28356 3652
rect 16356 3556 17448 3584
rect 16356 3544 16362 3556
rect 17494 3544 17500 3596
rect 17552 3584 17558 3596
rect 21910 3584 21916 3596
rect 17552 3556 17597 3584
rect 21871 3556 21916 3584
rect 17552 3544 17558 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 22094 3584 22100 3596
rect 22055 3556 22100 3584
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 23014 3544 23020 3596
rect 23072 3584 23078 3596
rect 23109 3587 23167 3593
rect 23109 3584 23121 3587
rect 23072 3556 23121 3584
rect 23072 3544 23078 3556
rect 23109 3553 23121 3556
rect 23155 3584 23167 3587
rect 26344 3584 26372 3624
rect 28350 3612 28356 3624
rect 28408 3652 28414 3664
rect 29822 3652 29828 3664
rect 28408 3624 29828 3652
rect 28408 3612 28414 3624
rect 23155 3556 26372 3584
rect 23155 3553 23167 3556
rect 23109 3547 23167 3553
rect 26418 3544 26424 3596
rect 26476 3584 26482 3596
rect 26476 3556 27016 3584
rect 26476 3544 26482 3556
rect 14553 3519 14611 3525
rect 14553 3516 14565 3519
rect 12452 3488 14565 3516
rect 14553 3485 14565 3488
rect 14599 3485 14611 3519
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 14553 3479 14611 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 17310 3516 17316 3528
rect 17271 3488 17316 3516
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 18414 3516 18420 3528
rect 18375 3488 18420 3516
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19242 3516 19248 3528
rect 19024 3488 19248 3516
rect 19024 3476 19030 3488
rect 19242 3476 19248 3488
rect 19300 3516 19306 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19300 3488 19533 3516
rect 19300 3476 19306 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20404 3488 20545 3516
rect 20404 3476 20410 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21174 3516 21180 3528
rect 20680 3488 21180 3516
rect 20680 3476 20686 3488
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 22186 3516 22192 3528
rect 22147 3488 22192 3516
rect 22186 3476 22192 3488
rect 22244 3476 22250 3528
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 22796 3488 23397 3516
rect 22796 3476 22802 3488
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 23385 3479 23443 3485
rect 23492 3488 25237 3516
rect 11072 3420 11192 3448
rect 10965 3411 11023 3417
rect 7650 3380 7656 3392
rect 6748 3352 7656 3380
rect 3053 3343 3111 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8386 3380 8392 3392
rect 8347 3352 8392 3380
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 11054 3380 11060 3392
rect 11015 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 11164 3380 11192 3420
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 14458 3448 14464 3460
rect 11480 3420 14320 3448
rect 14419 3420 14464 3448
rect 11480 3408 11486 3420
rect 12713 3383 12771 3389
rect 12713 3380 12725 3383
rect 11164 3352 12725 3380
rect 12713 3349 12725 3352
rect 12759 3349 12771 3383
rect 12713 3343 12771 3349
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 14292 3380 14320 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 17405 3451 17463 3457
rect 17405 3448 17417 3451
rect 14752 3420 17417 3448
rect 14752 3380 14780 3420
rect 17405 3417 17417 3420
rect 17451 3417 17463 3451
rect 23492 3448 23520 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 25372 3488 25421 3516
rect 25372 3476 25378 3488
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 26510 3516 26516 3528
rect 26471 3488 26516 3516
rect 25409 3479 25467 3485
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 26988 3525 27016 3556
rect 26973 3519 27031 3525
rect 26973 3485 26985 3519
rect 27019 3485 27031 3519
rect 27798 3516 27804 3528
rect 27759 3488 27804 3516
rect 26973 3479 27031 3485
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28828 3525 28856 3624
rect 29822 3612 29828 3624
rect 29880 3612 29886 3664
rect 31570 3652 31576 3664
rect 31531 3624 31576 3652
rect 31570 3612 31576 3624
rect 31628 3612 31634 3664
rect 31956 3624 32168 3652
rect 30282 3584 30288 3596
rect 28920 3556 30144 3584
rect 30243 3556 30288 3584
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 17405 3411 17463 3417
rect 22066 3420 23520 3448
rect 12860 3352 12905 3380
rect 14292 3352 14780 3380
rect 12860 3340 12866 3352
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17920 3352 18245 3380
rect 17920 3340 17926 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 21361 3383 21419 3389
rect 21361 3349 21373 3383
rect 21407 3380 21419 3383
rect 22066 3380 22094 3420
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 24581 3451 24639 3457
rect 24581 3448 24593 3451
rect 24268 3420 24593 3448
rect 24268 3408 24274 3420
rect 24581 3417 24593 3420
rect 24627 3417 24639 3451
rect 24762 3448 24768 3460
rect 24723 3420 24768 3448
rect 24581 3411 24639 3417
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 26786 3408 26792 3460
rect 26844 3448 26850 3460
rect 28629 3451 28687 3457
rect 28629 3448 28641 3451
rect 26844 3420 28641 3448
rect 26844 3408 26850 3420
rect 28629 3417 28641 3420
rect 28675 3417 28687 3451
rect 28629 3411 28687 3417
rect 23290 3380 23296 3392
rect 21407 3352 22094 3380
rect 23251 3352 23296 3380
rect 21407 3349 21419 3352
rect 21361 3343 21419 3349
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 25590 3380 25596 3392
rect 25551 3352 25596 3380
rect 25590 3340 25596 3352
rect 25648 3340 25654 3392
rect 26050 3340 26056 3392
rect 26108 3380 26114 3392
rect 26329 3383 26387 3389
rect 26329 3380 26341 3383
rect 26108 3352 26341 3380
rect 26108 3340 26114 3352
rect 26329 3349 26341 3352
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 26878 3340 26884 3392
rect 26936 3380 26942 3392
rect 27157 3383 27215 3389
rect 27157 3380 27169 3383
rect 26936 3352 27169 3380
rect 26936 3340 26942 3352
rect 27157 3349 27169 3352
rect 27203 3349 27215 3383
rect 27157 3343 27215 3349
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 27985 3383 28043 3389
rect 27985 3380 27997 3383
rect 27764 3352 27997 3380
rect 27764 3340 27770 3352
rect 27985 3349 27997 3352
rect 28031 3349 28043 3383
rect 27985 3343 28043 3349
rect 28166 3340 28172 3392
rect 28224 3380 28230 3392
rect 28920 3380 28948 3556
rect 29914 3476 29920 3528
rect 29972 3516 29978 3528
rect 30009 3519 30067 3525
rect 30009 3516 30021 3519
rect 29972 3488 30021 3516
rect 29972 3476 29978 3488
rect 30009 3485 30021 3488
rect 30055 3485 30067 3519
rect 30116 3516 30144 3556
rect 30282 3544 30288 3556
rect 30340 3544 30346 3596
rect 31956 3584 31984 3624
rect 30392 3556 31984 3584
rect 32140 3584 32168 3624
rect 34146 3612 34152 3664
rect 34204 3652 34210 3664
rect 36173 3655 36231 3661
rect 36173 3652 36185 3655
rect 34204 3624 36185 3652
rect 34204 3612 34210 3624
rect 36173 3621 36185 3624
rect 36219 3621 36231 3655
rect 36173 3615 36231 3621
rect 37274 3584 37280 3596
rect 32140 3556 37280 3584
rect 30392 3516 30420 3556
rect 37274 3544 37280 3556
rect 37332 3544 37338 3596
rect 37642 3544 37648 3596
rect 37700 3584 37706 3596
rect 37829 3587 37887 3593
rect 37829 3584 37841 3587
rect 37700 3556 37841 3584
rect 37700 3544 37706 3556
rect 37829 3553 37841 3556
rect 37875 3553 37887 3587
rect 37829 3547 37887 3553
rect 38105 3587 38163 3593
rect 38105 3553 38117 3587
rect 38151 3584 38163 3587
rect 38194 3584 38200 3596
rect 38151 3556 38200 3584
rect 38151 3553 38163 3556
rect 38105 3547 38163 3553
rect 38194 3544 38200 3556
rect 38252 3544 38258 3596
rect 30116 3488 30420 3516
rect 30009 3479 30067 3485
rect 30742 3476 30748 3528
rect 30800 3516 30806 3528
rect 31389 3519 31447 3525
rect 31389 3516 31401 3519
rect 30800 3488 31401 3516
rect 30800 3476 30806 3488
rect 31389 3485 31401 3488
rect 31435 3516 31447 3519
rect 31754 3516 31760 3528
rect 31435 3488 31760 3516
rect 31435 3485 31447 3488
rect 31389 3479 31447 3485
rect 31754 3476 31760 3488
rect 31812 3476 31818 3528
rect 32030 3476 32036 3528
rect 32088 3516 32094 3528
rect 32769 3519 32827 3525
rect 32088 3488 32133 3516
rect 32088 3476 32094 3488
rect 32769 3485 32781 3519
rect 32815 3485 32827 3519
rect 32769 3479 32827 3485
rect 28997 3451 29055 3457
rect 28997 3417 29009 3451
rect 29043 3448 29055 3451
rect 31662 3448 31668 3460
rect 29043 3420 31668 3448
rect 29043 3417 29055 3420
rect 28997 3411 29055 3417
rect 31662 3408 31668 3420
rect 31720 3408 31726 3460
rect 31938 3408 31944 3460
rect 31996 3448 32002 3460
rect 32784 3448 32812 3479
rect 33686 3476 33692 3528
rect 33744 3516 33750 3528
rect 33873 3519 33931 3525
rect 33873 3516 33885 3519
rect 33744 3488 33885 3516
rect 33744 3476 33750 3488
rect 33873 3485 33885 3488
rect 33919 3485 33931 3519
rect 33873 3479 33931 3485
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35253 3519 35311 3525
rect 35253 3516 35265 3519
rect 34848 3488 35265 3516
rect 34848 3476 34854 3488
rect 35253 3485 35265 3488
rect 35299 3516 35311 3519
rect 35434 3516 35440 3528
rect 35299 3488 35440 3516
rect 35299 3485 35311 3488
rect 35253 3479 35311 3485
rect 35434 3476 35440 3488
rect 35492 3476 35498 3528
rect 36357 3519 36415 3525
rect 36357 3485 36369 3519
rect 36403 3516 36415 3519
rect 38378 3516 38384 3528
rect 36403 3488 38384 3516
rect 36403 3485 36415 3488
rect 36357 3479 36415 3485
rect 38378 3476 38384 3488
rect 38436 3476 38442 3528
rect 31996 3420 32812 3448
rect 31996 3408 32002 3420
rect 34514 3408 34520 3460
rect 34572 3448 34578 3460
rect 35069 3451 35127 3457
rect 35069 3448 35081 3451
rect 34572 3420 35081 3448
rect 34572 3408 34578 3420
rect 35069 3417 35081 3420
rect 35115 3417 35127 3451
rect 35069 3411 35127 3417
rect 35158 3408 35164 3460
rect 35216 3448 35222 3460
rect 38930 3448 38936 3460
rect 35216 3420 38936 3448
rect 35216 3408 35222 3420
rect 38930 3408 38936 3420
rect 38988 3408 38994 3460
rect 28224 3352 28948 3380
rect 28224 3340 28230 3352
rect 31018 3340 31024 3392
rect 31076 3380 31082 3392
rect 32217 3383 32275 3389
rect 32217 3380 32229 3383
rect 31076 3352 32229 3380
rect 31076 3340 31082 3352
rect 32217 3349 32229 3352
rect 32263 3349 32275 3383
rect 32217 3343 32275 3349
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 32953 3383 33011 3389
rect 32953 3380 32965 3383
rect 32732 3352 32965 3380
rect 32732 3340 32738 3352
rect 32953 3349 32965 3352
rect 32999 3349 33011 3383
rect 32953 3343 33011 3349
rect 34057 3383 34115 3389
rect 34057 3349 34069 3383
rect 34103 3380 34115 3383
rect 34330 3380 34336 3392
rect 34103 3352 34336 3380
rect 34103 3349 34115 3352
rect 34057 3343 34115 3349
rect 34330 3340 34336 3352
rect 34388 3340 34394 3392
rect 34422 3340 34428 3392
rect 34480 3380 34486 3392
rect 38562 3380 38568 3392
rect 34480 3352 38568 3380
rect 34480 3340 34486 3352
rect 38562 3340 38568 3352
rect 38620 3340 38626 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 3384 3148 3433 3176
rect 3384 3136 3390 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 4522 3176 4528 3188
rect 3421 3139 3479 3145
rect 3988 3148 4528 3176
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 3988 3108 4016 3148
rect 4522 3136 4528 3148
rect 4580 3176 4586 3188
rect 5534 3176 5540 3188
rect 4580 3148 5540 3176
rect 4580 3136 4586 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 8202 3176 8208 3188
rect 5859 3148 8208 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 9548 3148 9597 3176
rect 9548 3136 9554 3148
rect 9585 3145 9597 3148
rect 9631 3145 9643 3179
rect 9585 3139 9643 3145
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 13688 3148 13737 3176
rect 13688 3136 13694 3148
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 13725 3139 13783 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15930 3176 15936 3188
rect 15891 3148 15936 3176
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 18598 3176 18604 3188
rect 17736 3148 18092 3176
rect 18559 3148 18604 3176
rect 17736 3136 17742 3148
rect 4154 3108 4160 3120
rect 3099 3080 4016 3108
rect 4115 3080 4160 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4890 3108 4896 3120
rect 4851 3080 4896 3108
rect 4890 3068 4896 3080
rect 4948 3068 4954 3120
rect 5074 3068 5080 3120
rect 5132 3108 5138 3120
rect 11422 3108 11428 3120
rect 5132 3080 11428 3108
rect 5132 3068 5138 3080
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 12406 3080 13216 3108
rect 1118 3000 1124 3052
rect 1176 3040 1182 3052
rect 1394 3040 1400 3052
rect 1176 3012 1400 3040
rect 1176 3000 1182 3012
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3694 3040 3700 3052
rect 3384 3012 3700 3040
rect 3384 3000 3390 3012
rect 3694 3000 3700 3012
rect 3752 3040 3758 3052
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3752 3012 3985 3040
rect 3752 3000 3758 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 4706 3040 4712 3052
rect 4619 3012 4712 3040
rect 3973 3003 4031 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 5810 3040 5816 3052
rect 5675 3012 5816 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6546 3040 6552 3052
rect 6288 3012 6552 3040
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 1673 2935 1731 2941
rect 1688 2904 1716 2935
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 4724 2972 4752 3000
rect 6288 2972 6316 3012
rect 6546 3000 6552 3012
rect 6604 3040 6610 3052
rect 6789 3043 6847 3049
rect 6789 3040 6801 3043
rect 6604 3012 6801 3040
rect 6604 3000 6610 3012
rect 6789 3009 6801 3012
rect 6835 3009 6847 3043
rect 6789 3003 6847 3009
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 8076 3012 8125 3040
rect 8076 3000 8082 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 9401 3043 9459 3049
rect 8113 3003 8171 3009
rect 8312 3012 9352 3040
rect 3936 2944 4752 2972
rect 5552 2944 6316 2972
rect 7009 2975 7067 2981
rect 3936 2932 3942 2944
rect 4430 2904 4436 2916
rect 1688 2876 4436 2904
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 5442 2904 5448 2916
rect 4764 2876 5448 2904
rect 4764 2864 4770 2876
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 5552 2848 5580 2944
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 8312 2972 8340 3012
rect 7055 2944 8340 2972
rect 8389 2975 8447 2981
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 9214 2972 9220 2984
rect 8435 2944 9220 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9324 2972 9352 3012
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 10134 3040 10140 3052
rect 9447 3012 10140 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 10134 3000 10140 3012
rect 10192 3040 10198 3052
rect 10594 3040 10600 3052
rect 10192 3012 10600 3040
rect 10192 3000 10198 3012
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 11606 3040 11612 3052
rect 11563 3012 11612 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 11848 3012 12265 3040
rect 11848 3000 11854 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 9858 2972 9864 2984
rect 9324 2944 9864 2972
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 10008 2944 10057 2972
rect 10008 2932 10014 2944
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 12406 2972 12434 3080
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12676 3012 13001 3040
rect 12676 3000 12682 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 13188 3040 13216 3080
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 15746 3108 15752 3120
rect 13320 3080 15752 3108
rect 13320 3068 13326 3080
rect 15746 3068 15752 3080
rect 15804 3108 15810 3120
rect 17954 3108 17960 3120
rect 15804 3080 16160 3108
rect 17915 3080 17960 3108
rect 15804 3068 15810 3080
rect 13906 3040 13912 3052
rect 13188 3012 13768 3040
rect 13867 3012 13912 3040
rect 12989 3003 13047 3009
rect 10367 2944 12434 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 10778 2904 10784 2916
rect 5684 2876 10784 2904
rect 5684 2864 5690 2876
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 13173 2907 13231 2913
rect 13173 2904 13185 2907
rect 11388 2876 13185 2904
rect 11388 2864 11394 2876
rect 13173 2873 13185 2876
rect 13219 2873 13231 2907
rect 13740 2904 13768 3012
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14366 3040 14372 3052
rect 14279 3012 14372 3040
rect 14366 3000 14372 3012
rect 14424 3040 14430 3052
rect 14642 3040 14648 3052
rect 14424 3012 14648 3040
rect 14424 3000 14430 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15102 3000 15108 3052
rect 15160 3040 15166 3052
rect 16132 3049 16160 3080
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18064 3108 18092 3148
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 20036 3148 20085 3176
rect 20036 3136 20042 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 24026 3176 24032 3188
rect 20073 3139 20131 3145
rect 22066 3148 24032 3176
rect 22066 3108 22094 3148
rect 24026 3136 24032 3148
rect 24084 3136 24090 3188
rect 24857 3179 24915 3185
rect 24857 3145 24869 3179
rect 24903 3176 24915 3179
rect 35158 3176 35164 3188
rect 24903 3148 35164 3176
rect 24903 3145 24915 3148
rect 24857 3139 24915 3145
rect 35158 3136 35164 3148
rect 35216 3136 35222 3188
rect 36354 3136 36360 3188
rect 36412 3176 36418 3188
rect 36633 3179 36691 3185
rect 36633 3176 36645 3179
rect 36412 3148 36645 3176
rect 36412 3136 36418 3148
rect 36633 3145 36645 3148
rect 36679 3145 36691 3179
rect 36633 3139 36691 3145
rect 28166 3108 28172 3120
rect 18064 3080 22094 3108
rect 22940 3080 28172 3108
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 15160 3012 15209 3040
rect 15160 3000 15166 3012
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 17218 3040 17224 3052
rect 16715 3012 17224 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16684 2972 16712 3003
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 17736 3012 17785 3040
rect 17736 3000 17742 3012
rect 17773 3009 17785 3012
rect 17819 3040 17831 3043
rect 18046 3040 18052 3052
rect 17819 3012 18052 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 18380 3012 18429 3040
rect 18380 3000 18386 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 18417 3003 18475 3009
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3040 19947 3043
rect 20162 3040 20168 3052
rect 19935 3012 20168 3040
rect 19935 3009 19947 3012
rect 19889 3003 19947 3009
rect 15988 2944 16712 2972
rect 15988 2932 15994 2944
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 18340 2972 18368 3000
rect 16816 2944 18368 2972
rect 16816 2932 16822 2944
rect 18966 2932 18972 2984
rect 19024 2972 19030 2984
rect 19904 2972 19932 3003
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 20990 3040 20996 3052
rect 20951 3012 20996 3040
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 22094 3040 22100 3052
rect 22055 3012 22100 3040
rect 22094 3000 22100 3012
rect 22152 3000 22158 3052
rect 22940 3049 22968 3080
rect 28166 3068 28172 3080
rect 28224 3068 28230 3120
rect 28350 3108 28356 3120
rect 28311 3080 28356 3108
rect 28350 3068 28356 3080
rect 28408 3068 28414 3120
rect 28810 3108 28816 3120
rect 28771 3080 28816 3108
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 28902 3068 28908 3120
rect 28960 3108 28966 3120
rect 29549 3111 29607 3117
rect 29549 3108 29561 3111
rect 28960 3080 29561 3108
rect 28960 3068 28966 3080
rect 29549 3077 29561 3080
rect 29595 3077 29607 3111
rect 34422 3108 34428 3120
rect 29549 3071 29607 3077
rect 31036 3080 34428 3108
rect 22925 3043 22983 3049
rect 22925 3009 22937 3043
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 23750 3040 23756 3052
rect 23164 3012 23756 3040
rect 23164 3000 23170 3012
rect 23750 3000 23756 3012
rect 23808 3040 23814 3052
rect 24029 3043 24087 3049
rect 24029 3040 24041 3043
rect 23808 3012 24041 3040
rect 23808 3000 23814 3012
rect 24029 3009 24041 3012
rect 24075 3009 24087 3043
rect 24486 3040 24492 3052
rect 24029 3003 24087 3009
rect 24136 3012 24492 3040
rect 19024 2944 19932 2972
rect 19024 2932 19030 2944
rect 19978 2932 19984 2984
rect 20036 2972 20042 2984
rect 20346 2972 20352 2984
rect 20036 2944 20352 2972
rect 20036 2932 20042 2944
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 22612 2944 22661 2972
rect 22612 2932 22618 2944
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 23382 2932 23388 2984
rect 23440 2972 23446 2984
rect 24136 2972 24164 3012
rect 24486 3000 24492 3012
rect 24544 3040 24550 3052
rect 24765 3043 24823 3049
rect 24765 3040 24777 3043
rect 24544 3012 24777 3040
rect 24544 3000 24550 3012
rect 24765 3009 24777 3012
rect 24811 3009 24823 3043
rect 25406 3040 25412 3052
rect 25367 3012 25412 3040
rect 24765 3003 24823 3009
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 26145 3043 26203 3049
rect 26145 3040 26157 3043
rect 25924 3012 26157 3040
rect 25924 3000 25930 3012
rect 26145 3009 26157 3012
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 27430 3000 27436 3052
rect 27488 3040 27494 3052
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 27488 3012 27721 3040
rect 27488 3000 27494 3012
rect 27709 3009 27721 3012
rect 27755 3040 27767 3043
rect 27982 3040 27988 3052
rect 27755 3012 27988 3040
rect 27755 3009 27767 3012
rect 27709 3003 27767 3009
rect 27982 3000 27988 3012
rect 28040 3000 28046 3052
rect 28074 3000 28080 3052
rect 28132 3040 28138 3052
rect 28997 3043 29055 3049
rect 28997 3040 29009 3043
rect 28132 3012 29009 3040
rect 28132 3000 28138 3012
rect 28997 3009 29009 3012
rect 29043 3009 29055 3043
rect 28997 3003 29055 3009
rect 29733 3043 29791 3049
rect 29733 3009 29745 3043
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 23440 2944 24164 2972
rect 24213 2975 24271 2981
rect 23440 2932 23446 2944
rect 24213 2941 24225 2975
rect 24259 2972 24271 2975
rect 24259 2944 28856 2972
rect 24259 2941 24271 2944
rect 24213 2935 24271 2941
rect 18230 2904 18236 2916
rect 13740 2876 18236 2904
rect 13173 2867 13231 2873
rect 18230 2864 18236 2876
rect 18288 2864 18294 2916
rect 24486 2864 24492 2916
rect 24544 2904 24550 2916
rect 25593 2907 25651 2913
rect 25593 2904 25605 2907
rect 24544 2876 25605 2904
rect 24544 2864 24550 2876
rect 25593 2873 25605 2876
rect 25639 2873 25651 2907
rect 26329 2907 26387 2913
rect 26329 2904 26341 2907
rect 25593 2867 25651 2873
rect 25700 2876 26341 2904
rect 106 2796 112 2848
rect 164 2836 170 2848
rect 1394 2836 1400 2848
rect 164 2808 1400 2836
rect 164 2796 170 2808
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 5534 2796 5540 2848
rect 5592 2796 5598 2848
rect 7558 2836 7564 2848
rect 7519 2808 7564 2836
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 8904 2808 11713 2836
rect 8904 2796 8910 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 11701 2799 11759 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12492 2808 12537 2836
rect 12492 2796 12498 2808
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 19245 2839 19303 2845
rect 19245 2836 19257 2839
rect 18748 2808 19257 2836
rect 18748 2796 18754 2808
rect 19245 2805 19257 2808
rect 19291 2805 19303 2839
rect 19245 2799 19303 2805
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20404 2808 20821 2836
rect 20404 2796 20410 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 21913 2839 21971 2845
rect 21913 2836 21925 2839
rect 21232 2808 21925 2836
rect 21232 2796 21238 2808
rect 21913 2805 21925 2808
rect 21959 2805 21971 2839
rect 21913 2799 21971 2805
rect 25314 2796 25320 2848
rect 25372 2836 25378 2848
rect 25700 2836 25728 2876
rect 26329 2873 26341 2876
rect 26375 2873 26387 2907
rect 26329 2867 26387 2873
rect 26418 2864 26424 2916
rect 26476 2904 26482 2916
rect 27522 2904 27528 2916
rect 26476 2876 27384 2904
rect 27483 2876 27528 2904
rect 26476 2864 26482 2876
rect 25372 2808 25728 2836
rect 25372 2796 25378 2808
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 25832 2808 26985 2836
rect 25832 2796 25838 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 27356 2836 27384 2876
rect 27522 2864 27528 2876
rect 27580 2864 27586 2916
rect 28828 2904 28856 2944
rect 28902 2932 28908 2984
rect 28960 2972 28966 2984
rect 29086 2972 29092 2984
rect 28960 2944 29092 2972
rect 28960 2932 28966 2944
rect 29086 2932 29092 2944
rect 29144 2972 29150 2984
rect 29748 2972 29776 3003
rect 30466 3000 30472 3052
rect 30524 3040 30530 3052
rect 30561 3043 30619 3049
rect 30561 3040 30573 3043
rect 30524 3012 30573 3040
rect 30524 3000 30530 3012
rect 30561 3009 30573 3012
rect 30607 3009 30619 3043
rect 30834 3040 30840 3052
rect 30795 3012 30840 3040
rect 30561 3003 30619 3009
rect 30834 3000 30840 3012
rect 30892 3000 30898 3052
rect 29144 2944 29776 2972
rect 29144 2932 29150 2944
rect 31036 2904 31064 3080
rect 34422 3068 34428 3080
rect 34480 3068 34486 3120
rect 34882 3108 34888 3120
rect 34843 3080 34888 3108
rect 34882 3068 34888 3080
rect 34940 3068 34946 3120
rect 35434 3068 35440 3120
rect 35492 3108 35498 3120
rect 35710 3108 35716 3120
rect 35492 3080 35716 3108
rect 35492 3068 35498 3080
rect 35710 3068 35716 3080
rect 35768 3068 35774 3120
rect 38286 3108 38292 3120
rect 36280 3080 38292 3108
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 32493 3043 32551 3049
rect 32493 3040 32505 3043
rect 32456 3012 32505 3040
rect 32456 3000 32462 3012
rect 32493 3009 32505 3012
rect 32539 3040 32551 3043
rect 32582 3040 32588 3052
rect 32539 3012 32588 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 32582 3000 32588 3012
rect 32640 3000 32646 3052
rect 33778 3040 33784 3052
rect 33739 3012 33784 3040
rect 33778 3000 33784 3012
rect 33836 3000 33842 3052
rect 32122 2932 32128 2984
rect 32180 2972 32186 2984
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 32180 2944 32781 2972
rect 32180 2932 32186 2944
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 34900 2972 34928 3068
rect 35069 3043 35127 3049
rect 35069 3009 35081 3043
rect 35115 3040 35127 3043
rect 36280 3040 36308 3080
rect 38286 3068 38292 3080
rect 38344 3068 38350 3120
rect 36446 3040 36452 3052
rect 35115 3012 36308 3040
rect 36407 3012 36452 3040
rect 35115 3009 35127 3012
rect 35069 3003 35127 3009
rect 36446 3000 36452 3012
rect 36504 3000 36510 3052
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 37458 3040 37464 3052
rect 37323 3012 37464 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 37458 3000 37464 3012
rect 37516 3000 37522 3052
rect 34900 2944 37320 2972
rect 32769 2935 32827 2941
rect 35529 2907 35587 2913
rect 35529 2904 35541 2907
rect 28828 2876 31064 2904
rect 31726 2876 35541 2904
rect 31726 2836 31754 2876
rect 35529 2873 35541 2876
rect 35575 2873 35587 2907
rect 37292 2904 37320 2944
rect 37366 2932 37372 2984
rect 37424 2972 37430 2984
rect 37553 2975 37611 2981
rect 37553 2972 37565 2975
rect 37424 2944 37565 2972
rect 37424 2932 37430 2944
rect 37553 2941 37565 2944
rect 37599 2941 37611 2975
rect 37553 2935 37611 2941
rect 38746 2904 38752 2916
rect 37292 2876 38752 2904
rect 35529 2867 35587 2873
rect 38746 2864 38752 2876
rect 38804 2864 38810 2916
rect 27356 2808 31754 2836
rect 26973 2799 27031 2805
rect 33502 2796 33508 2848
rect 33560 2836 33566 2848
rect 33965 2839 34023 2845
rect 33965 2836 33977 2839
rect 33560 2808 33977 2836
rect 33560 2796 33566 2808
rect 33965 2805 33977 2808
rect 34011 2805 34023 2839
rect 33965 2799 34023 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 6595 2635 6653 2641
rect 6595 2601 6607 2635
rect 6641 2632 6653 2635
rect 6641 2604 6914 2632
rect 6641 2601 6653 2604
rect 6595 2595 6653 2601
rect 6886 2564 6914 2604
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 9732 2604 12817 2632
rect 9732 2592 9738 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 15933 2635 15991 2641
rect 15933 2601 15945 2635
rect 15979 2632 15991 2635
rect 21910 2632 21916 2644
rect 15979 2604 20116 2632
rect 21871 2604 21916 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 10042 2564 10048 2576
rect 6886 2536 10048 2564
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 14918 2564 14924 2576
rect 10152 2536 14924 2564
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 3050 2496 3056 2508
rect 1719 2468 3056 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 4488 2468 4537 2496
rect 4488 2456 4494 2468
rect 4525 2465 4537 2468
rect 4571 2496 4583 2499
rect 4614 2496 4620 2508
rect 4571 2468 4620 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 9030 2496 9036 2508
rect 4847 2468 9036 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 9217 2499 9275 2505
rect 9217 2496 9229 2499
rect 9180 2468 9229 2496
rect 9180 2456 9186 2468
rect 9217 2465 9229 2468
rect 9263 2496 9275 2499
rect 9582 2496 9588 2508
rect 9263 2468 9588 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2590 2428 2596 2440
rect 2280 2400 2596 2428
rect 2280 2388 2286 2400
rect 2590 2388 2596 2400
rect 2648 2428 2654 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2648 2400 2789 2428
rect 2648 2388 2654 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 2924 2400 3893 2428
rect 2924 2388 2930 2400
rect 3881 2397 3893 2400
rect 3927 2428 3939 2431
rect 4062 2428 4068 2440
rect 3927 2400 4068 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5040 2400 6377 2428
rect 5040 2388 5046 2400
rect 6365 2397 6377 2400
rect 6411 2428 6423 2431
rect 6454 2428 6460 2440
rect 6411 2400 6460 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 6886 2400 7757 2428
rect 1394 2320 1400 2372
rect 1452 2360 1458 2372
rect 1762 2360 1768 2372
rect 1452 2332 1768 2360
rect 1452 2320 1458 2332
rect 1762 2320 1768 2332
rect 1820 2320 1826 2372
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4798 2360 4804 2372
rect 4212 2332 4804 2360
rect 4212 2320 4218 2332
rect 4798 2320 4804 2332
rect 4856 2320 4862 2372
rect 6086 2320 6092 2372
rect 6144 2360 6150 2372
rect 6886 2360 6914 2400
rect 7745 2397 7757 2400
rect 7791 2428 7803 2431
rect 8110 2428 8116 2440
rect 7791 2400 8116 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 10152 2428 10180 2536
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 18509 2567 18567 2573
rect 18509 2533 18521 2567
rect 18555 2564 18567 2567
rect 18782 2564 18788 2576
rect 18555 2536 18788 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 18782 2524 18788 2536
rect 18840 2524 18846 2576
rect 20088 2564 20116 2604
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 23566 2632 23572 2644
rect 22020 2604 23572 2632
rect 22020 2564 22048 2604
rect 23566 2592 23572 2604
rect 23624 2592 23630 2644
rect 23842 2632 23848 2644
rect 23803 2604 23848 2632
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 31386 2632 31392 2644
rect 24412 2604 31392 2632
rect 20088 2536 22048 2564
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10376 2468 12664 2496
rect 10376 2456 10382 2468
rect 9539 2400 10180 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10284 2400 10609 2428
rect 10284 2388 10290 2400
rect 10597 2397 10609 2400
rect 10643 2428 10655 2431
rect 10686 2428 10692 2440
rect 10643 2400 10692 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 12636 2437 12664 2468
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 24412 2496 24440 2604
rect 31386 2592 31392 2604
rect 31444 2592 31450 2644
rect 31726 2604 34100 2632
rect 25774 2524 25780 2576
rect 25832 2564 25838 2576
rect 31726 2564 31754 2604
rect 25832 2536 31754 2564
rect 34072 2564 34100 2604
rect 34698 2592 34704 2644
rect 34756 2632 34762 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34756 2604 34897 2632
rect 34756 2592 34762 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 36446 2564 36452 2576
rect 34072 2536 36452 2564
rect 25832 2524 25838 2536
rect 36446 2524 36452 2536
rect 36504 2524 36510 2576
rect 14516 2468 24440 2496
rect 24673 2499 24731 2505
rect 14516 2456 14522 2468
rect 24673 2465 24685 2499
rect 24719 2496 24731 2499
rect 30009 2499 30067 2505
rect 24719 2468 29868 2496
rect 24719 2465 24731 2468
rect 24673 2459 24731 2465
rect 12621 2431 12679 2437
rect 10836 2400 10881 2428
rect 10836 2388 10842 2400
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 12621 2391 12679 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15712 2400 15761 2428
rect 15712 2388 15718 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 16482 2388 16488 2440
rect 16540 2428 16546 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16540 2400 16681 2428
rect 16540 2388 16546 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17310 2388 17316 2440
rect 17368 2428 17374 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17368 2400 17509 2428
rect 17368 2388 17374 2400
rect 17497 2397 17509 2400
rect 17543 2428 17555 2431
rect 17586 2428 17592 2440
rect 17543 2400 17592 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 20349 2431 20407 2437
rect 20349 2428 20361 2431
rect 20312 2400 20361 2428
rect 20312 2388 20318 2400
rect 20349 2397 20361 2400
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22336 2400 22385 2428
rect 22336 2388 22342 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 23661 2431 23719 2437
rect 23661 2397 23673 2431
rect 23707 2397 23719 2431
rect 24394 2428 24400 2440
rect 24355 2400 24400 2428
rect 23661 2391 23719 2397
rect 6144 2332 6914 2360
rect 6144 2320 6150 2332
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 11238 2360 11244 2372
rect 8352 2332 11244 2360
rect 8352 2320 8358 2332
rect 11238 2320 11244 2332
rect 11296 2360 11302 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11296 2332 11989 2360
rect 11296 2320 11302 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 12161 2363 12219 2369
rect 12161 2329 12173 2363
rect 12207 2360 12219 2363
rect 12526 2360 12532 2372
rect 12207 2332 12532 2360
rect 12207 2329 12219 2332
rect 12161 2323 12219 2329
rect 12526 2320 12532 2332
rect 12584 2320 12590 2372
rect 13814 2360 13820 2372
rect 12728 2332 13820 2360
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 7837 2295 7895 2301
rect 7837 2261 7849 2295
rect 7883 2292 7895 2295
rect 12728 2292 12756 2332
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 18138 2320 18144 2372
rect 18196 2360 18202 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 18196 2332 18337 2360
rect 18196 2320 18202 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 18325 2323 18383 2329
rect 18414 2320 18420 2372
rect 18472 2360 18478 2372
rect 19150 2360 19156 2372
rect 18472 2332 19156 2360
rect 18472 2320 18478 2332
rect 19150 2320 19156 2332
rect 19208 2360 19214 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19208 2332 19717 2360
rect 19208 2320 19214 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 19889 2363 19947 2369
rect 19889 2329 19901 2363
rect 19935 2360 19947 2363
rect 20622 2360 20628 2372
rect 19935 2332 20628 2360
rect 19935 2329 19947 2332
rect 19889 2323 19947 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 23676 2360 23704 2391
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 27246 2388 27252 2440
rect 27304 2428 27310 2440
rect 27525 2431 27583 2437
rect 27525 2428 27537 2431
rect 27304 2400 27537 2428
rect 27304 2388 27310 2400
rect 27525 2397 27537 2400
rect 27571 2397 27583 2431
rect 28074 2428 28080 2440
rect 28035 2400 28080 2428
rect 27525 2391 27583 2397
rect 28074 2388 28080 2400
rect 28132 2388 28138 2440
rect 28994 2428 29000 2440
rect 28955 2400 29000 2428
rect 28994 2388 29000 2400
rect 29052 2388 29058 2440
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29840 2428 29868 2468
rect 30009 2465 30021 2499
rect 30055 2496 30067 2499
rect 30098 2496 30104 2508
rect 30055 2468 30104 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 30098 2456 30104 2468
rect 30156 2456 30162 2508
rect 32214 2496 32220 2508
rect 32175 2468 32220 2496
rect 32214 2456 32220 2468
rect 32272 2456 32278 2508
rect 32490 2496 32496 2508
rect 32451 2468 32496 2496
rect 32490 2456 32496 2468
rect 32548 2456 32554 2508
rect 35897 2499 35955 2505
rect 35897 2465 35909 2499
rect 35943 2496 35955 2499
rect 36078 2496 36084 2508
rect 35943 2468 36084 2496
rect 35943 2465 35955 2468
rect 35897 2459 35955 2465
rect 36078 2456 36084 2468
rect 36136 2496 36142 2508
rect 36538 2496 36544 2508
rect 36136 2468 36544 2496
rect 36136 2456 36142 2468
rect 36538 2456 36544 2468
rect 36596 2456 36602 2508
rect 37550 2496 37556 2508
rect 37511 2468 37556 2496
rect 37550 2456 37556 2468
rect 37608 2456 37614 2508
rect 34057 2431 34115 2437
rect 29840 2400 34008 2428
rect 29733 2391 29791 2397
rect 24762 2360 24768 2372
rect 21315 2332 24768 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 26145 2363 26203 2369
rect 26145 2360 26157 2363
rect 24912 2332 26157 2360
rect 24912 2320 24918 2332
rect 26145 2329 26157 2332
rect 26191 2329 26203 2363
rect 26145 2323 26203 2329
rect 26329 2363 26387 2369
rect 26329 2329 26341 2363
rect 26375 2360 26387 2363
rect 26694 2360 26700 2372
rect 26375 2332 26700 2360
rect 26375 2329 26387 2332
rect 26329 2323 26387 2329
rect 26694 2320 26700 2332
rect 26752 2320 26758 2372
rect 27338 2360 27344 2372
rect 27299 2332 27344 2360
rect 27338 2320 27344 2332
rect 27396 2320 27402 2372
rect 28261 2363 28319 2369
rect 28261 2329 28273 2363
rect 28307 2329 28319 2363
rect 28261 2323 28319 2329
rect 7883 2264 12756 2292
rect 7883 2261 7895 2264
rect 7837 2255 7895 2261
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 13449 2295 13507 2301
rect 13449 2292 13461 2295
rect 12860 2264 13461 2292
rect 12860 2252 12866 2264
rect 13449 2261 13461 2264
rect 13495 2292 13507 2295
rect 13538 2292 13544 2304
rect 13495 2264 13544 2292
rect 13495 2261 13507 2264
rect 13449 2255 13507 2261
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 14274 2292 14280 2304
rect 14235 2264 14280 2292
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 15068 2264 15117 2292
rect 15068 2252 15074 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 16850 2292 16856 2304
rect 16811 2264 16856 2292
rect 15105 2255 15163 2261
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 17589 2295 17647 2301
rect 17589 2261 17601 2295
rect 17635 2292 17647 2295
rect 19334 2292 19340 2304
rect 17635 2264 19340 2292
rect 17635 2261 17647 2264
rect 17589 2255 17647 2261
rect 19334 2252 19340 2264
rect 19392 2252 19398 2304
rect 19426 2252 19432 2304
rect 19484 2292 19490 2304
rect 20533 2295 20591 2301
rect 20533 2292 20545 2295
rect 19484 2264 20545 2292
rect 19484 2252 19490 2264
rect 20533 2261 20545 2264
rect 20579 2261 20591 2295
rect 20533 2255 20591 2261
rect 22603 2295 22661 2301
rect 22603 2261 22615 2295
rect 22649 2292 22661 2295
rect 25774 2292 25780 2304
rect 22649 2264 25780 2292
rect 22649 2261 22661 2264
rect 22603 2255 22661 2261
rect 25774 2252 25780 2264
rect 25832 2252 25838 2304
rect 27154 2252 27160 2304
rect 27212 2292 27218 2304
rect 28276 2292 28304 2323
rect 30006 2320 30012 2372
rect 30064 2360 30070 2372
rect 31205 2363 31263 2369
rect 31205 2360 31217 2363
rect 30064 2332 31217 2360
rect 30064 2320 30070 2332
rect 31205 2329 31217 2332
rect 31251 2329 31263 2363
rect 31205 2323 31263 2329
rect 31386 2320 31392 2372
rect 31444 2360 31450 2372
rect 33873 2363 33931 2369
rect 33873 2360 33885 2363
rect 31444 2332 33885 2360
rect 31444 2320 31450 2332
rect 33873 2329 33885 2332
rect 33919 2329 33931 2363
rect 33873 2323 33931 2329
rect 27212 2264 28304 2292
rect 27212 2252 27218 2264
rect 28718 2252 28724 2304
rect 28776 2292 28782 2304
rect 28813 2295 28871 2301
rect 28813 2292 28825 2295
rect 28776 2264 28825 2292
rect 28776 2252 28782 2264
rect 28813 2261 28825 2264
rect 28859 2261 28871 2295
rect 31110 2292 31116 2304
rect 31071 2264 31116 2292
rect 28813 2255 28871 2261
rect 31110 2252 31116 2264
rect 31168 2252 31174 2304
rect 33980 2292 34008 2400
rect 34057 2397 34069 2431
rect 34103 2428 34115 2431
rect 34238 2428 34244 2440
rect 34103 2400 34244 2428
rect 34103 2397 34115 2400
rect 34057 2391 34115 2397
rect 34238 2388 34244 2400
rect 34296 2388 34302 2440
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34664 2400 34713 2428
rect 34664 2388 34670 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 36170 2428 36176 2440
rect 36131 2400 36176 2428
rect 34701 2391 34759 2397
rect 36170 2388 36176 2400
rect 36228 2388 36234 2440
rect 37277 2431 37335 2437
rect 37277 2397 37289 2431
rect 37323 2428 37335 2431
rect 37826 2428 37832 2440
rect 37323 2400 37832 2428
rect 37323 2397 37335 2400
rect 37277 2391 37335 2397
rect 37826 2388 37832 2400
rect 37884 2388 37890 2440
rect 34256 2360 34284 2388
rect 35710 2360 35716 2372
rect 34256 2332 35716 2360
rect 35710 2320 35716 2332
rect 35768 2320 35774 2372
rect 36722 2292 36728 2304
rect 33980 2264 36728 2292
rect 36722 2252 36728 2264
rect 36780 2252 36786 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 7558 2048 7564 2100
rect 7616 2088 7622 2100
rect 31110 2088 31116 2100
rect 7616 2060 31116 2088
rect 7616 2048 7622 2060
rect 31110 2048 31116 2060
rect 31168 2048 31174 2100
rect 2866 1980 2872 2032
rect 2924 2020 2930 2032
rect 12342 2020 12348 2032
rect 2924 1992 12348 2020
rect 2924 1980 2930 1992
rect 12342 1980 12348 1992
rect 12400 1980 12406 2032
rect 13538 1980 13544 2032
rect 13596 2020 13602 2032
rect 13596 1992 31754 2020
rect 13596 1980 13602 1992
rect 3970 1912 3976 1964
rect 4028 1952 4034 1964
rect 14182 1952 14188 1964
rect 4028 1924 14188 1952
rect 4028 1912 4034 1924
rect 14182 1912 14188 1924
rect 14240 1912 14246 1964
rect 22094 1912 22100 1964
rect 22152 1952 22158 1964
rect 28718 1952 28724 1964
rect 22152 1924 28724 1952
rect 22152 1912 22158 1924
rect 28718 1912 28724 1924
rect 28776 1912 28782 1964
rect 12526 1844 12532 1896
rect 12584 1884 12590 1896
rect 23014 1884 23020 1896
rect 12584 1856 23020 1884
rect 12584 1844 12590 1856
rect 23014 1844 23020 1856
rect 23072 1844 23078 1896
rect 26602 1884 26608 1896
rect 23860 1856 26608 1884
rect 12434 1776 12440 1828
rect 12492 1816 12498 1828
rect 13906 1816 13912 1828
rect 12492 1788 13912 1816
rect 12492 1776 12498 1788
rect 13906 1776 13912 1788
rect 13964 1776 13970 1828
rect 16850 1776 16856 1828
rect 16908 1816 16914 1828
rect 23860 1816 23888 1856
rect 26602 1844 26608 1856
rect 26660 1844 26666 1896
rect 31726 1884 31754 1992
rect 34514 1884 34520 1896
rect 31726 1856 34520 1884
rect 34514 1844 34520 1856
rect 34572 1844 34578 1896
rect 16908 1788 23888 1816
rect 16908 1776 16914 1788
rect 23934 1776 23940 1828
rect 23992 1816 23998 1828
rect 24394 1816 24400 1828
rect 23992 1788 24400 1816
rect 23992 1776 23998 1788
rect 24394 1776 24400 1788
rect 24452 1776 24458 1828
rect 16114 1708 16120 1760
rect 16172 1748 16178 1760
rect 36170 1748 36176 1760
rect 16172 1720 36176 1748
rect 16172 1708 16178 1720
rect 36170 1708 36176 1720
rect 36228 1708 36234 1760
rect 19334 1640 19340 1692
rect 19392 1680 19398 1692
rect 19392 1652 22094 1680
rect 19392 1640 19398 1652
rect 22066 1612 22094 1652
rect 26418 1640 26424 1692
rect 26476 1680 26482 1692
rect 27246 1680 27252 1692
rect 26476 1652 27252 1680
rect 26476 1640 26482 1652
rect 27246 1640 27252 1652
rect 27304 1640 27310 1692
rect 29086 1640 29092 1692
rect 29144 1680 29150 1692
rect 30006 1680 30012 1692
rect 29144 1652 30012 1680
rect 29144 1640 29150 1652
rect 30006 1640 30012 1652
rect 30064 1640 30070 1692
rect 28442 1612 28448 1624
rect 22066 1584 28448 1612
rect 28442 1572 28448 1584
rect 28500 1572 28506 1624
<< via1 >>
rect 9680 37612 9732 37664
rect 16028 37612 16080 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 4896 37408 4948 37460
rect 9680 37451 9732 37460
rect 9680 37417 9689 37451
rect 9689 37417 9723 37451
rect 9723 37417 9732 37451
rect 9680 37408 9732 37417
rect 14556 37408 14608 37460
rect 16028 37408 16080 37460
rect 29092 37408 29144 37460
rect 7656 37340 7708 37392
rect 28448 37340 28500 37392
rect 3516 37272 3568 37324
rect 5080 37272 5132 37324
rect 14924 37272 14976 37324
rect 16028 37272 16080 37324
rect 17408 37272 17460 37324
rect 18880 37272 18932 37324
rect 22652 37272 22704 37324
rect 1124 37204 1176 37256
rect 1768 37204 1820 37256
rect 2136 37204 2188 37256
rect 2596 37204 2648 37256
rect 3240 37204 3292 37256
rect 4068 37204 4120 37256
rect 5724 37204 5776 37256
rect 6368 37204 6420 37256
rect 7472 37204 7524 37256
rect 8484 37204 8536 37256
rect 9404 37247 9456 37256
rect 9404 37213 9413 37247
rect 9413 37213 9447 37247
rect 9447 37213 9456 37247
rect 9404 37204 9456 37213
rect 10140 37204 10192 37256
rect 10600 37204 10652 37256
rect 12164 37204 12216 37256
rect 13820 37204 13872 37256
rect 14556 37247 14608 37256
rect 14556 37213 14565 37247
rect 14565 37213 14599 37247
rect 14599 37213 14608 37247
rect 14556 37204 14608 37213
rect 14832 37204 14884 37256
rect 15292 37247 15344 37256
rect 15292 37213 15301 37247
rect 15301 37213 15335 37247
rect 15335 37213 15344 37247
rect 15292 37204 15344 37213
rect 17960 37204 18012 37256
rect 19064 37204 19116 37256
rect 19248 37247 19300 37256
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 20076 37204 20128 37256
rect 20904 37247 20956 37256
rect 20904 37213 20913 37247
rect 20913 37213 20947 37247
rect 20947 37213 20956 37247
rect 20904 37204 20956 37213
rect 21088 37204 21140 37256
rect 30656 37315 30708 37324
rect 30656 37281 30665 37315
rect 30665 37281 30699 37315
rect 30699 37281 30708 37315
rect 30656 37272 30708 37281
rect 32312 37272 32364 37324
rect 4160 37136 4212 37188
rect 5264 37136 5316 37188
rect 11612 37136 11664 37188
rect 13728 37136 13780 37188
rect 15844 37136 15896 37188
rect 17500 37136 17552 37188
rect 22192 37136 22244 37188
rect 24308 37204 24360 37256
rect 25320 37204 25372 37256
rect 25504 37204 25556 37256
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 27068 37204 27120 37256
rect 28540 37204 28592 37256
rect 28908 37204 28960 37256
rect 29460 37204 29512 37256
rect 30564 37204 30616 37256
rect 29644 37136 29696 37188
rect 31208 37136 31260 37188
rect 31760 37204 31812 37256
rect 32772 37204 32824 37256
rect 33508 37247 33560 37256
rect 33508 37213 33517 37247
rect 33517 37213 33551 37247
rect 33551 37213 33560 37247
rect 33508 37204 33560 37213
rect 33784 37204 33836 37256
rect 35440 37204 35492 37256
rect 35716 37247 35768 37256
rect 35716 37213 35725 37247
rect 35725 37213 35759 37247
rect 35759 37213 35768 37247
rect 35716 37204 35768 37213
rect 35900 37204 35952 37256
rect 37280 37247 37332 37256
rect 37280 37213 37289 37247
rect 37289 37213 37323 37247
rect 37323 37213 37332 37247
rect 37280 37204 37332 37213
rect 1952 37111 2004 37120
rect 1952 37077 1961 37111
rect 1961 37077 1995 37111
rect 1995 37077 2004 37111
rect 1952 37068 2004 37077
rect 2780 37068 2832 37120
rect 7840 37111 7892 37120
rect 7840 37077 7849 37111
rect 7849 37077 7883 37111
rect 7883 37077 7892 37111
rect 7840 37068 7892 37077
rect 10600 37068 10652 37120
rect 12072 37111 12124 37120
rect 12072 37077 12081 37111
rect 12081 37077 12115 37111
rect 12115 37077 12124 37111
rect 12072 37068 12124 37077
rect 20168 37068 20220 37120
rect 20352 37111 20404 37120
rect 20352 37077 20361 37111
rect 20361 37077 20395 37111
rect 20395 37077 20404 37111
rect 20352 37068 20404 37077
rect 20444 37068 20496 37120
rect 23020 37068 23072 37120
rect 24584 37111 24636 37120
rect 24584 37077 24593 37111
rect 24593 37077 24627 37111
rect 24627 37077 24636 37111
rect 24584 37068 24636 37077
rect 25596 37111 25648 37120
rect 25596 37077 25605 37111
rect 25605 37077 25639 37111
rect 25639 37077 25648 37111
rect 25596 37068 25648 37077
rect 25688 37068 25740 37120
rect 26792 37068 26844 37120
rect 27804 37068 27856 37120
rect 28724 37111 28776 37120
rect 28724 37077 28733 37111
rect 28733 37077 28767 37111
rect 28767 37077 28776 37111
rect 28724 37068 28776 37077
rect 29736 37111 29788 37120
rect 29736 37077 29745 37111
rect 29745 37077 29779 37111
rect 29779 37077 29788 37111
rect 29736 37068 29788 37077
rect 31392 37111 31444 37120
rect 31392 37077 31401 37111
rect 31401 37077 31435 37111
rect 31435 37077 31444 37111
rect 31392 37068 31444 37077
rect 33692 37068 33744 37120
rect 34612 37068 34664 37120
rect 34888 37068 34940 37120
rect 36268 37111 36320 37120
rect 36268 37077 36277 37111
rect 36277 37077 36311 37111
rect 36311 37077 36320 37111
rect 36268 37068 36320 37077
rect 38384 37136 38436 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2504 36864 2556 36916
rect 3608 36864 3660 36916
rect 4620 36864 4672 36916
rect 4988 36864 5040 36916
rect 5816 36864 5868 36916
rect 7748 36864 7800 36916
rect 8852 36864 8904 36916
rect 10968 36864 11020 36916
rect 11980 36864 12032 36916
rect 13084 36864 13136 36916
rect 14096 36864 14148 36916
rect 15200 36864 15252 36916
rect 17224 36864 17276 36916
rect 18328 36864 18380 36916
rect 19340 36864 19392 36916
rect 19984 36864 20036 36916
rect 20812 36864 20864 36916
rect 21456 36864 21508 36916
rect 22560 36864 22612 36916
rect 23572 36864 23624 36916
rect 24860 36864 24912 36916
rect 25044 36864 25096 36916
rect 26240 36864 26292 36916
rect 27344 36864 27396 36916
rect 28172 36864 28224 36916
rect 29184 36864 29236 36916
rect 29920 36864 29972 36916
rect 30932 36864 30984 36916
rect 32036 36864 32088 36916
rect 33140 36864 33192 36916
rect 34152 36864 34204 36916
rect 34796 36864 34848 36916
rect 112 36796 164 36848
rect 1584 36796 1636 36848
rect 7472 36796 7524 36848
rect 12716 36796 12768 36848
rect 13728 36796 13780 36848
rect 16948 36796 17000 36848
rect 22836 36796 22888 36848
rect 31392 36796 31444 36848
rect 34336 36796 34388 36848
rect 34888 36796 34940 36848
rect 35348 36864 35400 36916
rect 36360 36864 36412 36916
rect 35716 36796 35768 36848
rect 38016 36796 38068 36848
rect 2780 36771 2832 36780
rect 2780 36737 2789 36771
rect 2789 36737 2823 36771
rect 2823 36737 2832 36771
rect 2780 36728 2832 36737
rect 3240 36771 3292 36780
rect 3240 36737 3249 36771
rect 3249 36737 3283 36771
rect 3283 36737 3292 36771
rect 3240 36728 3292 36737
rect 4620 36728 4672 36780
rect 5356 36728 5408 36780
rect 5540 36728 5592 36780
rect 5632 36728 5684 36780
rect 6184 36728 6236 36780
rect 7104 36771 7156 36780
rect 7104 36737 7113 36771
rect 7113 36737 7147 36771
rect 7147 36737 7156 36771
rect 7104 36728 7156 36737
rect 7932 36728 7984 36780
rect 8576 36771 8628 36780
rect 8576 36737 8585 36771
rect 8585 36737 8619 36771
rect 8619 36737 8628 36771
rect 8576 36728 8628 36737
rect 9772 36728 9824 36780
rect 10692 36771 10744 36780
rect 10692 36737 10701 36771
rect 10701 36737 10735 36771
rect 10735 36737 10744 36771
rect 10692 36728 10744 36737
rect 13360 36728 13412 36780
rect 14280 36771 14332 36780
rect 9404 36660 9456 36712
rect 14280 36737 14289 36771
rect 14289 36737 14323 36771
rect 14323 36737 14332 36771
rect 14280 36728 14332 36737
rect 16672 36728 16724 36780
rect 18052 36771 18104 36780
rect 18052 36737 18061 36771
rect 18061 36737 18095 36771
rect 18095 36737 18104 36771
rect 18052 36728 18104 36737
rect 19432 36728 19484 36780
rect 20168 36728 20220 36780
rect 20444 36771 20496 36780
rect 20444 36737 20453 36771
rect 20453 36737 20487 36771
rect 20487 36737 20496 36771
rect 20444 36728 20496 36737
rect 20536 36728 20588 36780
rect 20996 36728 21048 36780
rect 22560 36771 22612 36780
rect 22560 36737 22569 36771
rect 22569 36737 22603 36771
rect 22603 36737 22612 36771
rect 22560 36728 22612 36737
rect 23204 36728 23256 36780
rect 23480 36728 23532 36780
rect 23756 36728 23808 36780
rect 14832 36660 14884 36712
rect 15384 36660 15436 36712
rect 25412 36728 25464 36780
rect 26424 36771 26476 36780
rect 26424 36737 26433 36771
rect 26433 36737 26467 36771
rect 26467 36737 26476 36771
rect 26424 36728 26476 36737
rect 26884 36728 26936 36780
rect 27252 36728 27304 36780
rect 28632 36728 28684 36780
rect 28172 36660 28224 36712
rect 29368 36728 29420 36780
rect 31024 36771 31076 36780
rect 31024 36737 31033 36771
rect 31033 36737 31067 36771
rect 31067 36737 31076 36771
rect 31024 36728 31076 36737
rect 31944 36728 31996 36780
rect 33140 36771 33192 36780
rect 33140 36737 33149 36771
rect 33149 36737 33183 36771
rect 33183 36737 33192 36771
rect 33140 36728 33192 36737
rect 34244 36771 34296 36780
rect 34244 36737 34253 36771
rect 34253 36737 34287 36771
rect 34287 36737 34296 36771
rect 34244 36728 34296 36737
rect 34796 36728 34848 36780
rect 36176 36728 36228 36780
rect 2044 36635 2096 36644
rect 2044 36601 2053 36635
rect 2053 36601 2087 36635
rect 2087 36601 2096 36635
rect 2044 36592 2096 36601
rect 6644 36635 6696 36644
rect 6644 36601 6653 36635
rect 6653 36601 6687 36635
rect 6687 36601 6696 36635
rect 6644 36592 6696 36601
rect 6920 36592 6972 36644
rect 13636 36592 13688 36644
rect 18052 36592 18104 36644
rect 18604 36592 18656 36644
rect 37556 36592 37608 36644
rect 38568 36592 38620 36644
rect 1492 36524 1544 36576
rect 6368 36524 6420 36576
rect 6736 36524 6788 36576
rect 17224 36567 17276 36576
rect 17224 36533 17233 36567
rect 17233 36533 17267 36567
rect 17267 36533 17276 36567
rect 17224 36524 17276 36533
rect 23388 36567 23440 36576
rect 23388 36533 23397 36567
rect 23397 36533 23431 36567
rect 23431 36533 23440 36567
rect 23388 36524 23440 36533
rect 26240 36567 26292 36576
rect 26240 36533 26249 36567
rect 26249 36533 26283 36567
rect 26283 36533 26292 36567
rect 26240 36524 26292 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 388 36320 440 36372
rect 1860 36320 1912 36372
rect 2872 36320 2924 36372
rect 3884 36320 3936 36372
rect 5356 36363 5408 36372
rect 5356 36329 5365 36363
rect 5365 36329 5399 36363
rect 5399 36329 5408 36363
rect 5356 36320 5408 36329
rect 6000 36320 6052 36372
rect 7196 36320 7248 36372
rect 7932 36363 7984 36372
rect 7932 36329 7941 36363
rect 7941 36329 7975 36363
rect 7975 36329 7984 36363
rect 7932 36320 7984 36329
rect 8300 36320 8352 36372
rect 9864 36320 9916 36372
rect 10232 36320 10284 36372
rect 11336 36320 11388 36372
rect 12440 36320 12492 36372
rect 13452 36320 13504 36372
rect 14464 36320 14516 36372
rect 16212 36320 16264 36372
rect 16580 36320 16632 36372
rect 17592 36320 17644 36372
rect 19340 36363 19392 36372
rect 19340 36329 19349 36363
rect 19349 36329 19383 36363
rect 19383 36329 19392 36363
rect 19340 36320 19392 36329
rect 20536 36320 20588 36372
rect 20996 36320 21048 36372
rect 21824 36320 21876 36372
rect 23756 36320 23808 36372
rect 23940 36320 23992 36372
rect 25320 36363 25372 36372
rect 25320 36329 25329 36363
rect 25329 36329 25363 36363
rect 25363 36329 25372 36363
rect 25320 36320 25372 36329
rect 26424 36320 26476 36372
rect 27068 36320 27120 36372
rect 27252 36363 27304 36372
rect 27252 36329 27261 36363
rect 27261 36329 27295 36363
rect 27295 36329 27304 36363
rect 27252 36320 27304 36329
rect 28172 36363 28224 36372
rect 28172 36329 28181 36363
rect 28181 36329 28215 36363
rect 28215 36329 28224 36363
rect 28172 36320 28224 36329
rect 28632 36363 28684 36372
rect 28632 36329 28641 36363
rect 28641 36329 28675 36363
rect 28675 36329 28684 36363
rect 28632 36320 28684 36329
rect 28908 36320 28960 36372
rect 31300 36320 31352 36372
rect 34520 36320 34572 36372
rect 35440 36363 35492 36372
rect 35440 36329 35449 36363
rect 35449 36329 35483 36363
rect 35483 36329 35492 36363
rect 35440 36320 35492 36329
rect 22836 36252 22888 36304
rect 26240 36252 26292 36304
rect 27896 36252 27948 36304
rect 15292 36184 15344 36236
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 3056 36116 3108 36168
rect 4988 36116 5040 36168
rect 3148 36048 3200 36100
rect 7012 36116 7064 36168
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 8024 36116 8076 36168
rect 9220 36159 9272 36168
rect 9220 36125 9229 36159
rect 9229 36125 9263 36159
rect 9263 36125 9272 36159
rect 9220 36116 9272 36125
rect 10232 36159 10284 36168
rect 10232 36125 10241 36159
rect 10241 36125 10275 36159
rect 10275 36125 10284 36159
rect 10232 36116 10284 36125
rect 11704 36159 11756 36168
rect 6460 36048 6512 36100
rect 11704 36125 11713 36159
rect 11713 36125 11747 36159
rect 11747 36125 11756 36159
rect 11704 36116 11756 36125
rect 12256 36048 12308 36100
rect 13452 36116 13504 36168
rect 13912 36116 13964 36168
rect 14556 36116 14608 36168
rect 16856 36116 16908 36168
rect 17132 36116 17184 36168
rect 18052 36116 18104 36168
rect 12900 36048 12952 36100
rect 19984 36159 20036 36168
rect 19984 36125 19993 36159
rect 19993 36125 20027 36159
rect 20027 36125 20036 36159
rect 19984 36116 20036 36125
rect 20720 36116 20772 36168
rect 21916 36159 21968 36168
rect 21916 36125 21925 36159
rect 21925 36125 21959 36159
rect 21959 36125 21968 36159
rect 21916 36116 21968 36125
rect 20260 36048 20312 36100
rect 18052 35980 18104 36032
rect 23112 36048 23164 36100
rect 24860 36116 24912 36168
rect 26608 36116 26660 36168
rect 27068 36159 27120 36168
rect 27068 36125 27077 36159
rect 27077 36125 27111 36159
rect 27111 36125 27120 36159
rect 27068 36116 27120 36125
rect 27896 36048 27948 36100
rect 23204 35980 23256 36032
rect 23664 35980 23716 36032
rect 23848 35980 23900 36032
rect 29000 36184 29052 36236
rect 29552 36116 29604 36168
rect 30196 36159 30248 36168
rect 30196 36125 30205 36159
rect 30205 36125 30239 36159
rect 30239 36125 30248 36159
rect 30196 36116 30248 36125
rect 37464 36184 37516 36236
rect 37556 36227 37608 36236
rect 37556 36193 37565 36227
rect 37565 36193 37599 36227
rect 37599 36193 37608 36227
rect 37556 36184 37608 36193
rect 31668 36159 31720 36168
rect 31668 36125 31677 36159
rect 31677 36125 31711 36159
rect 31711 36125 31720 36159
rect 31668 36116 31720 36125
rect 34704 36159 34756 36168
rect 34704 36125 34713 36159
rect 34713 36125 34747 36159
rect 34747 36125 34756 36159
rect 34704 36116 34756 36125
rect 38476 36116 38528 36168
rect 30472 36048 30524 36100
rect 30932 36048 30984 36100
rect 32680 36048 32732 36100
rect 34152 36048 34204 36100
rect 28448 35980 28500 36032
rect 28908 35980 28960 36032
rect 30104 35980 30156 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 756 35776 808 35828
rect 3148 35776 3200 35828
rect 4068 35776 4120 35828
rect 5264 35776 5316 35828
rect 7104 35776 7156 35828
rect 8576 35819 8628 35828
rect 8576 35785 8585 35819
rect 8585 35785 8619 35819
rect 8619 35785 8628 35819
rect 8576 35776 8628 35785
rect 9312 35776 9364 35828
rect 10692 35776 10744 35828
rect 11704 35776 11756 35828
rect 14280 35776 14332 35828
rect 14832 35819 14884 35828
rect 14832 35785 14841 35819
rect 14841 35785 14875 35819
rect 14875 35785 14884 35819
rect 14832 35776 14884 35785
rect 15476 35776 15528 35828
rect 16672 35819 16724 35828
rect 16672 35785 16681 35819
rect 16681 35785 16715 35819
rect 16715 35785 16724 35819
rect 16672 35776 16724 35785
rect 16856 35776 16908 35828
rect 18696 35776 18748 35828
rect 19340 35776 19392 35828
rect 20904 35776 20956 35828
rect 22192 35776 22244 35828
rect 22928 35776 22980 35828
rect 23480 35776 23532 35828
rect 24308 35819 24360 35828
rect 24308 35785 24317 35819
rect 24317 35785 24351 35819
rect 24351 35785 24360 35819
rect 24308 35776 24360 35785
rect 26976 35776 27028 35828
rect 28816 35776 28868 35828
rect 29736 35776 29788 35828
rect 30288 35776 30340 35828
rect 31208 35819 31260 35828
rect 31208 35785 31217 35819
rect 31217 35785 31251 35819
rect 31251 35785 31260 35819
rect 31208 35776 31260 35785
rect 32404 35776 32456 35828
rect 35532 35776 35584 35828
rect 37280 35819 37332 35828
rect 37280 35785 37289 35819
rect 37289 35785 37323 35819
rect 37323 35785 37332 35819
rect 37280 35776 37332 35785
rect 27436 35708 27488 35760
rect 3148 35640 3200 35692
rect 3700 35640 3752 35692
rect 8852 35640 8904 35692
rect 11060 35640 11112 35692
rect 11704 35640 11756 35692
rect 12624 35640 12676 35692
rect 14188 35640 14240 35692
rect 14740 35640 14792 35692
rect 15936 35640 15988 35692
rect 16764 35640 16816 35692
rect 17868 35640 17920 35692
rect 11244 35572 11296 35624
rect 16672 35572 16724 35624
rect 22836 35640 22888 35692
rect 26148 35640 26200 35692
rect 26884 35640 26936 35692
rect 27160 35640 27212 35692
rect 30564 35708 30616 35760
rect 31300 35640 31352 35692
rect 32772 35683 32824 35692
rect 32772 35649 32781 35683
rect 32781 35649 32815 35683
rect 32815 35649 32824 35683
rect 32772 35640 32824 35649
rect 33968 35640 34020 35692
rect 34060 35683 34112 35692
rect 34060 35649 34069 35683
rect 34069 35649 34103 35683
rect 34103 35649 34112 35683
rect 34060 35640 34112 35649
rect 8116 35504 8168 35556
rect 22560 35504 22612 35556
rect 24952 35504 25004 35556
rect 35440 35640 35492 35692
rect 36360 35640 36412 35692
rect 37832 35640 37884 35692
rect 39028 35640 39080 35692
rect 35532 35572 35584 35624
rect 29460 35504 29512 35556
rect 33416 35504 33468 35556
rect 36544 35504 36596 35556
rect 37372 35504 37424 35556
rect 3700 35436 3752 35488
rect 5724 35479 5776 35488
rect 5724 35445 5733 35479
rect 5733 35445 5767 35479
rect 5767 35445 5776 35479
rect 5724 35436 5776 35445
rect 8024 35479 8076 35488
rect 8024 35445 8033 35479
rect 8033 35445 8067 35479
rect 8067 35445 8076 35479
rect 8024 35436 8076 35445
rect 12624 35436 12676 35488
rect 13452 35479 13504 35488
rect 13452 35445 13461 35479
rect 13461 35445 13495 35479
rect 13495 35445 13504 35479
rect 13452 35436 13504 35445
rect 17868 35436 17920 35488
rect 19984 35436 20036 35488
rect 20720 35479 20772 35488
rect 20720 35445 20729 35479
rect 20729 35445 20763 35479
rect 20763 35445 20772 35479
rect 20720 35436 20772 35445
rect 21916 35479 21968 35488
rect 21916 35445 21925 35479
rect 21925 35445 21959 35479
rect 21959 35445 21968 35479
rect 21916 35436 21968 35445
rect 24860 35479 24912 35488
rect 24860 35445 24869 35479
rect 24869 35445 24903 35479
rect 24903 35445 24912 35479
rect 24860 35436 24912 35445
rect 25412 35479 25464 35488
rect 25412 35445 25421 35479
rect 25421 35445 25455 35479
rect 25455 35445 25464 35479
rect 25412 35436 25464 35445
rect 28172 35479 28224 35488
rect 28172 35445 28181 35479
rect 28181 35445 28215 35479
rect 28215 35445 28224 35479
rect 28172 35436 28224 35445
rect 29644 35436 29696 35488
rect 38752 35436 38804 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1584 35275 1636 35284
rect 1584 35241 1593 35275
rect 1593 35241 1627 35275
rect 1627 35241 1636 35275
rect 1584 35232 1636 35241
rect 1768 35232 1820 35284
rect 6184 35275 6236 35284
rect 6184 35241 6193 35275
rect 6193 35241 6227 35275
rect 6227 35241 6236 35275
rect 6184 35232 6236 35241
rect 6736 35275 6788 35284
rect 6736 35241 6745 35275
rect 6745 35241 6779 35275
rect 6779 35241 6788 35275
rect 6736 35232 6788 35241
rect 7472 35232 7524 35284
rect 9588 35232 9640 35284
rect 10140 35232 10192 35284
rect 10232 35232 10284 35284
rect 12164 35275 12216 35284
rect 12164 35241 12173 35275
rect 12173 35241 12207 35275
rect 12207 35241 12216 35275
rect 12164 35232 12216 35241
rect 12716 35275 12768 35284
rect 12716 35241 12725 35275
rect 12725 35241 12759 35275
rect 12759 35241 12768 35275
rect 12716 35232 12768 35241
rect 15384 35232 15436 35284
rect 17500 35275 17552 35284
rect 17500 35241 17509 35275
rect 17509 35241 17543 35275
rect 17543 35241 17552 35275
rect 17500 35232 17552 35241
rect 17960 35232 18012 35284
rect 18604 35275 18656 35284
rect 18604 35241 18613 35275
rect 18613 35241 18647 35275
rect 18647 35241 18656 35275
rect 18604 35232 18656 35241
rect 19248 35275 19300 35284
rect 19248 35241 19257 35275
rect 19257 35241 19291 35275
rect 19291 35241 19300 35275
rect 19248 35232 19300 35241
rect 20076 35275 20128 35284
rect 20076 35241 20085 35275
rect 20085 35241 20119 35275
rect 20119 35241 20128 35275
rect 20076 35232 20128 35241
rect 29552 35275 29604 35284
rect 29552 35241 29561 35275
rect 29561 35241 29595 35275
rect 29595 35241 29604 35275
rect 29552 35232 29604 35241
rect 33508 35275 33560 35284
rect 33508 35241 33517 35275
rect 33517 35241 33551 35275
rect 33551 35241 33560 35275
rect 33508 35232 33560 35241
rect 35624 35232 35676 35284
rect 38292 35232 38344 35284
rect 1676 35164 1728 35216
rect 28172 35164 28224 35216
rect 25504 35096 25556 35148
rect 28448 35096 28500 35148
rect 10600 35071 10652 35080
rect 10600 35037 10609 35071
rect 10609 35037 10643 35071
rect 10643 35037 10652 35071
rect 10600 35028 10652 35037
rect 15108 35071 15160 35080
rect 15108 35037 15117 35071
rect 15117 35037 15151 35071
rect 15151 35037 15160 35071
rect 15108 35028 15160 35037
rect 15752 35071 15804 35080
rect 15752 35037 15761 35071
rect 15761 35037 15795 35071
rect 15795 35037 15804 35071
rect 15752 35028 15804 35037
rect 13360 35003 13412 35012
rect 13360 34969 13369 35003
rect 13369 34969 13403 35003
rect 13403 34969 13412 35003
rect 29644 35028 29696 35080
rect 35992 35071 36044 35080
rect 13360 34960 13412 34969
rect 20444 34960 20496 35012
rect 26240 34960 26292 35012
rect 30564 34960 30616 35012
rect 31668 34960 31720 35012
rect 3884 34935 3936 34944
rect 3884 34901 3893 34935
rect 3893 34901 3927 34935
rect 3927 34901 3936 34935
rect 3884 34892 3936 34901
rect 4712 34892 4764 34944
rect 5080 34892 5132 34944
rect 5540 34935 5592 34944
rect 5540 34901 5549 34935
rect 5549 34901 5583 34935
rect 5583 34901 5592 34935
rect 5540 34892 5592 34901
rect 7104 34892 7156 34944
rect 8852 34892 8904 34944
rect 11060 34935 11112 34944
rect 11060 34901 11069 34935
rect 11069 34901 11103 34935
rect 11103 34901 11112 34935
rect 11060 34892 11112 34901
rect 11704 34935 11756 34944
rect 11704 34901 11713 34935
rect 11713 34901 11747 34935
rect 11747 34901 11756 34935
rect 11704 34892 11756 34901
rect 14188 34892 14240 34944
rect 16764 34892 16816 34944
rect 19432 34892 19484 34944
rect 20536 34935 20588 34944
rect 20536 34901 20545 34935
rect 20545 34901 20579 34935
rect 20579 34901 20588 34935
rect 20536 34892 20588 34901
rect 21088 34935 21140 34944
rect 21088 34901 21097 34935
rect 21097 34901 21131 34935
rect 21131 34901 21140 34935
rect 21088 34892 21140 34901
rect 22192 34892 22244 34944
rect 22836 34935 22888 34944
rect 22836 34901 22845 34935
rect 22845 34901 22879 34935
rect 22879 34901 22888 34935
rect 22836 34892 22888 34901
rect 26332 34892 26384 34944
rect 29920 34935 29972 34944
rect 29920 34901 29929 34935
rect 29929 34901 29963 34935
rect 29963 34901 29972 34935
rect 29920 34892 29972 34901
rect 30380 34892 30432 34944
rect 31024 34892 31076 34944
rect 31944 34935 31996 34944
rect 31944 34901 31953 34935
rect 31953 34901 31987 34935
rect 31987 34901 31996 34935
rect 31944 34892 31996 34901
rect 32772 34892 32824 34944
rect 33232 34892 33284 34944
rect 34244 34892 34296 34944
rect 34704 34935 34756 34944
rect 34704 34901 34713 34935
rect 34713 34901 34747 34935
rect 34747 34901 34756 34935
rect 34704 34892 34756 34901
rect 35992 35037 36001 35071
rect 36001 35037 36035 35071
rect 36035 35037 36044 35071
rect 35992 35028 36044 35037
rect 36084 35028 36136 35080
rect 37280 35028 37332 35080
rect 38292 35028 38344 35080
rect 36452 34960 36504 35012
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2596 34731 2648 34740
rect 2596 34697 2605 34731
rect 2605 34697 2639 34731
rect 2639 34697 2648 34731
rect 2596 34688 2648 34697
rect 9220 34731 9272 34740
rect 9220 34697 9229 34731
rect 9229 34697 9263 34731
rect 9263 34697 9272 34731
rect 9220 34688 9272 34697
rect 12256 34688 12308 34740
rect 12900 34731 12952 34740
rect 12900 34697 12909 34731
rect 12909 34697 12943 34731
rect 12943 34697 12952 34731
rect 12900 34688 12952 34697
rect 15108 34688 15160 34740
rect 16948 34731 17000 34740
rect 16948 34697 16957 34731
rect 16957 34697 16991 34731
rect 16991 34697 17000 34731
rect 16948 34688 17000 34697
rect 20260 34688 20312 34740
rect 3056 34620 3108 34672
rect 2872 34484 2924 34536
rect 3240 34484 3292 34536
rect 4160 34484 4212 34536
rect 9496 34620 9548 34672
rect 19064 34620 19116 34672
rect 19984 34620 20036 34672
rect 5264 34552 5316 34604
rect 13912 34595 13964 34604
rect 13912 34561 13921 34595
rect 13921 34561 13955 34595
rect 13955 34561 13964 34595
rect 13912 34552 13964 34561
rect 14280 34552 14332 34604
rect 14556 34595 14608 34604
rect 14556 34561 14565 34595
rect 14565 34561 14599 34595
rect 14599 34561 14608 34595
rect 14556 34552 14608 34561
rect 14740 34552 14792 34604
rect 18328 34595 18380 34604
rect 18328 34561 18362 34595
rect 18362 34561 18380 34595
rect 18328 34552 18380 34561
rect 9772 34527 9824 34536
rect 9772 34493 9781 34527
rect 9781 34493 9815 34527
rect 9815 34493 9824 34527
rect 9772 34484 9824 34493
rect 10600 34484 10652 34536
rect 11244 34484 11296 34536
rect 13728 34484 13780 34536
rect 20260 34484 20312 34536
rect 23848 34688 23900 34740
rect 27160 34688 27212 34740
rect 35808 34688 35860 34740
rect 23112 34620 23164 34672
rect 26240 34620 26292 34672
rect 27528 34620 27580 34672
rect 37280 34688 37332 34740
rect 37924 34688 37976 34740
rect 39396 34688 39448 34740
rect 37188 34620 37240 34672
rect 39764 34620 39816 34672
rect 35256 34595 35308 34604
rect 35256 34561 35265 34595
rect 35265 34561 35299 34595
rect 35299 34561 35308 34595
rect 35256 34552 35308 34561
rect 36176 34552 36228 34604
rect 37556 34552 37608 34604
rect 25504 34484 25556 34536
rect 32956 34527 33008 34536
rect 32956 34493 32965 34527
rect 32965 34493 32999 34527
rect 32999 34493 33008 34527
rect 32956 34484 33008 34493
rect 33968 34484 34020 34536
rect 36912 34484 36964 34536
rect 5816 34391 5868 34400
rect 5816 34357 5825 34391
rect 5825 34357 5859 34391
rect 5859 34357 5868 34391
rect 5816 34348 5868 34357
rect 19432 34391 19484 34400
rect 19432 34357 19441 34391
rect 19441 34357 19475 34391
rect 19475 34357 19484 34391
rect 19432 34348 19484 34357
rect 22376 34391 22428 34400
rect 22376 34357 22385 34391
rect 22385 34357 22419 34391
rect 22419 34357 22428 34391
rect 23940 34416 23992 34468
rect 22376 34348 22428 34357
rect 35808 34348 35860 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 18052 34187 18104 34196
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 31300 34187 31352 34196
rect 31300 34153 31309 34187
rect 31309 34153 31343 34187
rect 31343 34153 31352 34187
rect 31300 34144 31352 34153
rect 35992 34144 36044 34196
rect 36084 34144 36136 34196
rect 37188 34187 37240 34196
rect 37188 34153 37197 34187
rect 37197 34153 37231 34187
rect 37231 34153 37240 34187
rect 37188 34144 37240 34153
rect 37648 34144 37700 34196
rect 9496 33940 9548 33992
rect 10140 33872 10192 33924
rect 10784 33847 10836 33856
rect 10784 33813 10793 33847
rect 10793 33813 10827 33847
rect 10827 33813 10836 33847
rect 10784 33804 10836 33813
rect 32128 33940 32180 33992
rect 36728 34008 36780 34060
rect 36636 33940 36688 33992
rect 37740 33983 37792 33992
rect 37740 33949 37749 33983
rect 37749 33949 37783 33983
rect 37783 33949 37792 33983
rect 37740 33940 37792 33949
rect 13728 33804 13780 33856
rect 15936 33847 15988 33856
rect 15936 33813 15945 33847
rect 15945 33813 15979 33847
rect 15979 33813 15988 33847
rect 15936 33804 15988 33813
rect 17132 33847 17184 33856
rect 17132 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17184 33847
rect 17132 33804 17184 33813
rect 23940 33804 23992 33856
rect 33600 33804 33652 33856
rect 34060 33804 34112 33856
rect 34612 33804 34664 33856
rect 35440 33804 35492 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 5264 33643 5316 33652
rect 5264 33609 5273 33643
rect 5273 33609 5307 33643
rect 5307 33609 5316 33643
rect 5264 33600 5316 33609
rect 10140 33643 10192 33652
rect 10140 33609 10149 33643
rect 10149 33609 10183 33643
rect 10183 33609 10192 33643
rect 10140 33600 10192 33609
rect 10784 33600 10836 33652
rect 11796 33600 11848 33652
rect 18328 33600 18380 33652
rect 29368 33643 29420 33652
rect 29368 33609 29377 33643
rect 29377 33609 29411 33643
rect 29411 33609 29420 33643
rect 29368 33600 29420 33609
rect 36728 33643 36780 33652
rect 36728 33609 36737 33643
rect 36737 33609 36771 33643
rect 36771 33609 36780 33643
rect 36728 33600 36780 33609
rect 37832 33600 37884 33652
rect 38660 33600 38712 33652
rect 6828 33464 6880 33516
rect 4896 33396 4948 33448
rect 5172 33396 5224 33448
rect 5816 33396 5868 33448
rect 6368 33396 6420 33448
rect 4804 33260 4856 33312
rect 7656 33260 7708 33312
rect 10784 33464 10836 33516
rect 19524 33464 19576 33516
rect 27528 33507 27580 33516
rect 27528 33473 27537 33507
rect 27537 33473 27571 33507
rect 27571 33473 27580 33507
rect 27528 33464 27580 33473
rect 29184 33507 29236 33516
rect 29184 33473 29193 33507
rect 29193 33473 29227 33507
rect 29227 33473 29236 33507
rect 29184 33464 29236 33473
rect 37832 33507 37884 33516
rect 37832 33473 37841 33507
rect 37841 33473 37875 33507
rect 37875 33473 37884 33507
rect 37832 33464 37884 33473
rect 19432 33396 19484 33448
rect 27804 33439 27856 33448
rect 27804 33405 27813 33439
rect 27813 33405 27847 33439
rect 27847 33405 27856 33439
rect 27804 33396 27856 33405
rect 19340 33328 19392 33380
rect 19248 33260 19300 33312
rect 35532 33260 35584 33312
rect 36360 33260 36412 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19524 33099 19576 33108
rect 19524 33065 19533 33099
rect 19533 33065 19567 33099
rect 19567 33065 19576 33099
rect 19524 33056 19576 33065
rect 28448 33031 28500 33040
rect 28448 32997 28457 33031
rect 28457 32997 28491 33031
rect 28491 32997 28500 33031
rect 28448 32988 28500 32997
rect 19248 32895 19300 32904
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 19432 32852 19484 32904
rect 27804 32852 27856 32904
rect 32864 32852 32916 32904
rect 38108 32895 38160 32904
rect 38108 32861 38117 32895
rect 38117 32861 38151 32895
rect 38151 32861 38160 32895
rect 38108 32852 38160 32861
rect 19340 32716 19392 32768
rect 19984 32759 20036 32768
rect 19984 32725 19993 32759
rect 19993 32725 20027 32759
rect 20027 32725 20036 32759
rect 19984 32716 20036 32725
rect 36544 32716 36596 32768
rect 36912 32716 36964 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 6828 32555 6880 32564
rect 6828 32521 6837 32555
rect 6837 32521 6871 32555
rect 6871 32521 6880 32555
rect 6828 32512 6880 32521
rect 26148 32555 26200 32564
rect 26148 32521 26157 32555
rect 26157 32521 26191 32555
rect 26191 32521 26200 32555
rect 26148 32512 26200 32521
rect 32128 32555 32180 32564
rect 32128 32521 32137 32555
rect 32137 32521 32171 32555
rect 32171 32521 32180 32555
rect 32128 32512 32180 32521
rect 38108 32487 38160 32496
rect 38108 32453 38117 32487
rect 38117 32453 38151 32487
rect 38151 32453 38160 32487
rect 38108 32444 38160 32453
rect 7656 32376 7708 32428
rect 13728 32376 13780 32428
rect 14372 32419 14424 32428
rect 14372 32385 14406 32419
rect 14406 32385 14424 32419
rect 14372 32376 14424 32385
rect 25320 32376 25372 32428
rect 26240 32376 26292 32428
rect 18788 32240 18840 32292
rect 34244 32376 34296 32428
rect 32864 32308 32916 32360
rect 7472 32215 7524 32224
rect 7472 32181 7481 32215
rect 7481 32181 7515 32215
rect 7515 32181 7524 32215
rect 7472 32172 7524 32181
rect 15200 32172 15252 32224
rect 25320 32215 25372 32224
rect 25320 32181 25329 32215
rect 25329 32181 25363 32215
rect 25363 32181 25372 32215
rect 25320 32172 25372 32181
rect 37740 32172 37792 32224
rect 38660 32172 38712 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 26608 31968 26660 32020
rect 29184 31968 29236 32020
rect 26240 31832 26292 31884
rect 25872 31764 25924 31816
rect 27528 31832 27580 31884
rect 26700 31764 26752 31816
rect 28448 31764 28500 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 33048 31288 33100 31340
rect 35992 31356 36044 31408
rect 36452 31331 36504 31340
rect 36452 31297 36470 31331
rect 36470 31297 36504 31331
rect 36452 31288 36504 31297
rect 38108 31331 38160 31340
rect 38108 31297 38117 31331
rect 38117 31297 38151 31331
rect 38151 31297 38160 31331
rect 38108 31288 38160 31297
rect 34244 31152 34296 31204
rect 33140 31084 33192 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 27068 30923 27120 30932
rect 27068 30889 27077 30923
rect 27077 30889 27111 30923
rect 27111 30889 27120 30923
rect 27068 30880 27120 30889
rect 33048 30923 33100 30932
rect 33048 30889 33057 30923
rect 33057 30889 33091 30923
rect 33091 30889 33100 30923
rect 33048 30880 33100 30889
rect 34428 30880 34480 30932
rect 35992 30880 36044 30932
rect 27528 30812 27580 30864
rect 32864 30855 32916 30864
rect 32864 30821 32873 30855
rect 32873 30821 32907 30855
rect 32907 30821 32916 30855
rect 32864 30812 32916 30821
rect 4068 30676 4120 30728
rect 4804 30719 4856 30728
rect 4804 30685 4813 30719
rect 4813 30685 4847 30719
rect 4847 30685 4856 30719
rect 4804 30676 4856 30685
rect 3608 30608 3660 30660
rect 4068 30540 4120 30592
rect 4896 30583 4948 30592
rect 4896 30549 4905 30583
rect 4905 30549 4939 30583
rect 4939 30549 4948 30583
rect 4896 30540 4948 30549
rect 22744 30608 22796 30660
rect 37188 30676 37240 30728
rect 27160 30608 27212 30660
rect 32588 30651 32640 30660
rect 32588 30617 32597 30651
rect 32597 30617 32631 30651
rect 32631 30617 32640 30651
rect 32588 30608 32640 30617
rect 6920 30540 6972 30592
rect 7472 30540 7524 30592
rect 8208 30540 8260 30592
rect 22284 30583 22336 30592
rect 22284 30549 22293 30583
rect 22293 30549 22327 30583
rect 22327 30549 22336 30583
rect 22284 30540 22336 30549
rect 27344 30540 27396 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4804 30336 4856 30388
rect 3608 30311 3660 30320
rect 3608 30277 3617 30311
rect 3617 30277 3651 30311
rect 3651 30277 3660 30311
rect 3608 30268 3660 30277
rect 1584 30200 1636 30252
rect 4896 30200 4948 30252
rect 5632 30268 5684 30320
rect 6368 30311 6420 30320
rect 6368 30277 6377 30311
rect 6377 30277 6411 30311
rect 6411 30277 6420 30311
rect 6368 30268 6420 30277
rect 7656 30268 7708 30320
rect 10968 30268 11020 30320
rect 11520 30311 11572 30320
rect 11520 30277 11529 30311
rect 11529 30277 11563 30311
rect 11563 30277 11572 30311
rect 11888 30336 11940 30388
rect 15384 30336 15436 30388
rect 22744 30379 22796 30388
rect 22744 30345 22753 30379
rect 22753 30345 22787 30379
rect 22787 30345 22796 30379
rect 22744 30336 22796 30345
rect 32404 30379 32456 30388
rect 32404 30345 32413 30379
rect 32413 30345 32447 30379
rect 32447 30345 32456 30379
rect 32404 30336 32456 30345
rect 32588 30336 32640 30388
rect 11520 30268 11572 30277
rect 4068 30175 4120 30184
rect 4068 30141 4077 30175
rect 4077 30141 4111 30175
rect 4111 30141 4120 30175
rect 14372 30311 14424 30320
rect 14372 30277 14381 30311
rect 14381 30277 14415 30311
rect 14415 30277 14424 30311
rect 14372 30268 14424 30277
rect 4068 30132 4120 30141
rect 6184 30064 6236 30116
rect 4804 29996 4856 30048
rect 4896 29996 4948 30048
rect 11428 30132 11480 30184
rect 11612 30064 11664 30116
rect 15200 30200 15252 30252
rect 15384 30243 15436 30252
rect 15384 30209 15393 30243
rect 15393 30209 15427 30243
rect 15427 30209 15436 30243
rect 15384 30200 15436 30209
rect 19248 30268 19300 30320
rect 15476 30132 15528 30184
rect 17500 30175 17552 30184
rect 17500 30141 17509 30175
rect 17509 30141 17543 30175
rect 17543 30141 17552 30175
rect 17500 30132 17552 30141
rect 18696 30200 18748 30252
rect 19432 30268 19484 30320
rect 32036 30268 32088 30320
rect 33140 30268 33192 30320
rect 20168 30243 20220 30252
rect 20168 30209 20177 30243
rect 20177 30209 20211 30243
rect 20211 30209 20220 30243
rect 20168 30200 20220 30209
rect 22928 30200 22980 30252
rect 30288 30200 30340 30252
rect 19432 30132 19484 30184
rect 22284 30175 22336 30184
rect 22284 30141 22293 30175
rect 22293 30141 22327 30175
rect 22327 30141 22336 30175
rect 22284 30132 22336 30141
rect 32128 30175 32180 30184
rect 32128 30141 32137 30175
rect 32137 30141 32171 30175
rect 32171 30141 32180 30175
rect 32128 30132 32180 30141
rect 18328 30064 18380 30116
rect 11796 29996 11848 30048
rect 15476 29996 15528 30048
rect 18420 29996 18472 30048
rect 19432 29996 19484 30048
rect 22284 29996 22336 30048
rect 30840 29996 30892 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 8208 29792 8260 29844
rect 15384 29792 15436 29844
rect 17500 29792 17552 29844
rect 20168 29792 20220 29844
rect 32864 29792 32916 29844
rect 37188 29792 37240 29844
rect 9496 29724 9548 29776
rect 11520 29724 11572 29776
rect 10968 29588 11020 29640
rect 11796 29588 11848 29640
rect 22284 29588 22336 29640
rect 10140 29520 10192 29572
rect 11336 29563 11388 29572
rect 11336 29529 11345 29563
rect 11345 29529 11379 29563
rect 11379 29529 11388 29563
rect 11336 29520 11388 29529
rect 25228 29563 25280 29572
rect 25228 29529 25237 29563
rect 25237 29529 25271 29563
rect 25271 29529 25280 29563
rect 25228 29520 25280 29529
rect 31576 29588 31628 29640
rect 32404 29699 32456 29708
rect 32404 29665 32413 29699
rect 32413 29665 32447 29699
rect 32447 29665 32456 29699
rect 32404 29656 32456 29665
rect 32588 29656 32640 29708
rect 32036 29588 32088 29640
rect 38108 29631 38160 29640
rect 32128 29520 32180 29572
rect 38108 29597 38117 29631
rect 38117 29597 38151 29631
rect 38151 29597 38160 29631
rect 38108 29588 38160 29597
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9496 29248 9548 29300
rect 22928 29291 22980 29300
rect 22928 29257 22937 29291
rect 22937 29257 22971 29291
rect 22971 29257 22980 29291
rect 22928 29248 22980 29257
rect 8392 29112 8444 29164
rect 11520 29155 11572 29164
rect 11520 29121 11529 29155
rect 11529 29121 11563 29155
rect 11563 29121 11572 29155
rect 11520 29112 11572 29121
rect 11612 29155 11664 29164
rect 11612 29121 11621 29155
rect 11621 29121 11655 29155
rect 11655 29121 11664 29155
rect 11612 29112 11664 29121
rect 15384 29112 15436 29164
rect 25228 29112 25280 29164
rect 30288 29112 30340 29164
rect 13084 29044 13136 29096
rect 11336 28976 11388 29028
rect 31576 28976 31628 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6184 28747 6236 28756
rect 6184 28713 6193 28747
rect 6193 28713 6227 28747
rect 6227 28713 6236 28747
rect 6184 28704 6236 28713
rect 6920 28747 6972 28756
rect 6920 28713 6929 28747
rect 6929 28713 6963 28747
rect 6963 28713 6972 28747
rect 6920 28704 6972 28713
rect 18328 28679 18380 28688
rect 18328 28645 18337 28679
rect 18337 28645 18371 28679
rect 18371 28645 18380 28679
rect 18328 28636 18380 28645
rect 6184 28500 6236 28552
rect 6736 28543 6788 28552
rect 6736 28509 6745 28543
rect 6745 28509 6779 28543
rect 6779 28509 6788 28543
rect 6736 28500 6788 28509
rect 18420 28543 18472 28552
rect 18420 28509 18429 28543
rect 18429 28509 18463 28543
rect 18463 28509 18472 28543
rect 18420 28500 18472 28509
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 29000 28432 29052 28484
rect 18420 28407 18472 28416
rect 17592 28364 17644 28373
rect 18420 28373 18429 28407
rect 18429 28373 18463 28407
rect 18463 28373 18472 28407
rect 18420 28364 18472 28373
rect 26424 28364 26476 28416
rect 30748 28407 30800 28416
rect 30748 28373 30757 28407
rect 30757 28373 30791 28407
rect 30791 28373 30800 28407
rect 30748 28364 30800 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 30288 28160 30340 28212
rect 31576 28160 31628 28212
rect 30748 28092 30800 28144
rect 34428 28092 34480 28144
rect 25228 28024 25280 28076
rect 26148 28067 26200 28076
rect 26148 28033 26157 28067
rect 26157 28033 26191 28067
rect 26191 28033 26200 28067
rect 26148 28024 26200 28033
rect 26240 28067 26292 28076
rect 26240 28033 26249 28067
rect 26249 28033 26283 28067
rect 26283 28033 26292 28067
rect 26424 28067 26476 28076
rect 26240 28024 26292 28033
rect 26424 28033 26433 28067
rect 26433 28033 26467 28067
rect 26467 28033 26476 28067
rect 26424 28024 26476 28033
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 27436 28067 27488 28076
rect 27436 28033 27470 28067
rect 27470 28033 27488 28067
rect 27436 28024 27488 28033
rect 31760 28024 31812 28076
rect 32588 28024 32640 28076
rect 38108 28067 38160 28076
rect 38108 28033 38117 28067
rect 38117 28033 38151 28067
rect 38151 28033 38160 28067
rect 38108 28024 38160 28033
rect 27068 27820 27120 27872
rect 32404 27863 32456 27872
rect 32404 27829 32413 27863
rect 32413 27829 32447 27863
rect 32447 27829 32456 27863
rect 32404 27820 32456 27829
rect 34796 27820 34848 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 27436 27616 27488 27668
rect 4804 27591 4856 27600
rect 4804 27557 4813 27591
rect 4813 27557 4847 27591
rect 4847 27557 4856 27591
rect 4804 27548 4856 27557
rect 5632 27480 5684 27532
rect 4804 27412 4856 27464
rect 6920 27548 6972 27600
rect 18696 27591 18748 27600
rect 18696 27557 18705 27591
rect 18705 27557 18739 27591
rect 18739 27557 18748 27591
rect 18696 27548 18748 27557
rect 26148 27548 26200 27600
rect 31760 27616 31812 27668
rect 32588 27548 32640 27600
rect 34428 27548 34480 27600
rect 37556 27591 37608 27600
rect 31760 27523 31812 27532
rect 31760 27489 31769 27523
rect 31769 27489 31803 27523
rect 31803 27489 31812 27523
rect 31760 27480 31812 27489
rect 37556 27557 37565 27591
rect 37565 27557 37599 27591
rect 37599 27557 37608 27591
rect 37556 27548 37608 27557
rect 4896 27344 4948 27396
rect 5356 27319 5408 27328
rect 5356 27285 5365 27319
rect 5365 27285 5399 27319
rect 5399 27285 5408 27319
rect 5356 27276 5408 27285
rect 15476 27276 15528 27328
rect 18420 27412 18472 27464
rect 26240 27412 26292 27464
rect 27068 27412 27120 27464
rect 30840 27412 30892 27464
rect 31576 27455 31628 27464
rect 31576 27421 31585 27455
rect 31585 27421 31619 27455
rect 31619 27421 31628 27455
rect 32404 27455 32456 27464
rect 31576 27412 31628 27421
rect 32404 27421 32413 27455
rect 32413 27421 32447 27455
rect 32447 27421 32456 27455
rect 32404 27412 32456 27421
rect 35716 27480 35768 27532
rect 36268 27344 36320 27396
rect 30840 27319 30892 27328
rect 30840 27285 30849 27319
rect 30849 27285 30883 27319
rect 30883 27285 30892 27319
rect 30840 27276 30892 27285
rect 32496 27319 32548 27328
rect 32496 27285 32505 27319
rect 32505 27285 32539 27319
rect 32539 27285 32548 27319
rect 32496 27276 32548 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 34428 27072 34480 27124
rect 32496 27004 32548 27056
rect 36268 27004 36320 27056
rect 15844 26936 15896 26988
rect 35716 26979 35768 26988
rect 35716 26945 35725 26979
rect 35725 26945 35759 26979
rect 35759 26945 35768 26979
rect 35716 26936 35768 26945
rect 16580 26868 16632 26920
rect 16764 26868 16816 26920
rect 13084 26732 13136 26784
rect 17592 26800 17644 26852
rect 32588 26800 32640 26852
rect 15844 26775 15896 26784
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 15844 26732 15896 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5632 26528 5684 26580
rect 15844 26528 15896 26580
rect 30840 26528 30892 26580
rect 5356 26392 5408 26444
rect 4252 26367 4304 26376
rect 4252 26333 4261 26367
rect 4261 26333 4295 26367
rect 4295 26333 4304 26367
rect 4252 26324 4304 26333
rect 4896 26324 4948 26376
rect 3792 26231 3844 26240
rect 3792 26197 3801 26231
rect 3801 26197 3835 26231
rect 3835 26197 3844 26231
rect 3792 26188 3844 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4160 25984 4212 26036
rect 8392 25984 8444 26036
rect 26424 25984 26476 26036
rect 30840 26027 30892 26036
rect 30840 25993 30849 26027
rect 30849 25993 30883 26027
rect 30883 25993 30892 26027
rect 30840 25984 30892 25993
rect 3792 25848 3844 25900
rect 27160 25916 27212 25968
rect 22100 25891 22152 25900
rect 22100 25857 22134 25891
rect 22134 25857 22152 25891
rect 30748 25959 30800 25968
rect 30748 25925 30757 25959
rect 30757 25925 30791 25959
rect 30791 25925 30800 25959
rect 30748 25916 30800 25925
rect 22100 25848 22152 25857
rect 8392 25712 8444 25764
rect 15476 25712 15528 25764
rect 38108 25755 38160 25764
rect 14464 25644 14516 25696
rect 38108 25721 38117 25755
rect 38117 25721 38151 25755
rect 38151 25721 38160 25755
rect 38108 25712 38160 25721
rect 23112 25644 23164 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 13084 25483 13136 25492
rect 8392 25236 8444 25288
rect 11520 25372 11572 25424
rect 13084 25449 13093 25483
rect 13093 25449 13127 25483
rect 13127 25449 13136 25483
rect 13084 25440 13136 25449
rect 22100 25440 22152 25492
rect 14464 25372 14516 25424
rect 15476 25347 15528 25356
rect 15476 25313 15485 25347
rect 15485 25313 15519 25347
rect 15519 25313 15528 25347
rect 15476 25304 15528 25313
rect 23112 25279 23164 25288
rect 7932 25168 7984 25220
rect 6736 25100 6788 25152
rect 10968 25168 11020 25220
rect 12992 25168 13044 25220
rect 22008 25168 22060 25220
rect 23112 25245 23121 25279
rect 23121 25245 23155 25279
rect 23155 25245 23164 25279
rect 23112 25236 23164 25245
rect 30932 25440 30984 25492
rect 31392 25304 31444 25356
rect 23296 25236 23348 25288
rect 34796 25236 34848 25288
rect 29000 25211 29052 25220
rect 9680 25143 9732 25152
rect 9680 25109 9689 25143
rect 9689 25109 9723 25143
rect 9723 25109 9732 25143
rect 9680 25100 9732 25109
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 19984 25100 20036 25152
rect 25688 25100 25740 25152
rect 26424 25100 26476 25152
rect 28172 25143 28224 25152
rect 28172 25109 28181 25143
rect 28181 25109 28215 25143
rect 28215 25109 28224 25143
rect 29000 25177 29009 25211
rect 29009 25177 29043 25211
rect 29043 25177 29052 25211
rect 29000 25168 29052 25177
rect 31576 25168 31628 25220
rect 28172 25100 28224 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7932 24939 7984 24948
rect 7932 24905 7941 24939
rect 7941 24905 7975 24939
rect 7975 24905 7984 24939
rect 7932 24896 7984 24905
rect 11520 24896 11572 24948
rect 12992 24939 13044 24948
rect 12992 24905 13001 24939
rect 13001 24905 13035 24939
rect 13035 24905 13044 24939
rect 12992 24896 13044 24905
rect 9680 24828 9732 24880
rect 10968 24760 11020 24812
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 12348 24828 12400 24880
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 12440 24692 12492 24744
rect 10140 24667 10192 24676
rect 10140 24633 10149 24667
rect 10149 24633 10183 24667
rect 10183 24633 10192 24667
rect 10140 24624 10192 24633
rect 13084 24760 13136 24812
rect 14096 24760 14148 24812
rect 20904 24760 20956 24812
rect 28172 24760 28224 24812
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 12440 24352 12492 24404
rect 20904 24395 20956 24404
rect 20904 24361 20913 24395
rect 20913 24361 20947 24395
rect 20947 24361 20956 24395
rect 20904 24352 20956 24361
rect 25688 24395 25740 24404
rect 25688 24361 25697 24395
rect 25697 24361 25731 24395
rect 25731 24361 25740 24395
rect 25688 24352 25740 24361
rect 8852 24284 8904 24336
rect 8024 24216 8076 24268
rect 10968 24148 11020 24200
rect 14096 24148 14148 24200
rect 23296 24148 23348 24200
rect 25688 24148 25740 24200
rect 31392 24148 31444 24200
rect 19432 24080 19484 24132
rect 30104 24080 30156 24132
rect 30840 24080 30892 24132
rect 38016 24123 38068 24132
rect 38016 24089 38025 24123
rect 38025 24089 38059 24123
rect 38059 24089 38068 24123
rect 38016 24080 38068 24089
rect 12532 24012 12584 24064
rect 25136 24055 25188 24064
rect 25136 24021 25145 24055
rect 25145 24021 25179 24055
rect 25179 24021 25188 24055
rect 25136 24012 25188 24021
rect 37924 24055 37976 24064
rect 37924 24021 37933 24055
rect 37933 24021 37967 24055
rect 37967 24021 37976 24055
rect 37924 24012 37976 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 37464 23808 37516 23860
rect 37556 23808 37608 23860
rect 10600 23740 10652 23792
rect 31392 23783 31444 23792
rect 31392 23749 31401 23783
rect 31401 23749 31435 23783
rect 31435 23749 31444 23783
rect 31392 23740 31444 23749
rect 18052 23672 18104 23724
rect 37648 23715 37700 23724
rect 20628 23536 20680 23588
rect 16764 23511 16816 23520
rect 16764 23477 16773 23511
rect 16773 23477 16807 23511
rect 16807 23477 16816 23511
rect 16764 23468 16816 23477
rect 19432 23511 19484 23520
rect 19432 23477 19441 23511
rect 19441 23477 19475 23511
rect 19475 23477 19484 23511
rect 19432 23468 19484 23477
rect 30104 23511 30156 23520
rect 30104 23477 30113 23511
rect 30113 23477 30147 23511
rect 30147 23477 30156 23511
rect 30104 23468 30156 23477
rect 37648 23681 37657 23715
rect 37657 23681 37691 23715
rect 37691 23681 37700 23715
rect 37648 23672 37700 23681
rect 35900 23604 35952 23656
rect 32312 23468 32364 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 17592 23264 17644 23316
rect 18052 23307 18104 23316
rect 18052 23273 18061 23307
rect 18061 23273 18095 23307
rect 18095 23273 18104 23307
rect 18052 23264 18104 23273
rect 17684 23128 17736 23180
rect 17960 23103 18012 23112
rect 17960 23069 17969 23103
rect 17969 23069 18003 23103
rect 18003 23069 18012 23103
rect 17960 23060 18012 23069
rect 31392 23128 31444 23180
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 28264 23060 28316 23112
rect 32404 23060 32456 23112
rect 20628 22992 20680 23044
rect 22008 22992 22060 23044
rect 26056 23035 26108 23044
rect 26056 23001 26090 23035
rect 26090 23001 26108 23035
rect 26056 22992 26108 23001
rect 27252 22924 27304 22976
rect 37556 22967 37608 22976
rect 37556 22933 37565 22967
rect 37565 22933 37599 22967
rect 37599 22933 37608 22967
rect 37556 22924 37608 22933
rect 37648 22924 37700 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 20536 22720 20588 22772
rect 20628 22652 20680 22704
rect 26056 22720 26108 22772
rect 32680 22720 32732 22772
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 25136 22584 25188 22636
rect 32680 22584 32732 22636
rect 34796 22584 34848 22636
rect 35900 22652 35952 22704
rect 37556 22652 37608 22704
rect 38200 22652 38252 22704
rect 27252 22516 27304 22568
rect 32128 22516 32180 22568
rect 32404 22516 32456 22568
rect 37924 22516 37976 22568
rect 17224 22448 17276 22500
rect 20996 22380 21048 22432
rect 26424 22380 26476 22432
rect 32036 22380 32088 22432
rect 32680 22423 32732 22432
rect 32680 22389 32689 22423
rect 32689 22389 32723 22423
rect 32723 22389 32732 22423
rect 32680 22380 32732 22389
rect 36084 22423 36136 22432
rect 36084 22389 36093 22423
rect 36093 22389 36127 22423
rect 36127 22389 36136 22423
rect 36084 22380 36136 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6920 22040 6972 22092
rect 17960 22040 18012 22092
rect 21272 22040 21324 22092
rect 23296 22040 23348 22092
rect 31392 22108 31444 22160
rect 6368 21904 6420 21956
rect 20628 21972 20680 22024
rect 20996 22015 21048 22024
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 20996 21972 21048 21981
rect 38108 22015 38160 22024
rect 38108 21981 38117 22015
rect 38117 21981 38151 22015
rect 38151 21981 38160 22015
rect 38108 21972 38160 21981
rect 34796 21904 34848 21956
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 30288 21836 30340 21888
rect 30472 21836 30524 21888
rect 33048 21836 33100 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4620 21632 4672 21684
rect 2780 21496 2832 21548
rect 23296 21564 23348 21616
rect 23664 21496 23716 21548
rect 6552 21292 6604 21344
rect 10416 21292 10468 21344
rect 33140 21292 33192 21344
rect 34704 21292 34756 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6368 21131 6420 21140
rect 6368 21097 6377 21131
rect 6377 21097 6411 21131
rect 6411 21097 6420 21131
rect 6368 21088 6420 21097
rect 5632 20952 5684 21004
rect 6552 20995 6604 21004
rect 6552 20961 6561 20995
rect 6561 20961 6595 20995
rect 6595 20961 6604 20995
rect 6552 20952 6604 20961
rect 10232 20952 10284 21004
rect 36084 20952 36136 21004
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 37096 20884 37148 20936
rect 11060 20816 11112 20868
rect 10416 20791 10468 20800
rect 10416 20757 10425 20791
rect 10425 20757 10459 20791
rect 10459 20757 10468 20791
rect 10416 20748 10468 20757
rect 13084 20748 13136 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 7012 20544 7064 20596
rect 11060 20544 11112 20596
rect 33048 20544 33100 20596
rect 4620 20476 4672 20528
rect 29000 20476 29052 20528
rect 7472 20408 7524 20460
rect 10232 20408 10284 20460
rect 15200 20451 15252 20460
rect 6920 20340 6972 20392
rect 7380 20340 7432 20392
rect 12256 20340 12308 20392
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15844 20408 15896 20460
rect 38108 20451 38160 20460
rect 38108 20417 38117 20451
rect 38117 20417 38151 20451
rect 38151 20417 38160 20451
rect 38108 20408 38160 20417
rect 25596 20272 25648 20324
rect 28264 20315 28316 20324
rect 28264 20281 28273 20315
rect 28273 20281 28307 20315
rect 28307 20281 28316 20315
rect 28264 20272 28316 20281
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6736 20000 6788 20052
rect 10048 20000 10100 20052
rect 10416 20000 10468 20052
rect 6920 19932 6972 19984
rect 4804 19864 4856 19916
rect 7472 19932 7524 19984
rect 8208 19932 8260 19984
rect 13084 19975 13136 19984
rect 13084 19941 13093 19975
rect 13093 19941 13127 19975
rect 13127 19941 13136 19975
rect 13084 19932 13136 19941
rect 4620 19796 4672 19848
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 7380 19796 7432 19848
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 12532 19796 12584 19848
rect 17960 20000 18012 20052
rect 23664 20000 23716 20052
rect 23296 19932 23348 19984
rect 27252 19975 27304 19984
rect 27252 19941 27261 19975
rect 27261 19941 27295 19975
rect 27295 19941 27304 19975
rect 27252 19932 27304 19941
rect 19984 19864 20036 19916
rect 25596 19864 25648 19916
rect 16764 19796 16816 19848
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 23112 19796 23164 19848
rect 27160 19796 27212 19848
rect 7564 19728 7616 19780
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 12900 19703 12952 19712
rect 12900 19669 12909 19703
rect 12909 19669 12943 19703
rect 12943 19669 12952 19703
rect 12900 19660 12952 19669
rect 17684 19660 17736 19712
rect 30196 19728 30248 19780
rect 33416 19796 33468 19848
rect 22836 19660 22888 19712
rect 26240 19660 26292 19712
rect 27252 19660 27304 19712
rect 30932 19703 30984 19712
rect 30932 19669 30941 19703
rect 30941 19669 30975 19703
rect 30975 19669 30984 19703
rect 30932 19660 30984 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 12256 19499 12308 19508
rect 12256 19465 12265 19499
rect 12265 19465 12299 19499
rect 12299 19465 12308 19499
rect 12256 19456 12308 19465
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 26424 19456 26476 19508
rect 30196 19499 30248 19508
rect 30196 19465 30205 19499
rect 30205 19465 30239 19499
rect 30239 19465 30248 19499
rect 30196 19456 30248 19465
rect 33416 19499 33468 19508
rect 33416 19465 33425 19499
rect 33425 19465 33459 19499
rect 33459 19465 33468 19499
rect 33416 19456 33468 19465
rect 35992 19456 36044 19508
rect 12532 19388 12584 19440
rect 12808 19388 12860 19440
rect 19892 19431 19944 19440
rect 19892 19397 19901 19431
rect 19901 19397 19935 19431
rect 19935 19397 19944 19431
rect 19892 19388 19944 19397
rect 23664 19388 23716 19440
rect 27160 19431 27212 19440
rect 13084 19320 13136 19372
rect 17776 19320 17828 19372
rect 19800 19363 19852 19372
rect 19800 19329 19809 19363
rect 19809 19329 19843 19363
rect 19843 19329 19852 19363
rect 19800 19320 19852 19329
rect 20628 19320 20680 19372
rect 23112 19320 23164 19372
rect 27160 19397 27171 19431
rect 27171 19397 27212 19431
rect 27160 19388 27212 19397
rect 27252 19388 27304 19440
rect 26240 19363 26292 19372
rect 26240 19329 26249 19363
rect 26249 19329 26283 19363
rect 26283 19329 26292 19363
rect 26240 19320 26292 19329
rect 12900 19252 12952 19304
rect 22836 19252 22888 19304
rect 20168 19227 20220 19236
rect 20168 19193 20177 19227
rect 20177 19193 20211 19227
rect 20211 19193 20220 19227
rect 20168 19184 20220 19193
rect 12532 19116 12584 19168
rect 26240 19116 26292 19168
rect 28264 19116 28316 19168
rect 30932 19320 30984 19372
rect 34704 19388 34756 19440
rect 33416 19320 33468 19372
rect 34796 19320 34848 19372
rect 37556 19320 37608 19372
rect 38476 19252 38528 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19892 18912 19944 18964
rect 23112 18955 23164 18964
rect 23112 18921 23121 18955
rect 23121 18921 23155 18955
rect 23155 18921 23164 18955
rect 23112 18912 23164 18921
rect 25596 18912 25648 18964
rect 34704 18955 34756 18964
rect 26424 18844 26476 18896
rect 34704 18921 34713 18955
rect 34713 18921 34747 18955
rect 34747 18921 34756 18955
rect 34704 18912 34756 18921
rect 22376 18708 22428 18760
rect 22836 18708 22888 18760
rect 23296 18751 23348 18760
rect 23296 18717 23305 18751
rect 23305 18717 23339 18751
rect 23339 18717 23348 18751
rect 23296 18708 23348 18717
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 38108 18751 38160 18760
rect 38108 18717 38117 18751
rect 38117 18717 38151 18751
rect 38151 18717 38160 18751
rect 38108 18708 38160 18717
rect 19800 18683 19852 18692
rect 19800 18649 19827 18683
rect 19827 18649 19852 18683
rect 19800 18640 19852 18649
rect 19984 18683 20036 18692
rect 19984 18649 19993 18683
rect 19993 18649 20027 18683
rect 20027 18649 20036 18683
rect 19984 18640 20036 18649
rect 34428 18640 34480 18692
rect 18052 18572 18104 18624
rect 18880 18572 18932 18624
rect 23480 18615 23532 18624
rect 23480 18581 23489 18615
rect 23489 18581 23523 18615
rect 23523 18581 23532 18615
rect 23480 18572 23532 18581
rect 26056 18572 26108 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2780 18368 2832 18420
rect 17960 18368 18012 18420
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 3148 18232 3200 18241
rect 17684 18275 17736 18284
rect 17684 18241 17693 18275
rect 17693 18241 17727 18275
rect 17727 18241 17736 18275
rect 17684 18232 17736 18241
rect 18052 18232 18104 18284
rect 4804 18164 4856 18216
rect 3976 18028 4028 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3148 17824 3200 17876
rect 7380 17824 7432 17876
rect 4804 17688 4856 17740
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 7380 17620 7432 17672
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 8484 17620 8536 17672
rect 15200 17824 15252 17876
rect 22376 17867 22428 17876
rect 22376 17833 22385 17867
rect 22385 17833 22419 17867
rect 22419 17833 22428 17867
rect 22376 17824 22428 17833
rect 23480 17663 23532 17672
rect 23480 17629 23498 17663
rect 23498 17629 23532 17663
rect 23480 17620 23532 17629
rect 38108 17663 38160 17672
rect 4620 17484 4672 17536
rect 4896 17484 4948 17536
rect 12440 17484 12492 17536
rect 38108 17629 38117 17663
rect 38117 17629 38151 17663
rect 38151 17629 38160 17663
rect 38108 17620 38160 17629
rect 25780 17484 25832 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8484 17323 8536 17332
rect 8484 17289 8493 17323
rect 8493 17289 8527 17323
rect 8527 17289 8536 17323
rect 8484 17280 8536 17289
rect 26608 17280 26660 17332
rect 34336 17280 34388 17332
rect 7380 17144 7432 17196
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 17684 17212 17736 17264
rect 12440 17144 12492 17153
rect 12808 17144 12860 17196
rect 17776 17144 17828 17196
rect 33968 17144 34020 17196
rect 7012 17008 7064 17060
rect 12348 17076 12400 17128
rect 34152 17119 34204 17128
rect 12532 17008 12584 17060
rect 34152 17085 34161 17119
rect 34161 17085 34195 17119
rect 34195 17085 34204 17119
rect 34152 17076 34204 17085
rect 7288 16940 7340 16992
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4804 16736 4856 16788
rect 7012 16779 7064 16788
rect 7012 16745 7021 16779
rect 7021 16745 7055 16779
rect 7055 16745 7064 16779
rect 7012 16736 7064 16745
rect 12808 16736 12860 16788
rect 18696 16668 18748 16720
rect 17776 16600 17828 16652
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 12532 16575 12584 16584
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 17684 16575 17736 16584
rect 12532 16532 12584 16541
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 31944 16600 31996 16652
rect 31392 16575 31444 16584
rect 31392 16541 31401 16575
rect 31401 16541 31435 16575
rect 31435 16541 31444 16575
rect 31392 16532 31444 16541
rect 7196 16507 7248 16516
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 8208 16396 8260 16448
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 37740 16396 37792 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 30564 16192 30616 16244
rect 34152 16192 34204 16244
rect 34428 16235 34480 16244
rect 34428 16201 34437 16235
rect 34437 16201 34471 16235
rect 34471 16201 34480 16235
rect 34428 16192 34480 16201
rect 37832 16235 37884 16244
rect 37832 16201 37841 16235
rect 37841 16201 37875 16235
rect 37875 16201 37884 16235
rect 37832 16192 37884 16201
rect 4896 16124 4948 16176
rect 30380 16124 30432 16176
rect 6828 16056 6880 16108
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 20168 16056 20220 16108
rect 29000 16056 29052 16108
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 33416 16056 33468 16108
rect 37740 16099 37792 16108
rect 37740 16065 37749 16099
rect 37749 16065 37783 16099
rect 37783 16065 37792 16099
rect 37740 16056 37792 16065
rect 38936 16056 38988 16108
rect 31944 15988 31996 16040
rect 37924 15988 37976 16040
rect 3976 15852 4028 15904
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 33416 15895 33468 15904
rect 33416 15861 33425 15895
rect 33425 15861 33459 15895
rect 33459 15861 33468 15895
rect 33416 15852 33468 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4620 15648 4672 15700
rect 12532 15648 12584 15700
rect 20168 15648 20220 15700
rect 27252 15648 27304 15700
rect 31392 15648 31444 15700
rect 32220 15648 32272 15700
rect 34796 15691 34848 15700
rect 34796 15657 34805 15691
rect 34805 15657 34839 15691
rect 34839 15657 34848 15691
rect 34796 15648 34848 15657
rect 37924 15691 37976 15700
rect 37924 15657 37933 15691
rect 37933 15657 37967 15691
rect 37967 15657 37976 15691
rect 37924 15648 37976 15657
rect 18512 15512 18564 15564
rect 31944 15555 31996 15564
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4160 15444 4212 15496
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 6920 15308 6972 15360
rect 10048 15308 10100 15360
rect 31944 15521 31953 15555
rect 31953 15521 31987 15555
rect 31987 15521 31996 15555
rect 31944 15512 31996 15521
rect 25780 15487 25832 15496
rect 25780 15453 25789 15487
rect 25789 15453 25823 15487
rect 25823 15453 25832 15487
rect 25780 15444 25832 15453
rect 28264 15444 28316 15496
rect 29184 15444 29236 15496
rect 34704 15444 34756 15496
rect 38016 15487 38068 15496
rect 38016 15453 38025 15487
rect 38025 15453 38059 15487
rect 38059 15453 38068 15487
rect 38016 15444 38068 15453
rect 12072 15376 12124 15428
rect 18788 15376 18840 15428
rect 26056 15419 26108 15428
rect 26056 15385 26090 15419
rect 26090 15385 26108 15419
rect 26056 15376 26108 15385
rect 36452 15419 36504 15428
rect 36452 15385 36461 15419
rect 36461 15385 36495 15419
rect 36495 15385 36504 15419
rect 36452 15376 36504 15385
rect 31484 15351 31536 15360
rect 31484 15317 31493 15351
rect 31493 15317 31527 15351
rect 31527 15317 31536 15351
rect 31484 15308 31536 15317
rect 36636 15308 36688 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 7564 15104 7616 15156
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 23204 15147 23256 15156
rect 23204 15113 23213 15147
rect 23213 15113 23247 15147
rect 23247 15113 23256 15147
rect 23204 15104 23256 15113
rect 29000 15104 29052 15156
rect 30564 15104 30616 15156
rect 36544 15104 36596 15156
rect 38016 15147 38068 15156
rect 38016 15113 38025 15147
rect 38025 15113 38059 15147
rect 38059 15113 38068 15147
rect 38016 15104 38068 15113
rect 21916 15036 21968 15088
rect 29184 15079 29236 15088
rect 29184 15045 29193 15079
rect 29193 15045 29227 15079
rect 29227 15045 29236 15079
rect 29184 15036 29236 15045
rect 4068 14968 4120 15020
rect 7196 14968 7248 15020
rect 16948 14968 17000 15020
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 8300 14900 8352 14952
rect 23664 14832 23716 14884
rect 28540 14832 28592 14884
rect 29460 14875 29512 14884
rect 29460 14841 29469 14875
rect 29469 14841 29503 14875
rect 29503 14841 29512 14875
rect 29460 14832 29512 14841
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 20260 14764 20312 14816
rect 35992 14968 36044 15020
rect 37372 14968 37424 15020
rect 35992 14807 36044 14816
rect 35992 14773 36001 14807
rect 36001 14773 36035 14807
rect 36035 14773 36044 14807
rect 35992 14764 36044 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 13728 14560 13780 14612
rect 14740 14560 14792 14612
rect 6828 14424 6880 14476
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 8300 14356 8352 14408
rect 34704 14560 34756 14612
rect 15844 14424 15896 14476
rect 23204 14424 23256 14476
rect 24860 14492 24912 14544
rect 29000 14424 29052 14476
rect 36728 14424 36780 14476
rect 22468 14356 22520 14408
rect 23664 14399 23716 14408
rect 23664 14365 23673 14399
rect 23673 14365 23707 14399
rect 23707 14365 23716 14399
rect 23664 14356 23716 14365
rect 24124 14356 24176 14408
rect 29460 14356 29512 14408
rect 37280 14399 37332 14408
rect 37280 14365 37289 14399
rect 37289 14365 37323 14399
rect 37323 14365 37332 14399
rect 37280 14356 37332 14365
rect 14648 14288 14700 14340
rect 18420 14288 18472 14340
rect 31392 14288 31444 14340
rect 7196 14220 7248 14272
rect 24308 14220 24360 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 15844 14016 15896 14068
rect 16120 14016 16172 14068
rect 26332 14059 26384 14068
rect 6920 13948 6972 14000
rect 14280 13948 14332 14000
rect 15936 13948 15988 14000
rect 17960 13948 18012 14000
rect 24124 13948 24176 14000
rect 24308 13991 24360 14000
rect 24308 13957 24317 13991
rect 24317 13957 24351 13991
rect 24351 13957 24360 13991
rect 24308 13948 24360 13957
rect 25412 13948 25464 14000
rect 26332 14025 26341 14059
rect 26341 14025 26375 14059
rect 26375 14025 26384 14059
rect 26332 14016 26384 14025
rect 31392 14059 31444 14068
rect 31392 14025 31401 14059
rect 31401 14025 31435 14059
rect 31435 14025 31444 14059
rect 31392 14016 31444 14025
rect 31484 13991 31536 14000
rect 31484 13957 31493 13991
rect 31493 13957 31527 13991
rect 31527 13957 31536 13991
rect 31484 13948 31536 13957
rect 38292 13948 38344 14000
rect 3792 13880 3844 13932
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 17132 13880 17184 13932
rect 23572 13880 23624 13932
rect 37740 13923 37792 13932
rect 37740 13889 37749 13923
rect 37749 13889 37783 13923
rect 37783 13889 37792 13923
rect 37740 13880 37792 13889
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 15568 13812 15620 13864
rect 13728 13744 13780 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 22560 13472 22612 13524
rect 23572 13472 23624 13524
rect 36728 13472 36780 13524
rect 11152 13336 11204 13388
rect 10692 13268 10744 13320
rect 23664 13336 23716 13388
rect 13268 13132 13320 13184
rect 14648 13132 14700 13184
rect 22284 13243 22336 13252
rect 22284 13209 22293 13243
rect 22293 13209 22327 13243
rect 22327 13209 22336 13243
rect 22284 13200 22336 13209
rect 23204 13243 23256 13252
rect 23204 13209 23213 13243
rect 23213 13209 23247 13243
rect 23247 13209 23256 13243
rect 23204 13200 23256 13209
rect 23572 13268 23624 13320
rect 33692 13268 33744 13320
rect 31852 13200 31904 13252
rect 23112 13132 23164 13184
rect 37740 13132 37792 13184
rect 38476 13132 38528 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 20536 12928 20588 12980
rect 23480 12928 23532 12980
rect 23664 12971 23716 12980
rect 23664 12937 23673 12971
rect 23673 12937 23707 12971
rect 23707 12937 23716 12971
rect 23664 12928 23716 12937
rect 23848 12928 23900 12980
rect 13912 12860 13964 12912
rect 29000 12860 29052 12912
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7196 12835 7248 12844
rect 7196 12801 7230 12835
rect 7230 12801 7248 12835
rect 7196 12792 7248 12801
rect 13176 12792 13228 12844
rect 27528 12792 27580 12844
rect 32128 12835 32180 12844
rect 32128 12801 32137 12835
rect 32137 12801 32171 12835
rect 32171 12801 32180 12835
rect 32128 12792 32180 12801
rect 32404 12767 32456 12776
rect 32404 12733 32413 12767
rect 32413 12733 32447 12767
rect 32447 12733 32456 12767
rect 32404 12724 32456 12733
rect 9772 12656 9824 12708
rect 19800 12631 19852 12640
rect 19800 12597 19809 12631
rect 19809 12597 19843 12631
rect 19843 12597 19852 12631
rect 19800 12588 19852 12597
rect 33692 12588 33744 12640
rect 38108 12631 38160 12640
rect 38108 12597 38117 12631
rect 38117 12597 38151 12631
rect 38151 12597 38160 12631
rect 38108 12588 38160 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 20720 12384 20772 12436
rect 4620 12316 4672 12368
rect 11704 12316 11756 12368
rect 22652 12384 22704 12436
rect 7748 12248 7800 12300
rect 16304 12248 16356 12300
rect 4712 12112 4764 12164
rect 11428 12180 11480 12232
rect 14556 12044 14608 12096
rect 18236 12044 18288 12096
rect 19340 12112 19392 12164
rect 19800 12112 19852 12164
rect 23848 12112 23900 12164
rect 31392 12155 31444 12164
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 22008 12044 22060 12096
rect 28356 12044 28408 12096
rect 31392 12121 31401 12155
rect 31401 12121 31435 12155
rect 31435 12121 31444 12155
rect 31392 12112 31444 12121
rect 37924 12044 37976 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 16672 11840 16724 11892
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 19156 11840 19208 11892
rect 3056 11772 3108 11824
rect 5080 11772 5132 11824
rect 7840 11772 7892 11824
rect 22008 11772 22060 11824
rect 22192 11840 22244 11892
rect 27528 11840 27580 11892
rect 31392 11840 31444 11892
rect 24584 11772 24636 11824
rect 27988 11772 28040 11824
rect 32404 11772 32456 11824
rect 2412 11704 2464 11756
rect 3332 11704 3384 11756
rect 20444 11704 20496 11756
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 10876 11636 10928 11688
rect 9864 11568 9916 11620
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 12532 11543 12584 11552
rect 12532 11509 12541 11543
rect 12541 11509 12575 11543
rect 12575 11509 12584 11543
rect 12532 11500 12584 11509
rect 15016 11568 15068 11620
rect 19340 11636 19392 11688
rect 27068 11568 27120 11620
rect 28356 11611 28408 11620
rect 28356 11577 28365 11611
rect 28365 11577 28399 11611
rect 28399 11577 28408 11611
rect 28356 11568 28408 11577
rect 19156 11500 19208 11552
rect 28448 11500 28500 11552
rect 29000 11500 29052 11552
rect 30564 11568 30616 11620
rect 31944 11500 31996 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 15108 11296 15160 11348
rect 16304 11296 16356 11348
rect 27068 11339 27120 11348
rect 27068 11305 27077 11339
rect 27077 11305 27111 11339
rect 27111 11305 27120 11339
rect 27068 11296 27120 11305
rect 33232 11339 33284 11348
rect 33232 11305 33241 11339
rect 33241 11305 33275 11339
rect 33275 11305 33284 11339
rect 33232 11296 33284 11305
rect 37924 11339 37976 11348
rect 37924 11305 37933 11339
rect 37933 11305 37967 11339
rect 37967 11305 37976 11339
rect 37924 11296 37976 11305
rect 19340 11228 19392 11280
rect 23112 11228 23164 11280
rect 27804 11228 27856 11280
rect 2044 11092 2096 11144
rect 10876 11092 10928 11144
rect 13636 11024 13688 11076
rect 16672 11160 16724 11212
rect 25596 11160 25648 11212
rect 27988 11203 28040 11212
rect 27988 11169 27997 11203
rect 27997 11169 28031 11203
rect 28031 11169 28040 11203
rect 27988 11160 28040 11169
rect 30012 11160 30064 11212
rect 14556 11092 14608 11144
rect 20352 11092 20404 11144
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 16672 11024 16724 11076
rect 3424 10956 3476 11008
rect 19340 11024 19392 11076
rect 22284 11024 22336 11076
rect 30380 11024 30432 11076
rect 19432 10956 19484 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3240 10752 3292 10804
rect 27804 10795 27856 10804
rect 5540 10684 5592 10736
rect 27804 10761 27813 10795
rect 27813 10761 27847 10795
rect 27847 10761 27856 10795
rect 27804 10752 27856 10761
rect 24400 10684 24452 10736
rect 4988 10616 5040 10668
rect 12532 10616 12584 10668
rect 18972 10616 19024 10668
rect 3700 10548 3752 10600
rect 25964 10548 26016 10600
rect 35900 10548 35952 10600
rect 21088 10480 21140 10532
rect 12992 10412 13044 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 37280 10412 37332 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 17868 10208 17920 10260
rect 7104 10140 7156 10192
rect 17408 10140 17460 10192
rect 35808 10072 35860 10124
rect 25688 10004 25740 10056
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 2780 9936 2832 9945
rect 6184 9936 6236 9988
rect 14280 9936 14332 9988
rect 13452 9868 13504 9920
rect 17500 9868 17552 9920
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 29736 9868 29788 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 17408 9664 17460 9716
rect 4620 9596 4672 9648
rect 26884 9596 26936 9648
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 13820 9528 13872 9580
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 15936 9528 15988 9580
rect 9588 9460 9640 9512
rect 22928 9460 22980 9512
rect 24400 9503 24452 9512
rect 24400 9469 24409 9503
rect 24409 9469 24443 9503
rect 24443 9469 24452 9503
rect 24400 9460 24452 9469
rect 25136 9528 25188 9580
rect 29000 9571 29052 9580
rect 29000 9537 29009 9571
rect 29009 9537 29043 9571
rect 29043 9537 29052 9571
rect 29000 9528 29052 9537
rect 30012 9571 30064 9580
rect 30012 9537 30021 9571
rect 30021 9537 30055 9571
rect 30055 9537 30064 9571
rect 30012 9528 30064 9537
rect 37740 9571 37792 9580
rect 37740 9537 37749 9571
rect 37749 9537 37783 9571
rect 37783 9537 37792 9571
rect 37740 9528 37792 9537
rect 25044 9460 25096 9512
rect 3884 9392 3936 9444
rect 24676 9392 24728 9444
rect 25412 9392 25464 9444
rect 31024 9392 31076 9444
rect 13728 9324 13780 9376
rect 15752 9324 15804 9376
rect 32220 9324 32272 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3516 9120 3568 9172
rect 5264 9120 5316 9172
rect 5816 9120 5868 9172
rect 34060 9120 34112 9172
rect 9588 9095 9640 9104
rect 9588 9061 9597 9095
rect 9597 9061 9631 9095
rect 9631 9061 9640 9095
rect 9588 9052 9640 9061
rect 11612 9052 11664 9104
rect 20996 9095 21048 9104
rect 20996 9061 21005 9095
rect 21005 9061 21039 9095
rect 21039 9061 21048 9095
rect 20996 9052 21048 9061
rect 12624 8984 12676 9036
rect 32312 8984 32364 9036
rect 36084 8984 36136 9036
rect 3056 8848 3108 8900
rect 5356 8848 5408 8900
rect 9036 8848 9088 8900
rect 20352 8916 20404 8968
rect 23848 8916 23900 8968
rect 25044 8916 25096 8968
rect 9496 8848 9548 8900
rect 20996 8848 21048 8900
rect 25228 8848 25280 8900
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 5908 8823 5960 8832
rect 5908 8789 5917 8823
rect 5917 8789 5951 8823
rect 5951 8789 5960 8823
rect 5908 8780 5960 8789
rect 9772 8780 9824 8832
rect 20168 8780 20220 8832
rect 21180 8780 21232 8832
rect 23388 8780 23440 8832
rect 24676 8823 24728 8832
rect 24676 8789 24685 8823
rect 24685 8789 24719 8823
rect 24719 8789 24728 8823
rect 24676 8780 24728 8789
rect 35808 8916 35860 8968
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 26976 8848 27028 8900
rect 34796 8848 34848 8900
rect 26332 8780 26384 8832
rect 36452 8780 36504 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2780 8576 2832 8628
rect 4620 8576 4672 8628
rect 5908 8576 5960 8628
rect 2964 8508 3016 8560
rect 6460 8508 6512 8560
rect 3424 8440 3476 8492
rect 5356 8440 5408 8492
rect 9956 8508 10008 8560
rect 16488 8508 16540 8560
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 21180 8576 21232 8628
rect 24860 8576 24912 8628
rect 25228 8576 25280 8628
rect 34612 8576 34664 8628
rect 37832 8576 37884 8628
rect 38568 8576 38620 8628
rect 20352 8508 20404 8560
rect 30380 8508 30432 8560
rect 32312 8551 32364 8560
rect 32312 8517 32321 8551
rect 32321 8517 32355 8551
rect 32355 8517 32364 8551
rect 32312 8508 32364 8517
rect 32772 8508 32824 8560
rect 11612 8372 11664 8424
rect 3056 8304 3108 8356
rect 11796 8304 11848 8356
rect 20168 8440 20220 8492
rect 20260 8304 20312 8356
rect 25228 8440 25280 8492
rect 25596 8440 25648 8492
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 20720 8304 20772 8356
rect 23480 8347 23532 8356
rect 23480 8313 23489 8347
rect 23489 8313 23523 8347
rect 23523 8313 23532 8347
rect 23480 8304 23532 8313
rect 32312 8372 32364 8424
rect 36084 8508 36136 8560
rect 33600 8483 33652 8492
rect 33600 8449 33609 8483
rect 33609 8449 33643 8483
rect 33643 8449 33652 8483
rect 33600 8440 33652 8449
rect 37924 8372 37976 8424
rect 26332 8304 26384 8356
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 37464 8347 37516 8356
rect 37464 8313 37473 8347
rect 37473 8313 37507 8347
rect 37507 8313 37516 8347
rect 37464 8304 37516 8313
rect 11520 8236 11572 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 36912 8032 36964 8084
rect 13360 7964 13412 8016
rect 32956 7964 33008 8016
rect 31852 7896 31904 7948
rect 9680 7828 9732 7880
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 32404 7871 32456 7880
rect 32404 7837 32413 7871
rect 32413 7837 32447 7871
rect 32447 7837 32456 7871
rect 32404 7828 32456 7837
rect 38108 7871 38160 7880
rect 38108 7837 38117 7871
rect 38117 7837 38151 7871
rect 38151 7837 38160 7871
rect 38108 7828 38160 7837
rect 11428 7803 11480 7812
rect 11428 7769 11437 7803
rect 11437 7769 11471 7803
rect 11471 7769 11480 7803
rect 11428 7760 11480 7769
rect 30012 7803 30064 7812
rect 30012 7769 30021 7803
rect 30021 7769 30055 7803
rect 30055 7769 30064 7803
rect 30012 7760 30064 7769
rect 32312 7760 32364 7812
rect 35716 7760 35768 7812
rect 36728 7760 36780 7812
rect 3424 7692 3476 7744
rect 20352 7735 20404 7744
rect 20352 7701 20361 7735
rect 20361 7701 20395 7735
rect 20395 7701 20404 7735
rect 20352 7692 20404 7701
rect 25872 7692 25924 7744
rect 35348 7692 35400 7744
rect 38200 7692 38252 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 25044 7488 25096 7540
rect 28632 7531 28684 7540
rect 8116 7420 8168 7472
rect 14188 7420 14240 7472
rect 28632 7497 28641 7531
rect 28641 7497 28675 7531
rect 28675 7497 28684 7531
rect 28632 7488 28684 7497
rect 6736 7284 6788 7336
rect 11520 7395 11572 7404
rect 6644 7216 6696 7268
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 16212 7352 16264 7404
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 17224 7284 17276 7336
rect 14924 7216 14976 7268
rect 12624 7148 12676 7200
rect 16212 7148 16264 7200
rect 16488 7148 16540 7200
rect 37832 7463 37884 7472
rect 37832 7429 37841 7463
rect 37841 7429 37875 7463
rect 37875 7429 37884 7463
rect 37832 7420 37884 7429
rect 33968 7352 34020 7404
rect 35992 7352 36044 7404
rect 36544 7352 36596 7404
rect 20444 7284 20496 7336
rect 37832 7284 37884 7336
rect 20536 7216 20588 7268
rect 27620 7216 27672 7268
rect 30932 7216 30984 7268
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 27804 7148 27856 7200
rect 34612 7191 34664 7200
rect 34612 7157 34621 7191
rect 34621 7157 34655 7191
rect 34655 7157 34664 7191
rect 34612 7148 34664 7157
rect 35992 7148 36044 7200
rect 36176 7191 36228 7200
rect 36176 7157 36185 7191
rect 36185 7157 36219 7191
rect 36219 7157 36228 7191
rect 36176 7148 36228 7157
rect 38108 7148 38160 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 14924 6987 14976 6996
rect 14924 6953 14933 6987
rect 14933 6953 14967 6987
rect 14967 6953 14976 6987
rect 14924 6944 14976 6953
rect 17224 6944 17276 6996
rect 28908 6944 28960 6996
rect 6644 6808 6696 6860
rect 16028 6851 16080 6860
rect 16028 6817 16037 6851
rect 16037 6817 16071 6851
rect 16071 6817 16080 6851
rect 20536 6876 20588 6928
rect 23204 6876 23256 6928
rect 30932 6876 30984 6928
rect 16028 6808 16080 6817
rect 20812 6740 20864 6792
rect 24952 6808 25004 6860
rect 16488 6672 16540 6724
rect 19984 6715 20036 6724
rect 19984 6681 19993 6715
rect 19993 6681 20027 6715
rect 20027 6681 20036 6715
rect 19984 6672 20036 6681
rect 24860 6715 24912 6724
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 19432 6604 19484 6656
rect 20444 6604 20496 6656
rect 20628 6604 20680 6656
rect 24860 6681 24869 6715
rect 24869 6681 24903 6715
rect 24903 6681 24912 6715
rect 24860 6672 24912 6681
rect 25044 6672 25096 6724
rect 28724 6808 28776 6860
rect 32312 6808 32364 6860
rect 35624 6740 35676 6792
rect 30012 6672 30064 6724
rect 34520 6672 34572 6724
rect 35348 6672 35400 6724
rect 37280 6740 37332 6792
rect 39580 6672 39632 6724
rect 28632 6604 28684 6656
rect 29920 6647 29972 6656
rect 29920 6613 29929 6647
rect 29929 6613 29963 6647
rect 29963 6613 29972 6647
rect 29920 6604 29972 6613
rect 30380 6604 30432 6656
rect 32312 6604 32364 6656
rect 32588 6647 32640 6656
rect 32588 6613 32597 6647
rect 32597 6613 32631 6647
rect 32631 6613 32640 6647
rect 32588 6604 32640 6613
rect 33876 6604 33928 6656
rect 35808 6604 35860 6656
rect 37372 6647 37424 6656
rect 37372 6613 37381 6647
rect 37381 6613 37415 6647
rect 37415 6613 37424 6647
rect 37372 6604 37424 6613
rect 38476 6604 38528 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 5172 6400 5224 6452
rect 15568 6443 15620 6452
rect 15568 6409 15577 6443
rect 15577 6409 15611 6443
rect 15611 6409 15620 6443
rect 15568 6400 15620 6409
rect 35900 6400 35952 6452
rect 37740 6400 37792 6452
rect 16580 6332 16632 6384
rect 35992 6332 36044 6384
rect 2780 6196 2832 6248
rect 15844 6264 15896 6316
rect 16488 6264 16540 6316
rect 17684 6264 17736 6316
rect 35256 6307 35308 6316
rect 35256 6273 35265 6307
rect 35265 6273 35299 6307
rect 35299 6273 35308 6307
rect 35256 6264 35308 6273
rect 35900 6264 35952 6316
rect 37372 6332 37424 6384
rect 38752 6332 38804 6384
rect 39028 6264 39080 6316
rect 25688 6196 25740 6248
rect 31852 6196 31904 6248
rect 30012 6128 30064 6180
rect 34520 6128 34572 6180
rect 1584 6060 1636 6112
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 15108 6103 15160 6112
rect 15108 6069 15117 6103
rect 15117 6069 15151 6103
rect 15151 6069 15160 6103
rect 15108 6060 15160 6069
rect 17684 6060 17736 6112
rect 29644 6103 29696 6112
rect 29644 6069 29653 6103
rect 29653 6069 29687 6103
rect 29687 6069 29696 6103
rect 29644 6060 29696 6069
rect 30472 6103 30524 6112
rect 30472 6069 30481 6103
rect 30481 6069 30515 6103
rect 30515 6069 30524 6103
rect 30472 6060 30524 6069
rect 30932 6103 30984 6112
rect 30932 6069 30941 6103
rect 30941 6069 30975 6103
rect 30975 6069 30984 6103
rect 30932 6060 30984 6069
rect 31760 6060 31812 6112
rect 32956 6103 33008 6112
rect 32956 6069 32965 6103
rect 32965 6069 32999 6103
rect 32999 6069 33008 6103
rect 32956 6060 33008 6069
rect 34060 6060 34112 6112
rect 37740 6103 37792 6112
rect 37740 6069 37749 6103
rect 37749 6069 37783 6103
rect 37783 6069 37792 6103
rect 37740 6060 37792 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4712 5856 4764 5908
rect 16120 5899 16172 5908
rect 16120 5865 16129 5899
rect 16129 5865 16163 5899
rect 16163 5865 16172 5899
rect 16120 5856 16172 5865
rect 18420 5856 18472 5908
rect 30656 5899 30708 5908
rect 30656 5865 30665 5899
rect 30665 5865 30699 5899
rect 30699 5865 30708 5899
rect 30656 5856 30708 5865
rect 31208 5899 31260 5908
rect 31208 5865 31217 5899
rect 31217 5865 31251 5899
rect 31251 5865 31260 5899
rect 31208 5856 31260 5865
rect 32680 5856 32732 5908
rect 33968 5899 34020 5908
rect 33968 5865 33977 5899
rect 33977 5865 34011 5899
rect 34011 5865 34020 5899
rect 33968 5856 34020 5865
rect 34796 5856 34848 5908
rect 39304 5856 39356 5908
rect 24032 5788 24084 5840
rect 37740 5788 37792 5840
rect 13820 5720 13872 5772
rect 22284 5720 22336 5772
rect 36084 5720 36136 5772
rect 6644 5652 6696 5704
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 30656 5652 30708 5704
rect 1768 5584 1820 5636
rect 2780 5584 2832 5636
rect 4712 5627 4764 5636
rect 4712 5593 4721 5627
rect 4721 5593 4755 5627
rect 4755 5593 4764 5627
rect 4712 5584 4764 5593
rect 1400 5559 1452 5568
rect 1400 5525 1409 5559
rect 1409 5525 1443 5559
rect 1443 5525 1452 5559
rect 1400 5516 1452 5525
rect 1676 5516 1728 5568
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 5080 5516 5132 5568
rect 5632 5516 5684 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 8024 5559 8076 5568
rect 6920 5516 6972 5525
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 11152 5516 11204 5568
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 24860 5584 24912 5636
rect 34060 5652 34112 5704
rect 35624 5652 35676 5704
rect 36636 5695 36688 5704
rect 36636 5661 36645 5695
rect 36645 5661 36679 5695
rect 36679 5661 36688 5695
rect 36636 5652 36688 5661
rect 37096 5695 37148 5704
rect 37096 5661 37105 5695
rect 37105 5661 37139 5695
rect 37139 5661 37148 5695
rect 37096 5652 37148 5661
rect 35808 5584 35860 5636
rect 38016 5627 38068 5636
rect 38016 5593 38025 5627
rect 38025 5593 38059 5627
rect 38059 5593 38068 5627
rect 38016 5584 38068 5593
rect 14188 5559 14240 5568
rect 14188 5525 14197 5559
rect 14197 5525 14231 5559
rect 14231 5525 14240 5559
rect 14188 5516 14240 5525
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 15660 5559 15712 5568
rect 15660 5525 15669 5559
rect 15669 5525 15703 5559
rect 15703 5525 15712 5559
rect 15660 5516 15712 5525
rect 20076 5516 20128 5568
rect 20904 5516 20956 5568
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 24492 5559 24544 5568
rect 24492 5525 24501 5559
rect 24501 5525 24535 5559
rect 24535 5525 24544 5559
rect 24492 5516 24544 5525
rect 25228 5559 25280 5568
rect 25228 5525 25237 5559
rect 25237 5525 25271 5559
rect 25271 5525 25280 5559
rect 25228 5516 25280 5525
rect 25412 5516 25464 5568
rect 26424 5516 26476 5568
rect 26516 5516 26568 5568
rect 26884 5559 26936 5568
rect 26884 5525 26893 5559
rect 26893 5525 26927 5559
rect 26927 5525 26936 5559
rect 26884 5516 26936 5525
rect 29092 5516 29144 5568
rect 31300 5516 31352 5568
rect 33232 5516 33284 5568
rect 36084 5516 36136 5568
rect 37740 5516 37792 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 26056 5312 26108 5364
rect 26608 5312 26660 5364
rect 29276 5355 29328 5364
rect 29276 5321 29285 5355
rect 29285 5321 29319 5355
rect 29319 5321 29328 5355
rect 29276 5312 29328 5321
rect 31944 5312 31996 5364
rect 32404 5312 32456 5364
rect 33600 5312 33652 5364
rect 34888 5355 34940 5364
rect 34888 5321 34897 5355
rect 34897 5321 34931 5355
rect 34931 5321 34940 5355
rect 34888 5312 34940 5321
rect 35532 5355 35584 5364
rect 35532 5321 35541 5355
rect 35541 5321 35575 5355
rect 35575 5321 35584 5355
rect 35532 5312 35584 5321
rect 37372 5355 37424 5364
rect 37372 5321 37381 5355
rect 37381 5321 37415 5355
rect 37415 5321 37424 5355
rect 37372 5312 37424 5321
rect 12256 5244 12308 5296
rect 13268 5244 13320 5296
rect 31300 5244 31352 5296
rect 30656 5176 30708 5228
rect 31208 5176 31260 5228
rect 32864 5244 32916 5296
rect 32956 5176 33008 5228
rect 33876 5176 33928 5228
rect 34244 5176 34296 5228
rect 36452 5219 36504 5228
rect 36452 5185 36461 5219
rect 36461 5185 36495 5219
rect 36495 5185 36504 5219
rect 36452 5176 36504 5185
rect 38108 5219 38160 5228
rect 38108 5185 38117 5219
rect 38117 5185 38151 5219
rect 38151 5185 38160 5219
rect 38108 5176 38160 5185
rect 11704 5108 11756 5160
rect 27436 5108 27488 5160
rect 4712 5040 4764 5092
rect 16396 5040 16448 5092
rect 27620 5040 27672 5092
rect 32036 5040 32088 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 2964 4972 3016 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 4620 4972 4672 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 7748 4972 7800 5024
rect 8208 4972 8260 5024
rect 8576 4972 8628 5024
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 11244 4972 11296 5024
rect 12532 4972 12584 5024
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 14096 4972 14148 5024
rect 14832 5015 14884 5024
rect 14832 4981 14841 5015
rect 14841 4981 14875 5015
rect 14875 4981 14884 5015
rect 14832 4972 14884 4981
rect 15752 5015 15804 5024
rect 15752 4981 15761 5015
rect 15761 4981 15795 5015
rect 15795 4981 15804 5015
rect 15752 4972 15804 4981
rect 16488 4972 16540 5024
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 18972 5015 19024 5024
rect 18972 4981 18981 5015
rect 18981 4981 19015 5015
rect 19015 4981 19024 5015
rect 18972 4972 19024 4981
rect 19156 4972 19208 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 21180 4972 21232 5024
rect 21456 4972 21508 5024
rect 22376 5015 22428 5024
rect 22376 4981 22385 5015
rect 22385 4981 22419 5015
rect 22419 4981 22428 5015
rect 22376 4972 22428 4981
rect 22560 4972 22612 5024
rect 24216 4972 24268 5024
rect 24400 4972 24452 5024
rect 25044 5015 25096 5024
rect 25044 4981 25053 5015
rect 25053 4981 25087 5015
rect 25087 4981 25096 5015
rect 25044 4972 25096 4981
rect 26700 4972 26752 5024
rect 27528 5015 27580 5024
rect 27528 4981 27537 5015
rect 27537 4981 27571 5015
rect 27571 4981 27580 5015
rect 27528 4972 27580 4981
rect 27988 5015 28040 5024
rect 27988 4981 27997 5015
rect 27997 4981 28031 5015
rect 28031 4981 28040 5015
rect 27988 4972 28040 4981
rect 28080 4972 28132 5024
rect 31944 4972 31996 5024
rect 36820 4972 36872 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 5172 4768 5224 4820
rect 2872 4700 2924 4752
rect 8484 4700 8536 4752
rect 12256 4743 12308 4752
rect 12256 4709 12265 4743
rect 12265 4709 12299 4743
rect 12299 4709 12308 4743
rect 12256 4700 12308 4709
rect 12716 4768 12768 4820
rect 25136 4811 25188 4820
rect 25136 4777 25145 4811
rect 25145 4777 25179 4811
rect 25179 4777 25188 4811
rect 25136 4768 25188 4777
rect 30564 4811 30616 4820
rect 19340 4700 19392 4752
rect 22192 4700 22244 4752
rect 1584 4564 1636 4616
rect 1768 4564 1820 4616
rect 2504 4564 2556 4616
rect 8300 4632 8352 4684
rect 5264 4564 5316 4616
rect 6920 4564 6972 4616
rect 7932 4564 7984 4616
rect 7748 4496 7800 4548
rect 9036 4539 9088 4548
rect 9036 4505 9045 4539
rect 9045 4505 9079 4539
rect 9079 4505 9088 4539
rect 9036 4496 9088 4505
rect 11152 4564 11204 4616
rect 12716 4564 12768 4616
rect 13360 4564 13412 4616
rect 13452 4564 13504 4616
rect 14188 4564 14240 4616
rect 16396 4564 16448 4616
rect 22468 4632 22520 4684
rect 25964 4675 26016 4684
rect 25964 4641 25973 4675
rect 25973 4641 26007 4675
rect 26007 4641 26016 4675
rect 25964 4632 26016 4641
rect 20076 4607 20128 4616
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 4160 4428 4212 4480
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 6552 4471 6604 4480
rect 6552 4437 6561 4471
rect 6561 4437 6595 4471
rect 6595 4437 6604 4471
rect 6552 4428 6604 4437
rect 8116 4428 8168 4480
rect 9956 4428 10008 4480
rect 17500 4496 17552 4548
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 21456 4564 21508 4616
rect 21732 4564 21784 4616
rect 22100 4564 22152 4616
rect 25044 4564 25096 4616
rect 26332 4564 26384 4616
rect 27252 4700 27304 4752
rect 30564 4777 30573 4811
rect 30573 4777 30607 4811
rect 30607 4777 30616 4811
rect 30564 4768 30616 4777
rect 33508 4768 33560 4820
rect 31852 4700 31904 4752
rect 33600 4700 33652 4752
rect 35440 4700 35492 4752
rect 27068 4632 27120 4684
rect 27620 4564 27672 4616
rect 30380 4607 30432 4616
rect 30380 4573 30389 4607
rect 30389 4573 30423 4607
rect 30423 4573 30432 4607
rect 30380 4564 30432 4573
rect 31024 4607 31076 4616
rect 31024 4573 31033 4607
rect 31033 4573 31067 4607
rect 31067 4573 31076 4607
rect 31024 4564 31076 4573
rect 20996 4496 21048 4548
rect 12348 4428 12400 4480
rect 13912 4428 13964 4480
rect 14464 4428 14516 4480
rect 15476 4428 15528 4480
rect 16212 4428 16264 4480
rect 17592 4471 17644 4480
rect 17592 4437 17601 4471
rect 17601 4437 17635 4471
rect 17635 4437 17644 4471
rect 17592 4428 17644 4437
rect 18052 4428 18104 4480
rect 20168 4428 20220 4480
rect 20536 4428 20588 4480
rect 26792 4496 26844 4548
rect 27160 4496 27212 4548
rect 28724 4496 28776 4548
rect 33968 4607 34020 4616
rect 33968 4573 33977 4607
rect 33977 4573 34011 4607
rect 34011 4573 34020 4607
rect 33968 4564 34020 4573
rect 36084 4607 36136 4616
rect 36084 4573 36093 4607
rect 36093 4573 36127 4607
rect 36127 4573 36136 4607
rect 36084 4564 36136 4573
rect 37096 4564 37148 4616
rect 33508 4496 33560 4548
rect 37188 4539 37240 4548
rect 37188 4505 37197 4539
rect 37197 4505 37231 4539
rect 37231 4505 37240 4539
rect 37188 4496 37240 4505
rect 37280 4496 37332 4548
rect 37924 4496 37976 4548
rect 22744 4428 22796 4480
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 26332 4428 26384 4480
rect 27436 4471 27488 4480
rect 27436 4437 27445 4471
rect 27445 4437 27479 4471
rect 27479 4437 27488 4471
rect 27436 4428 27488 4437
rect 29828 4428 29880 4480
rect 30196 4428 30248 4480
rect 34152 4471 34204 4480
rect 34152 4437 34161 4471
rect 34161 4437 34195 4471
rect 34195 4437 34204 4471
rect 34152 4428 34204 4437
rect 35992 4428 36044 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3884 4224 3936 4276
rect 8484 4224 8536 4276
rect 12256 4224 12308 4276
rect 572 4088 624 4140
rect 1952 4088 2004 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3240 4088 3292 4140
rect 5080 4156 5132 4208
rect 296 4020 348 4072
rect 1584 4020 1636 4072
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 4804 4088 4856 4140
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 5632 4156 5684 4208
rect 7196 4156 7248 4208
rect 8116 4156 8168 4208
rect 20536 4267 20588 4276
rect 20536 4233 20545 4267
rect 20545 4233 20579 4267
rect 20579 4233 20588 4267
rect 20536 4224 20588 4233
rect 20996 4224 21048 4276
rect 21916 4224 21968 4276
rect 24584 4224 24636 4276
rect 25964 4224 26016 4276
rect 27620 4267 27672 4276
rect 4896 4088 4948 4097
rect 5448 4088 5500 4140
rect 6368 4088 6420 4140
rect 11336 4088 11388 4140
rect 11704 4088 11756 4140
rect 11980 4088 12032 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 2412 3995 2464 4004
rect 2412 3961 2421 3995
rect 2421 3961 2455 3995
rect 2455 3961 2464 3995
rect 2412 3952 2464 3961
rect 3608 3952 3660 4004
rect 7564 4020 7616 4072
rect 8484 4020 8536 4072
rect 8576 4020 8628 4072
rect 9680 4020 9732 4072
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 12256 4020 12308 4072
rect 16120 4088 16172 4140
rect 19340 4131 19392 4140
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 27068 4156 27120 4208
rect 27620 4233 27629 4267
rect 27629 4233 27663 4267
rect 27663 4233 27672 4267
rect 27620 4224 27672 4233
rect 28264 4224 28316 4276
rect 22284 4088 22336 4140
rect 23020 4088 23072 4140
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 24032 4131 24084 4140
rect 24032 4097 24041 4131
rect 24041 4097 24075 4131
rect 24075 4097 24084 4131
rect 24032 4088 24084 4097
rect 2780 3884 2832 3936
rect 5632 3952 5684 4004
rect 7932 3952 7984 4004
rect 10600 3995 10652 4004
rect 10600 3961 10609 3995
rect 10609 3961 10643 3995
rect 10643 3961 10652 3995
rect 10600 3952 10652 3961
rect 11428 3952 11480 4004
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 5356 3884 5408 3936
rect 5540 3884 5592 3936
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 10968 3884 11020 3936
rect 12992 3952 13044 4004
rect 15568 4020 15620 4072
rect 19064 4063 19116 4072
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 19892 4020 19944 4072
rect 20444 4063 20496 4072
rect 20444 4029 20453 4063
rect 20453 4029 20487 4063
rect 20487 4029 20496 4063
rect 20444 4020 20496 4029
rect 15844 3952 15896 4004
rect 17316 3952 17368 4004
rect 12164 3884 12216 3936
rect 13728 3884 13780 3936
rect 14740 3884 14792 3936
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17040 3884 17092 3936
rect 18144 3884 18196 3936
rect 20812 3952 20864 4004
rect 22652 4020 22704 4072
rect 24584 4020 24636 4072
rect 25320 4020 25372 4072
rect 20996 3952 21048 4004
rect 26056 3995 26108 4004
rect 26056 3961 26065 3995
rect 26065 3961 26099 3995
rect 26099 3961 26108 3995
rect 26056 3952 26108 3961
rect 26976 3995 27028 4004
rect 26976 3961 26985 3995
rect 26985 3961 27019 3995
rect 27019 3961 27028 3995
rect 26976 3952 27028 3961
rect 22008 3884 22060 3936
rect 22836 3884 22888 3936
rect 23664 3884 23716 3936
rect 25780 3884 25832 3936
rect 27528 4088 27580 4140
rect 28632 4131 28684 4140
rect 28632 4097 28641 4131
rect 28641 4097 28675 4131
rect 28675 4097 28684 4131
rect 28632 4088 28684 4097
rect 29368 4088 29420 4140
rect 30380 4224 30432 4276
rect 31484 4224 31536 4276
rect 31668 4224 31720 4276
rect 34244 4224 34296 4276
rect 29828 4063 29880 4072
rect 29828 4029 29837 4063
rect 29837 4029 29871 4063
rect 29871 4029 29880 4063
rect 29828 4020 29880 4029
rect 30932 4156 30984 4208
rect 30748 4088 30800 4140
rect 32220 4088 32272 4140
rect 32312 4088 32364 4140
rect 33968 4131 34020 4140
rect 28540 3884 28592 3936
rect 29000 3884 29052 3936
rect 29552 3952 29604 4004
rect 32220 3952 32272 4004
rect 33968 4097 33977 4131
rect 33977 4097 34011 4131
rect 34011 4097 34020 4131
rect 33968 4088 34020 4097
rect 33140 4020 33192 4072
rect 36268 4156 36320 4208
rect 34152 4088 34204 4140
rect 37280 4131 37332 4140
rect 37280 4097 37289 4131
rect 37289 4097 37323 4131
rect 37323 4097 37332 4131
rect 37280 4088 37332 4097
rect 38384 4088 38436 4140
rect 30656 3884 30708 3936
rect 31852 3884 31904 3936
rect 33784 3884 33836 3936
rect 38660 3952 38712 4004
rect 34428 3884 34480 3936
rect 34796 3884 34848 3936
rect 35348 3884 35400 3936
rect 36452 3927 36504 3936
rect 36452 3893 36461 3927
rect 36461 3893 36495 3927
rect 36495 3893 36504 3927
rect 36452 3884 36504 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 6184 3723 6236 3732
rect 6184 3689 6193 3723
rect 6193 3689 6227 3723
rect 6227 3689 6236 3723
rect 6184 3680 6236 3689
rect 7564 3680 7616 3732
rect 11520 3723 11572 3732
rect 1952 3612 2004 3664
rect 3148 3612 3200 3664
rect 848 3544 900 3596
rect 2964 3544 3016 3596
rect 1676 3476 1728 3528
rect 5172 3544 5224 3596
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 8300 3612 8352 3664
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 13176 3723 13228 3732
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 14004 3680 14056 3732
rect 16948 3723 17000 3732
rect 16948 3689 16957 3723
rect 16957 3689 16991 3723
rect 16991 3689 17000 3723
rect 16948 3680 17000 3689
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 19892 3680 19944 3732
rect 20536 3680 20588 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 23388 3680 23440 3732
rect 23940 3680 23992 3732
rect 24032 3680 24084 3732
rect 36452 3680 36504 3732
rect 5540 3544 5592 3553
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 8392 3544 8444 3596
rect 2964 3340 3016 3392
rect 4436 3476 4488 3528
rect 4528 3451 4580 3460
rect 4528 3417 4537 3451
rect 4537 3417 4571 3451
rect 4571 3417 4580 3451
rect 4528 3408 4580 3417
rect 6092 3408 6144 3460
rect 7472 3476 7524 3528
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 9404 3476 9456 3528
rect 9864 3544 9916 3596
rect 10784 3544 10836 3596
rect 6828 3408 6880 3460
rect 9864 3408 9916 3460
rect 10876 3408 10928 3460
rect 12348 3476 12400 3528
rect 12532 3587 12584 3596
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 14188 3544 14240 3596
rect 15844 3587 15896 3596
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 17132 3612 17184 3664
rect 16304 3544 16356 3596
rect 26240 3612 26292 3664
rect 17500 3587 17552 3596
rect 17500 3553 17509 3587
rect 17509 3553 17543 3587
rect 17543 3553 17552 3587
rect 21916 3587 21968 3596
rect 17500 3544 17552 3553
rect 21916 3553 21925 3587
rect 21925 3553 21959 3587
rect 21959 3553 21968 3587
rect 21916 3544 21968 3553
rect 22100 3587 22152 3596
rect 22100 3553 22109 3587
rect 22109 3553 22143 3587
rect 22143 3553 22152 3587
rect 22100 3544 22152 3553
rect 23020 3544 23072 3596
rect 28356 3612 28408 3664
rect 26424 3544 26476 3596
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 18972 3476 19024 3528
rect 19248 3476 19300 3528
rect 20352 3476 20404 3528
rect 20628 3476 20680 3528
rect 21180 3519 21232 3528
rect 21180 3485 21189 3519
rect 21189 3485 21223 3519
rect 21223 3485 21232 3519
rect 21180 3476 21232 3485
rect 22192 3519 22244 3528
rect 22192 3485 22201 3519
rect 22201 3485 22235 3519
rect 22235 3485 22244 3519
rect 22192 3476 22244 3485
rect 22744 3476 22796 3528
rect 7656 3340 7708 3392
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 11428 3408 11480 3460
rect 14464 3451 14516 3460
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 14464 3417 14473 3451
rect 14473 3417 14507 3451
rect 14507 3417 14516 3451
rect 14464 3408 14516 3417
rect 25320 3476 25372 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 29828 3612 29880 3664
rect 31576 3655 31628 3664
rect 31576 3621 31585 3655
rect 31585 3621 31619 3655
rect 31619 3621 31628 3655
rect 31576 3612 31628 3621
rect 30288 3587 30340 3596
rect 12808 3340 12860 3349
rect 17868 3340 17920 3392
rect 24216 3408 24268 3460
rect 24768 3451 24820 3460
rect 24768 3417 24777 3451
rect 24777 3417 24811 3451
rect 24811 3417 24820 3451
rect 24768 3408 24820 3417
rect 26792 3408 26844 3460
rect 23296 3383 23348 3392
rect 23296 3349 23305 3383
rect 23305 3349 23339 3383
rect 23339 3349 23348 3383
rect 23296 3340 23348 3349
rect 25596 3383 25648 3392
rect 25596 3349 25605 3383
rect 25605 3349 25639 3383
rect 25639 3349 25648 3383
rect 25596 3340 25648 3349
rect 26056 3340 26108 3392
rect 26884 3340 26936 3392
rect 27712 3340 27764 3392
rect 28172 3340 28224 3392
rect 29920 3476 29972 3528
rect 30288 3553 30297 3587
rect 30297 3553 30331 3587
rect 30331 3553 30340 3587
rect 30288 3544 30340 3553
rect 34152 3612 34204 3664
rect 37280 3544 37332 3596
rect 37648 3544 37700 3596
rect 38200 3544 38252 3596
rect 30748 3476 30800 3528
rect 31760 3476 31812 3528
rect 32036 3519 32088 3528
rect 32036 3485 32045 3519
rect 32045 3485 32079 3519
rect 32079 3485 32088 3519
rect 32036 3476 32088 3485
rect 31668 3408 31720 3460
rect 31944 3408 31996 3460
rect 33692 3476 33744 3528
rect 34796 3476 34848 3528
rect 35440 3476 35492 3528
rect 38384 3476 38436 3528
rect 34520 3408 34572 3460
rect 35164 3408 35216 3460
rect 38936 3408 38988 3460
rect 31024 3340 31076 3392
rect 32680 3340 32732 3392
rect 34336 3340 34388 3392
rect 34428 3340 34480 3392
rect 38568 3340 38620 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3332 3136 3384 3188
rect 4528 3136 4580 3188
rect 5540 3136 5592 3188
rect 8208 3136 8260 3188
rect 9496 3136 9548 3188
rect 13636 3136 13688 3188
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17684 3136 17736 3188
rect 18604 3179 18656 3188
rect 4160 3111 4212 3120
rect 4160 3077 4169 3111
rect 4169 3077 4203 3111
rect 4203 3077 4212 3111
rect 4160 3068 4212 3077
rect 4896 3111 4948 3120
rect 4896 3077 4905 3111
rect 4905 3077 4939 3111
rect 4939 3077 4948 3111
rect 4896 3068 4948 3077
rect 5080 3068 5132 3120
rect 11428 3068 11480 3120
rect 1124 3000 1176 3052
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 3332 3000 3384 3052
rect 3700 3000 3752 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5816 3000 5868 3052
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 3884 2932 3936 2984
rect 6552 3000 6604 3052
rect 8024 3000 8076 3052
rect 4436 2864 4488 2916
rect 4712 2864 4764 2916
rect 5448 2864 5500 2916
rect 9220 2932 9272 2984
rect 10140 3000 10192 3052
rect 10600 3000 10652 3052
rect 11612 3000 11664 3052
rect 11796 3000 11848 3052
rect 9864 2932 9916 2984
rect 9956 2932 10008 2984
rect 12624 3000 12676 3052
rect 13268 3068 13320 3120
rect 15752 3068 15804 3120
rect 17960 3111 18012 3120
rect 13912 3043 13964 3052
rect 5632 2864 5684 2916
rect 10784 2864 10836 2916
rect 11336 2864 11388 2916
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14648 3000 14700 3052
rect 15108 3000 15160 3052
rect 17960 3077 17969 3111
rect 17969 3077 18003 3111
rect 18003 3077 18012 3111
rect 17960 3068 18012 3077
rect 18604 3145 18613 3179
rect 18613 3145 18647 3179
rect 18647 3145 18656 3179
rect 18604 3136 18656 3145
rect 19984 3136 20036 3188
rect 24032 3136 24084 3188
rect 35164 3136 35216 3188
rect 36360 3136 36412 3188
rect 15936 2932 15988 2984
rect 17224 3000 17276 3052
rect 17684 3000 17736 3052
rect 18052 3000 18104 3052
rect 18328 3000 18380 3052
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 16764 2932 16816 2984
rect 18972 2932 19024 2984
rect 20168 3000 20220 3052
rect 20996 3043 21048 3052
rect 20996 3009 21005 3043
rect 21005 3009 21039 3043
rect 21039 3009 21048 3043
rect 20996 3000 21048 3009
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 28172 3068 28224 3120
rect 28356 3111 28408 3120
rect 28356 3077 28365 3111
rect 28365 3077 28399 3111
rect 28399 3077 28408 3111
rect 28356 3068 28408 3077
rect 28816 3111 28868 3120
rect 28816 3077 28825 3111
rect 28825 3077 28859 3111
rect 28859 3077 28868 3111
rect 28816 3068 28868 3077
rect 28908 3068 28960 3120
rect 23112 3000 23164 3052
rect 23756 3000 23808 3052
rect 19984 2932 20036 2984
rect 20352 2932 20404 2984
rect 22560 2932 22612 2984
rect 23388 2932 23440 2984
rect 24492 3000 24544 3052
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 25872 3000 25924 3052
rect 27436 3000 27488 3052
rect 27988 3000 28040 3052
rect 28080 3000 28132 3052
rect 18236 2864 18288 2916
rect 24492 2864 24544 2916
rect 112 2796 164 2848
rect 1400 2796 1452 2848
rect 5540 2796 5592 2848
rect 7564 2839 7616 2848
rect 7564 2805 7573 2839
rect 7573 2805 7607 2839
rect 7607 2805 7616 2839
rect 7564 2796 7616 2805
rect 8852 2796 8904 2848
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 18696 2796 18748 2848
rect 20352 2796 20404 2848
rect 21180 2796 21232 2848
rect 25320 2796 25372 2848
rect 26424 2864 26476 2916
rect 27528 2907 27580 2916
rect 25780 2796 25832 2848
rect 27528 2873 27537 2907
rect 27537 2873 27571 2907
rect 27571 2873 27580 2907
rect 27528 2864 27580 2873
rect 28908 2932 28960 2984
rect 29092 2932 29144 2984
rect 30472 3000 30524 3052
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 34428 3068 34480 3120
rect 34888 3111 34940 3120
rect 34888 3077 34897 3111
rect 34897 3077 34931 3111
rect 34931 3077 34940 3111
rect 34888 3068 34940 3077
rect 35440 3068 35492 3120
rect 35716 3111 35768 3120
rect 35716 3077 35725 3111
rect 35725 3077 35759 3111
rect 35759 3077 35768 3111
rect 35716 3068 35768 3077
rect 32404 3000 32456 3052
rect 32588 3000 32640 3052
rect 33784 3043 33836 3052
rect 33784 3009 33793 3043
rect 33793 3009 33827 3043
rect 33827 3009 33836 3043
rect 33784 3000 33836 3009
rect 32128 2932 32180 2984
rect 38292 3068 38344 3120
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 37464 3000 37516 3052
rect 37372 2932 37424 2984
rect 38752 2864 38804 2916
rect 33508 2796 33560 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 9680 2592 9732 2644
rect 21916 2635 21968 2644
rect 10048 2524 10100 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 3056 2456 3108 2508
rect 4436 2456 4488 2508
rect 4620 2456 4672 2508
rect 9036 2456 9088 2508
rect 9128 2456 9180 2508
rect 9588 2456 9640 2508
rect 2228 2388 2280 2440
rect 2596 2388 2648 2440
rect 2872 2388 2924 2440
rect 4068 2388 4120 2440
rect 4988 2388 5040 2440
rect 6460 2388 6512 2440
rect 1400 2320 1452 2372
rect 1768 2320 1820 2372
rect 4160 2320 4212 2372
rect 4804 2320 4856 2372
rect 6092 2320 6144 2372
rect 8116 2388 8168 2440
rect 14924 2524 14976 2576
rect 18788 2524 18840 2576
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 23572 2592 23624 2644
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 10324 2456 10376 2508
rect 10232 2388 10284 2440
rect 10692 2388 10744 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 14464 2456 14516 2508
rect 31392 2592 31444 2644
rect 25780 2524 25832 2576
rect 34704 2592 34756 2644
rect 36452 2524 36504 2576
rect 10784 2388 10836 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14832 2388 14884 2440
rect 15660 2388 15712 2440
rect 16488 2388 16540 2440
rect 17316 2388 17368 2440
rect 17592 2388 17644 2440
rect 20260 2388 20312 2440
rect 22284 2388 22336 2440
rect 24400 2431 24452 2440
rect 8300 2320 8352 2372
rect 11244 2320 11296 2372
rect 12532 2320 12584 2372
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 13820 2320 13872 2372
rect 18144 2320 18196 2372
rect 18420 2320 18472 2372
rect 19156 2320 19208 2372
rect 20628 2320 20680 2372
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 27252 2388 27304 2440
rect 28080 2431 28132 2440
rect 28080 2397 28089 2431
rect 28089 2397 28123 2431
rect 28123 2397 28132 2431
rect 28080 2388 28132 2397
rect 29000 2431 29052 2440
rect 29000 2397 29009 2431
rect 29009 2397 29043 2431
rect 29043 2397 29052 2431
rect 29000 2388 29052 2397
rect 29644 2388 29696 2440
rect 30104 2456 30156 2508
rect 32220 2499 32272 2508
rect 32220 2465 32229 2499
rect 32229 2465 32263 2499
rect 32263 2465 32272 2499
rect 32220 2456 32272 2465
rect 32496 2499 32548 2508
rect 32496 2465 32505 2499
rect 32505 2465 32539 2499
rect 32539 2465 32548 2499
rect 32496 2456 32548 2465
rect 36084 2456 36136 2508
rect 36544 2456 36596 2508
rect 37556 2499 37608 2508
rect 37556 2465 37565 2499
rect 37565 2465 37599 2499
rect 37599 2465 37608 2499
rect 37556 2456 37608 2465
rect 24768 2320 24820 2372
rect 24860 2320 24912 2372
rect 26700 2320 26752 2372
rect 27344 2363 27396 2372
rect 27344 2329 27353 2363
rect 27353 2329 27387 2363
rect 27387 2329 27396 2363
rect 27344 2320 27396 2329
rect 12808 2252 12860 2304
rect 13544 2252 13596 2304
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 15016 2252 15068 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 19340 2252 19392 2304
rect 19432 2252 19484 2304
rect 25780 2252 25832 2304
rect 27160 2252 27212 2304
rect 30012 2320 30064 2372
rect 31392 2320 31444 2372
rect 28724 2252 28776 2304
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 34244 2388 34296 2440
rect 34612 2388 34664 2440
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 37832 2388 37884 2440
rect 35716 2320 35768 2372
rect 36728 2252 36780 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 7564 2048 7616 2100
rect 31116 2048 31168 2100
rect 2872 1980 2924 2032
rect 12348 1980 12400 2032
rect 13544 1980 13596 2032
rect 3976 1912 4028 1964
rect 14188 1912 14240 1964
rect 22100 1912 22152 1964
rect 28724 1912 28776 1964
rect 12532 1844 12584 1896
rect 23020 1844 23072 1896
rect 12440 1776 12492 1828
rect 13912 1776 13964 1828
rect 16856 1776 16908 1828
rect 26608 1844 26660 1896
rect 34520 1844 34572 1896
rect 23940 1776 23992 1828
rect 24400 1776 24452 1828
rect 16120 1708 16172 1760
rect 36176 1708 36228 1760
rect 19340 1640 19392 1692
rect 26424 1640 26476 1692
rect 27252 1640 27304 1692
rect 29092 1640 29144 1692
rect 30012 1640 30064 1692
rect 28448 1572 28500 1624
<< metal2 >>
rect 110 39200 166 40000
rect 386 39200 442 40000
rect 754 39200 810 40000
rect 1122 39200 1178 40000
rect 1490 39200 1546 40000
rect 1858 39200 1914 40000
rect 2134 39200 2190 40000
rect 2502 39200 2558 40000
rect 2870 39200 2926 40000
rect 3238 39200 3294 40000
rect 3606 39200 3662 40000
rect 3882 39200 3938 40000
rect 4250 39200 4306 40000
rect 4618 39200 4674 40000
rect 4986 39200 5042 40000
rect 5354 39200 5410 40000
rect 5722 39200 5778 40000
rect 5998 39200 6054 40000
rect 6366 39200 6422 40000
rect 6734 39200 6790 40000
rect 7102 39200 7158 40000
rect 7470 39200 7526 40000
rect 7746 39200 7802 40000
rect 8114 39200 8170 40000
rect 8482 39200 8538 40000
rect 8850 39200 8906 40000
rect 9218 39200 9274 40000
rect 9586 39200 9642 40000
rect 9862 39200 9918 40000
rect 10230 39200 10286 40000
rect 10598 39200 10654 40000
rect 10966 39200 11022 40000
rect 11334 39200 11390 40000
rect 11610 39200 11666 40000
rect 11978 39200 12034 40000
rect 12346 39200 12402 40000
rect 12714 39200 12770 40000
rect 13082 39200 13138 40000
rect 13450 39200 13506 40000
rect 13726 39200 13782 40000
rect 14094 39200 14150 40000
rect 14462 39200 14518 40000
rect 14830 39200 14886 40000
rect 15198 39200 15254 40000
rect 15474 39200 15530 40000
rect 15842 39200 15898 40000
rect 16210 39200 16266 40000
rect 16578 39200 16634 40000
rect 16946 39200 17002 40000
rect 17222 39200 17278 40000
rect 17590 39200 17646 40000
rect 17958 39200 18014 40000
rect 18326 39200 18382 40000
rect 18694 39200 18750 40000
rect 19062 39200 19118 40000
rect 19338 39200 19394 40000
rect 19706 39200 19762 40000
rect 19812 39222 20024 39250
rect 124 36854 152 39200
rect 112 36848 164 36854
rect 112 36790 164 36796
rect 400 36378 428 39200
rect 388 36372 440 36378
rect 388 36314 440 36320
rect 768 35834 796 39200
rect 1136 37262 1164 39200
rect 1124 37256 1176 37262
rect 1124 37198 1176 37204
rect 1504 36582 1532 39200
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1584 36848 1636 36854
rect 1584 36790 1636 36796
rect 1492 36576 1544 36582
rect 1492 36518 1544 36524
rect 756 35828 808 35834
rect 756 35770 808 35776
rect 1596 35290 1624 36790
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1584 35284 1636 35290
rect 1584 35226 1636 35232
rect 1688 35222 1716 36110
rect 1780 35290 1808 37198
rect 1872 36378 1900 39200
rect 2148 37262 2176 39200
rect 2136 37256 2188 37262
rect 2136 37198 2188 37204
rect 1952 37120 2004 37126
rect 1952 37062 2004 37068
rect 1860 36372 1912 36378
rect 1860 36314 1912 36320
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 1676 35216 1728 35222
rect 1676 35158 1728 35164
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 30025 1624 30194
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1596 29850 1624 29951
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1964 8401 1992 37062
rect 2516 36922 2544 39200
rect 2596 37256 2648 37262
rect 2596 37198 2648 37204
rect 2504 36916 2556 36922
rect 2504 36858 2556 36864
rect 2044 36644 2096 36650
rect 2044 36586 2096 36592
rect 2056 11354 2084 36586
rect 2608 34746 2636 37198
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2792 36786 2820 37062
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2884 36378 2912 39200
rect 3252 37262 3280 39200
rect 3516 37324 3568 37330
rect 3516 37266 3568 37272
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 3240 36780 3292 36786
rect 3240 36722 3292 36728
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 3056 36168 3108 36174
rect 3056 36110 3108 36116
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 3068 34678 3096 36110
rect 3148 36100 3200 36106
rect 3148 36042 3200 36048
rect 3160 35834 3188 36042
rect 3148 35828 3200 35834
rect 3148 35770 3200 35776
rect 3148 35692 3200 35698
rect 3148 35634 3200 35640
rect 3056 34672 3108 34678
rect 3056 34614 3108 34620
rect 2872 34536 2924 34542
rect 2872 34478 2924 34484
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2792 18426 2820 21490
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2056 11150 2084 11290
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1950 8392 2006 8401
rect 1950 8327 2006 8336
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 296 4072 348 4078
rect 296 4014 348 4020
rect 112 2848 164 2854
rect 112 2790 164 2796
rect 124 800 152 2790
rect 308 800 336 4014
rect 584 800 612 4082
rect 848 3596 900 3602
rect 848 3538 900 3544
rect 860 800 888 3538
rect 1412 3058 1440 5510
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1124 3052 1176 3058
rect 1124 2994 1176 3000
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1136 800 1164 2994
rect 1400 2848 1452 2854
rect 1504 2836 1532 4966
rect 1596 4622 1624 6054
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 4078 1624 4558
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1688 3534 1716 5510
rect 1780 4622 1808 5578
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1452 2808 1532 2836
rect 1400 2790 1452 2796
rect 1412 2514 1440 2790
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1412 800 1440 2314
rect 1688 800 1716 3470
rect 1780 2378 1808 4558
rect 1964 4146 1992 4966
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2424 4010 2452 11698
rect 2884 10266 2912 34478
rect 3068 11830 3096 34614
rect 3160 26234 3188 35634
rect 3252 34542 3280 36722
rect 3240 34536 3292 34542
rect 3240 34478 3292 34484
rect 3160 26206 3280 26234
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3160 17882 3188 18226
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3252 10810 3280 26206
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2792 8634 2820 9930
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2976 8566 3004 8774
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 3068 8362 3096 8842
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 4622 2544 6054
rect 2792 5642 2820 6190
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 1964 800 1992 3606
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 2516 800 2544 4558
rect 2608 2446 2636 4966
rect 2792 3942 2820 5578
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2884 4146 2912 4694
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 2990 2820 3878
rect 2976 3602 3004 4966
rect 3068 4078 3096 8298
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3194 3004 3334
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 3068 2514 3096 4014
rect 3160 3670 3188 5510
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 2596 2440 2648 2446
rect 2872 2440 2924 2446
rect 2596 2382 2648 2388
rect 2792 2388 2872 2394
rect 3252 2394 3280 4082
rect 3344 3194 3372 11698
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10033 3464 10950
rect 3422 10024 3478 10033
rect 3422 9959 3478 9968
rect 3528 9178 3556 37266
rect 3620 36922 3648 39200
rect 3608 36916 3660 36922
rect 3608 36858 3660 36864
rect 3896 36378 3924 39200
rect 4264 37754 4292 39200
rect 4080 37726 4292 37754
rect 4080 37346 4108 37726
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4080 37318 4200 37346
rect 4068 37256 4120 37262
rect 4068 37198 4120 37204
rect 3884 36372 3936 36378
rect 3884 36314 3936 36320
rect 4080 35834 4108 37198
rect 4172 37194 4200 37318
rect 4160 37188 4212 37194
rect 4160 37130 4212 37136
rect 4632 36922 4660 39200
rect 4896 37460 4948 37466
rect 4896 37402 4948 37408
rect 4620 36916 4672 36922
rect 4620 36858 4672 36864
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4632 35894 4660 36722
rect 4632 35866 4752 35894
rect 4068 35828 4120 35834
rect 4068 35770 4120 35776
rect 3700 35692 3752 35698
rect 3700 35634 3752 35640
rect 3712 35494 3740 35634
rect 3700 35488 3752 35494
rect 3700 35430 3752 35436
rect 3608 30660 3660 30666
rect 3608 30602 3660 30608
rect 3620 30326 3648 30602
rect 3608 30320 3660 30326
rect 3608 30262 3660 30268
rect 3712 10606 3740 35430
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4724 34950 4752 35866
rect 3884 34944 3936 34950
rect 3884 34886 3936 34892
rect 4712 34944 4764 34950
rect 4712 34886 4764 34892
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3804 25906 3832 26182
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 13938 3832 15302
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3896 9450 3924 34886
rect 4160 34536 4212 34542
rect 4080 34484 4160 34490
rect 4080 34478 4212 34484
rect 4080 34462 4200 34478
rect 4080 30734 4108 34462
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 4080 30190 4108 30534
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 4264 26234 4292 26318
rect 4172 26206 4292 26234
rect 4172 26042 4200 26206
rect 4160 26036 4212 26042
rect 4160 25978 4212 25984
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4632 20534 4660 21626
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4632 19854 4660 20470
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3988 17678 4016 18022
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3988 15502 4016 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4632 15706 4660 17478
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 3976 15496 4028 15502
rect 4160 15496 4212 15502
rect 3976 15438 4028 15444
rect 4080 15444 4160 15450
rect 4080 15438 4212 15444
rect 4080 15422 4200 15438
rect 4080 15026 4108 15422
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14074 4108 14962
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4724 12434 4752 34886
rect 4908 33454 4936 37402
rect 5000 36922 5028 39200
rect 5080 37324 5132 37330
rect 5080 37266 5132 37272
rect 4988 36916 5040 36922
rect 4988 36858 5040 36864
rect 4988 36168 5040 36174
rect 4988 36110 5040 36116
rect 5000 34932 5028 36110
rect 5092 35894 5120 37266
rect 5264 37188 5316 37194
rect 5264 37130 5316 37136
rect 5092 35866 5212 35894
rect 5080 34944 5132 34950
rect 5000 34904 5080 34932
rect 5080 34886 5132 34892
rect 4896 33448 4948 33454
rect 4896 33390 4948 33396
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 4816 30734 4844 33254
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4816 30394 4844 30670
rect 4896 30592 4948 30598
rect 4896 30534 4948 30540
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4908 30258 4936 30534
rect 4896 30252 4948 30258
rect 4896 30194 4948 30200
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4816 27606 4844 29990
rect 4804 27600 4856 27606
rect 4804 27542 4856 27548
rect 4816 27470 4844 27542
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 4908 27402 4936 29990
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 4908 26382 4936 27338
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4816 18222 4844 19858
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4816 17746 4844 18158
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4816 16794 4844 17682
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4908 16182 4936 17478
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4632 12406 4752 12434
rect 4632 12374 4660 12406
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 4632 8634 4660 9590
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3436 7750 3464 8434
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 2792 2382 2924 2388
rect 2792 2366 2912 2382
rect 3068 2366 3280 2394
rect 2792 800 2820 2366
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 2038 2912 2246
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 3068 800 3096 2366
rect 3344 800 3372 2994
rect 3436 2417 3464 7686
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4724 5914 4752 12106
rect 5092 11830 5120 34886
rect 5184 33538 5212 35866
rect 5276 35834 5304 37130
rect 5368 36938 5396 39200
rect 5736 37346 5764 39200
rect 5736 37318 5856 37346
rect 5724 37256 5776 37262
rect 5724 37198 5776 37204
rect 5368 36910 5672 36938
rect 5644 36786 5672 36910
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 5540 36780 5592 36786
rect 5540 36722 5592 36728
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 5368 36378 5396 36722
rect 5356 36372 5408 36378
rect 5356 36314 5408 36320
rect 5264 35828 5316 35834
rect 5264 35770 5316 35776
rect 5552 34950 5580 36722
rect 5736 35494 5764 37198
rect 5828 36922 5856 37318
rect 5816 36916 5868 36922
rect 5816 36858 5868 36864
rect 6012 36378 6040 39200
rect 6380 37262 6408 39200
rect 6368 37256 6420 37262
rect 6368 37198 6420 37204
rect 6184 36780 6236 36786
rect 6184 36722 6236 36728
rect 6000 36372 6052 36378
rect 6000 36314 6052 36320
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5540 34944 5592 34950
rect 5540 34886 5592 34892
rect 5264 34604 5316 34610
rect 5264 34546 5316 34552
rect 5276 33658 5304 34546
rect 5264 33652 5316 33658
rect 5264 33594 5316 33600
rect 5184 33510 5304 33538
rect 5172 33448 5224 33454
rect 5172 33390 5224 33396
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4710 5672 4766 5681
rect 4710 5607 4712 5616
rect 4764 5607 4766 5616
rect 4712 5578 4764 5584
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3422 2408 3478 2417
rect 3422 2343 3478 2352
rect 3620 800 3648 3946
rect 3712 3058 3740 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3884 4480 3936 4486
rect 3882 4448 3884 4457
rect 4160 4480 4212 4486
rect 3936 4448 3938 4457
rect 4160 4422 4212 4428
rect 3882 4383 3938 4392
rect 3896 4282 3924 4383
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 4172 4026 4200 4422
rect 4080 3998 4200 4026
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3896 800 3924 2926
rect 4080 2446 4108 3998
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4158 3360 4214 3369
rect 4158 3295 4214 3304
rect 4172 3126 4200 3295
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4448 2922 4476 3470
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4540 3194 4568 3402
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 2514 4660 4966
rect 4724 3058 4752 5034
rect 4816 4146 4844 6054
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3346 4936 4082
rect 5000 3738 5028 10610
rect 5184 6458 5212 33390
rect 5276 9178 5304 33510
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5368 26450 5396 27270
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5552 10742 5580 34886
rect 5632 30320 5684 30326
rect 5632 30262 5684 30268
rect 5644 27538 5672 30262
rect 5632 27532 5684 27538
rect 5632 27474 5684 27480
rect 5644 26586 5672 27474
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5644 21010 5672 26522
rect 5736 22094 5764 35430
rect 6196 35290 6224 36722
rect 6380 36582 6408 37198
rect 6748 36666 6776 39200
rect 7116 37210 7144 39200
rect 7484 37262 7512 39200
rect 7656 37392 7708 37398
rect 7656 37334 7708 37340
rect 7472 37256 7524 37262
rect 7116 37182 7236 37210
rect 7472 37198 7524 37204
rect 7104 36780 7156 36786
rect 7104 36722 7156 36728
rect 6748 36650 6960 36666
rect 6644 36644 6696 36650
rect 6748 36644 6972 36650
rect 6748 36638 6920 36644
rect 6644 36586 6696 36592
rect 6920 36586 6972 36592
rect 6368 36576 6420 36582
rect 6368 36518 6420 36524
rect 6460 36100 6512 36106
rect 6460 36042 6512 36048
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 5816 34400 5868 34406
rect 5816 34342 5868 34348
rect 5828 33454 5856 34342
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 6368 33448 6420 33454
rect 6368 33390 6420 33396
rect 6380 30326 6408 33390
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 6184 30116 6236 30122
rect 6184 30058 6236 30064
rect 6196 28762 6224 30058
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6196 28558 6224 28698
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 5736 22066 5856 22094
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5828 9178 5856 22066
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6380 21146 6408 21898
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8498 5396 8842
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5920 8634 5948 8774
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5092 4214 5120 5510
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4816 3318 4936 3346
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3988 1970 4016 2246
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 4172 800 4200 2314
rect 4448 800 4476 2450
rect 4724 800 4752 2858
rect 4816 2378 4844 3318
rect 4894 3224 4950 3233
rect 4894 3159 4950 3168
rect 4908 3126 4936 3159
rect 5092 3126 5120 3878
rect 5184 3602 5212 4762
rect 5276 4622 5304 6598
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 5000 800 5028 2382
rect 5276 800 5304 4558
rect 5368 3942 5396 8434
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 4146 5488 6054
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 4214 5672 5510
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5460 2922 5488 4082
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3602 5580 3878
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5552 2961 5580 3130
rect 5538 2952 5594 2961
rect 5448 2916 5500 2922
rect 5644 2922 5672 3946
rect 5828 3058 5856 4966
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 3777 6132 4422
rect 6090 3768 6146 3777
rect 6196 3738 6224 9930
rect 6472 8566 6500 36042
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21350 6592 21830
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6564 20602 6592 20946
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6656 7274 6684 36586
rect 6736 36576 6788 36582
rect 6736 36518 6788 36524
rect 6748 35290 6776 36518
rect 7012 36168 7064 36174
rect 7012 36110 7064 36116
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 7024 34932 7052 36110
rect 7116 35834 7144 36722
rect 7208 36378 7236 37182
rect 7484 36854 7512 37198
rect 7472 36848 7524 36854
rect 7472 36790 7524 36796
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7470 36272 7526 36281
rect 7470 36207 7526 36216
rect 7484 36174 7512 36207
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7104 35828 7156 35834
rect 7104 35770 7156 35776
rect 7484 35290 7512 36110
rect 7668 35894 7696 37334
rect 7760 36922 7788 39200
rect 7840 37120 7892 37126
rect 7840 37062 7892 37068
rect 7748 36916 7800 36922
rect 7748 36858 7800 36864
rect 7668 35866 7788 35894
rect 7472 35284 7524 35290
rect 7472 35226 7524 35232
rect 7104 34944 7156 34950
rect 7024 34904 7104 34932
rect 7104 34886 7156 34892
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6840 32570 6868 33458
rect 6828 32564 6880 32570
rect 6828 32506 6880 32512
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6932 28762 6960 30534
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6748 25158 6776 28494
rect 6932 27606 6960 28698
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20058 6776 20878
rect 6932 20398 6960 22034
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6932 19990 6960 20334
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 7024 19854 7052 20538
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 7024 16794 7052 17002
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16114 6868 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6840 14482 6868 16050
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6932 14006 6960 15302
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6932 12850 6960 13942
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7116 10198 7144 34886
rect 7656 33312 7708 33318
rect 7656 33254 7708 33260
rect 7668 32434 7696 33254
rect 7656 32428 7708 32434
rect 7656 32370 7708 32376
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 7484 30598 7512 32166
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7668 30326 7696 32370
rect 7656 30320 7708 30326
rect 7656 30262 7708 30268
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19854 7420 20334
rect 7484 19990 7512 20402
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7392 17882 7420 19790
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17678 7420 17818
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17202 7420 17614
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7576 17134 7604 19722
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 15026 7236 16458
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7300 14414 7328 16934
rect 7576 15162 7604 17070
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 12850 7236 14214
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7760 12306 7788 35866
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7852 11830 7880 37062
rect 7932 36780 7984 36786
rect 7932 36722 7984 36728
rect 7944 36378 7972 36722
rect 7932 36372 7984 36378
rect 8128 36360 8156 39200
rect 8496 37262 8524 39200
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8864 36922 8892 39200
rect 9232 37618 9260 39200
rect 9232 37590 9352 37618
rect 8852 36916 8904 36922
rect 8852 36858 8904 36864
rect 8576 36780 8628 36786
rect 8576 36722 8628 36728
rect 8300 36372 8352 36378
rect 8128 36332 8300 36360
rect 7932 36314 7984 36320
rect 8300 36314 8352 36320
rect 8024 36168 8076 36174
rect 8024 36110 8076 36116
rect 8036 35494 8064 36110
rect 8588 35834 8616 36722
rect 9232 36174 9260 36205
rect 9220 36168 9272 36174
rect 9218 36136 9220 36145
rect 9272 36136 9274 36145
rect 9218 36071 9274 36080
rect 8576 35828 8628 35834
rect 8576 35770 8628 35776
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 8116 35556 8168 35562
rect 8116 35498 8168 35504
rect 8024 35488 8076 35494
rect 8024 35430 8076 35436
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7944 24954 7972 25162
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 8036 24274 8064 35430
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 8128 7478 8156 35498
rect 8864 34950 8892 35634
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 8208 30592 8260 30598
rect 8208 30534 8260 30540
rect 8220 29850 8248 30534
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8404 26042 8432 29106
rect 8392 26036 8444 26042
rect 8392 25978 8444 25984
rect 8404 25770 8432 25978
rect 8392 25764 8444 25770
rect 8392 25706 8444 25712
rect 8404 25294 8432 25706
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8864 24342 8892 34886
rect 9232 34746 9260 36071
rect 9324 35834 9352 37590
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 9416 36718 9444 37198
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9312 35828 9364 35834
rect 9312 35770 9364 35776
rect 9600 35290 9628 39200
rect 9680 37664 9732 37670
rect 9680 37606 9732 37612
rect 9692 37466 9720 37606
rect 9680 37460 9732 37466
rect 9680 37402 9732 37408
rect 9772 36780 9824 36786
rect 9772 36722 9824 36728
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 9220 34740 9272 34746
rect 9220 34682 9272 34688
rect 9496 34672 9548 34678
rect 9496 34614 9548 34620
rect 9508 33998 9536 34614
rect 9784 34542 9812 36722
rect 9876 36378 9904 39200
rect 10140 37256 10192 37262
rect 10140 37198 10192 37204
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 10152 35290 10180 37198
rect 10244 36378 10272 39200
rect 10612 37262 10640 39200
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 10232 36372 10284 36378
rect 10232 36314 10284 36320
rect 10232 36168 10284 36174
rect 10232 36110 10284 36116
rect 10244 35290 10272 36110
rect 10140 35284 10192 35290
rect 10140 35226 10192 35232
rect 10232 35284 10284 35290
rect 10232 35226 10284 35232
rect 10612 35170 10640 37062
rect 10980 36922 11008 39200
rect 10968 36916 11020 36922
rect 10968 36858 11020 36864
rect 10692 36780 10744 36786
rect 10692 36722 10744 36728
rect 10704 35834 10732 36722
rect 11348 36378 11376 39200
rect 11624 37194 11652 39200
rect 11612 37188 11664 37194
rect 11612 37130 11664 37136
rect 11992 36922 12020 39200
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 12072 37120 12124 37126
rect 12072 37062 12124 37068
rect 11980 36916 12032 36922
rect 11980 36858 12032 36864
rect 11336 36372 11388 36378
rect 11336 36314 11388 36320
rect 11704 36168 11756 36174
rect 11704 36110 11756 36116
rect 11716 35834 11744 36110
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11060 35692 11112 35698
rect 11060 35634 11112 35640
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 10612 35142 10732 35170
rect 10600 35080 10652 35086
rect 10600 35022 10652 35028
rect 10612 34542 10640 35022
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 10600 34536 10652 34542
rect 10600 34478 10652 34484
rect 9496 33992 9548 33998
rect 9496 33934 9548 33940
rect 9508 29782 9536 33934
rect 9496 29776 9548 29782
rect 9496 29718 9548 29724
rect 9508 29306 9536 29718
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9692 24886 9720 25094
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8220 17678 8248 19926
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8220 16454 8248 17614
rect 8496 17338 8524 17614
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14414 8340 14894
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8312 12986 8340 14350
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 9784 12714 9812 34478
rect 10140 33924 10192 33930
rect 10140 33866 10192 33872
rect 10152 33658 10180 33866
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10152 24682 10180 29514
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10060 19718 10088 19994
rect 10152 19854 10180 24618
rect 10612 23798 10640 34478
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10244 20466 10272 20946
rect 10428 20806 10456 21286
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10428 20058 10456 20742
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 15366 10088 19654
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10704 13326 10732 35142
rect 11072 34950 11100 35634
rect 11244 35624 11296 35630
rect 11244 35566 11296 35572
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 10784 33856 10836 33862
rect 10784 33798 10836 33804
rect 10796 33658 10824 33798
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10796 33522 10824 33594
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10968 30320 11020 30326
rect 10968 30262 11020 30268
rect 10980 29646 11008 30262
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 10980 24818 11008 25162
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10980 24206 11008 24754
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 11072 22094 11100 34886
rect 11256 34542 11284 35566
rect 11716 34950 11744 35634
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11244 34536 11296 34542
rect 11244 34478 11296 34484
rect 11256 26234 11284 34478
rect 11520 30320 11572 30326
rect 11440 30268 11520 30274
rect 11440 30262 11572 30268
rect 11440 30246 11560 30262
rect 11440 30190 11468 30246
rect 11428 30184 11480 30190
rect 11348 30132 11428 30138
rect 11348 30126 11480 30132
rect 11348 30110 11468 30126
rect 11348 29578 11376 30110
rect 11440 30061 11468 30110
rect 11612 30116 11664 30122
rect 11612 30058 11664 30064
rect 11520 29776 11572 29782
rect 11520 29718 11572 29724
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 11348 29034 11376 29514
rect 11532 29170 11560 29718
rect 11624 29170 11652 30058
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11612 29164 11664 29170
rect 11612 29106 11664 29112
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 11716 26234 11744 34886
rect 11796 33652 11848 33658
rect 11796 33594 11848 33600
rect 11808 30410 11836 33594
rect 11808 30394 11928 30410
rect 11808 30388 11940 30394
rect 11808 30382 11888 30388
rect 11808 30054 11836 30382
rect 11888 30330 11940 30336
rect 11796 30048 11848 30054
rect 11796 29990 11848 29996
rect 11808 29646 11836 29990
rect 11796 29640 11848 29646
rect 11796 29582 11848 29588
rect 11256 26206 11468 26234
rect 11072 22066 11192 22094
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20602 11100 20810
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11164 13394 11192 22066
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 11440 12238 11468 26206
rect 11624 26206 11744 26234
rect 12084 26234 12112 37062
rect 12176 35290 12204 37198
rect 12254 36408 12310 36417
rect 12254 36343 12310 36352
rect 12360 36360 12388 39200
rect 12728 36854 12756 39200
rect 13096 36922 13124 39200
rect 13084 36916 13136 36922
rect 13084 36858 13136 36864
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 12440 36372 12492 36378
rect 12268 36106 12296 36343
rect 12360 36332 12440 36360
rect 12440 36314 12492 36320
rect 12256 36100 12308 36106
rect 12256 36042 12308 36048
rect 12164 35284 12216 35290
rect 12164 35226 12216 35232
rect 12268 34746 12296 36042
rect 12624 35692 12676 35698
rect 12624 35634 12676 35640
rect 12636 35494 12664 35634
rect 12624 35488 12676 35494
rect 12624 35430 12676 35436
rect 12256 34740 12308 34746
rect 12256 34682 12308 34688
rect 12084 26206 12204 26234
rect 11520 25424 11572 25430
rect 11520 25366 11572 25372
rect 11532 24954 11560 25366
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 11532 24818 11560 24890
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9600 9110 9628 9454
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6656 6866 6684 7210
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 4146 6408 5510
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6090 3703 6146 3712
rect 6184 3732 6236 3738
rect 6104 3466 6132 3703
rect 6184 3674 6236 3680
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5538 2887 5594 2896
rect 5632 2916 5684 2922
rect 5448 2858 5500 2864
rect 5632 2858 5684 2864
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 800 5580 2790
rect 5828 800 5856 2994
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6104 800 6132 2314
rect 6380 800 6408 4082
rect 6472 2446 6500 4966
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 3058 6592 4422
rect 6656 3942 6684 5646
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6748 3602 6776 7278
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 6932 4622 6960 5510
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6840 1714 6868 3402
rect 6656 1686 6868 1714
rect 6656 800 6684 1686
rect 6932 800 6960 4558
rect 7208 4214 7236 4966
rect 7760 4554 7788 4966
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7208 800 7236 4150
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7576 3738 7604 4014
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 800 7512 3470
rect 7656 3392 7708 3398
rect 7576 3340 7656 3346
rect 7576 3334 7708 3340
rect 7576 3318 7696 3334
rect 7576 2854 7604 3318
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7576 2106 7604 2790
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7760 800 7788 4490
rect 7944 4010 7972 4558
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 8036 3058 8064 5510
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4214 8156 4422
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8036 800 8064 2994
rect 8128 2446 8156 3878
rect 8220 3534 8248 4966
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 3754 8340 4626
rect 8496 4282 8524 4694
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8588 4078 8616 4966
rect 9048 4554 9076 8842
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8496 3913 8524 4014
rect 8482 3904 8538 3913
rect 8482 3839 8538 3848
rect 8312 3726 8432 3754
rect 8300 3664 8352 3670
rect 8298 3632 8300 3641
rect 8352 3632 8354 3641
rect 8404 3602 8432 3726
rect 8298 3567 8354 3576
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8392 3392 8444 3398
rect 8206 3360 8262 3369
rect 8392 3334 8444 3340
rect 8206 3295 8262 3304
rect 8220 3194 8248 3295
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8312 800 8340 2314
rect 8404 1601 8432 3334
rect 8390 1592 8446 1601
rect 8390 1527 8446 1536
rect 8588 800 8616 4014
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8864 800 8892 2790
rect 9048 2514 9076 4490
rect 9218 4176 9274 4185
rect 9218 4111 9274 4120
rect 9232 2990 9260 4111
rect 9416 3534 9444 5510
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9140 800 9168 2450
rect 9416 800 9444 3470
rect 9508 3194 9536 8842
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8498 9812 8774
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9600 2514 9628 4966
rect 9692 4078 9720 7822
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9876 3602 9904 11562
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9968 7857 9996 8502
rect 9954 7848 10010 7857
rect 9954 7783 10010 7792
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 2990 9904 3402
rect 9968 2990 9996 4422
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9692 800 9720 2586
rect 9968 800 9996 2926
rect 10060 2582 10088 4014
rect 10152 3058 10180 4966
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10336 2514 10364 11494
rect 10888 11150 10916 11630
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10598 4040 10654 4049
rect 10598 3975 10600 3984
rect 10652 3975 10654 3984
rect 10600 3946 10652 3952
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10506 2816 10562 2825
rect 10506 2751 10562 2760
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10244 800 10272 2382
rect 10520 800 10548 2751
rect 10612 2292 10640 2994
rect 10704 2446 10732 4966
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 2922 10824 3538
rect 10888 3466 10916 11086
rect 11624 9110 11652 26206
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 15434 12112 16390
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11428 7812 11480 7818
rect 11428 7754 11480 7760
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 4622 11192 5510
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3505 11008 3878
rect 10966 3496 11022 3505
rect 10876 3460 10928 3466
rect 10966 3431 11022 3440
rect 10876 3402 10928 3408
rect 11060 3392 11112 3398
rect 11058 3360 11060 3369
rect 11112 3360 11114 3369
rect 11058 3295 11114 3304
rect 11164 3210 11192 4558
rect 11072 3182 11192 3210
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10782 2680 10838 2689
rect 10782 2615 10838 2624
rect 10796 2446 10824 2615
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10612 2264 10824 2292
rect 10796 800 10824 2264
rect 11072 800 11100 3182
rect 11256 2378 11284 4966
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11348 3505 11376 4082
rect 11440 4010 11468 7754
rect 11532 7410 11560 8230
rect 11624 7886 11652 8366
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11716 6914 11744 12310
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11624 6886 11744 6914
rect 11518 4040 11574 4049
rect 11428 4004 11480 4010
rect 11518 3975 11574 3984
rect 11428 3946 11480 3952
rect 11532 3738 11560 3975
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11334 3496 11390 3505
rect 11334 3431 11390 3440
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11440 3126 11468 3402
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11624 3058 11652 6886
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11716 4146 11744 5102
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11716 2938 11744 4082
rect 11808 3058 11836 8298
rect 12176 6914 12204 26206
rect 12348 24880 12400 24886
rect 12348 24822 12400 24828
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12268 19514 12296 20334
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12360 17134 12388 24822
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12452 24410 12480 24686
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12544 24070 12572 24754
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12544 19854 12572 24006
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19446 12572 19790
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 17202 12480 17478
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12544 17066 12572 19110
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16590 12296 16934
rect 12544 16590 12572 17002
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12544 15706 12572 16526
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 10674 12572 11494
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12636 9042 12664 35430
rect 12728 35290 12756 36790
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 12900 36100 12952 36106
rect 12900 36042 12952 36048
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 12912 34746 12940 36042
rect 13372 35018 13400 36722
rect 13464 36378 13492 39200
rect 13740 37346 13768 39200
rect 13740 37318 13860 37346
rect 13832 37262 13860 37318
rect 13820 37256 13872 37262
rect 13820 37198 13872 37204
rect 13728 37188 13780 37194
rect 13728 37130 13780 37136
rect 13740 36854 13768 37130
rect 14108 36922 14136 39200
rect 14096 36916 14148 36922
rect 14096 36858 14148 36864
rect 13728 36848 13780 36854
rect 13728 36790 13780 36796
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 13636 36644 13688 36650
rect 13636 36586 13688 36592
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13452 36168 13504 36174
rect 13452 36110 13504 36116
rect 13464 35494 13492 36110
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13360 35012 13412 35018
rect 13360 34954 13412 34960
rect 12900 34740 12952 34746
rect 12900 34682 12952 34688
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 13096 26790 13124 29038
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13096 25498 13124 26726
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 13004 24954 13032 25162
rect 12992 24948 13044 24954
rect 12992 24890 13044 24896
rect 13096 24818 13124 25434
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13096 19990 13124 20742
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12820 19446 12848 19654
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12820 17202 12848 19382
rect 12912 19310 12940 19654
rect 13096 19378 13124 19926
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12084 6886 12204 6914
rect 12084 6225 12112 6886
rect 12070 6216 12126 6225
rect 12070 6151 12126 6160
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12268 4758 12296 5238
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12256 4752 12308 4758
rect 12308 4712 12480 4740
rect 12256 4694 12308 4700
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11992 4026 12020 4082
rect 12268 4078 12296 4218
rect 12256 4072 12308 4078
rect 11900 3998 12020 4026
rect 12070 4040 12126 4049
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11624 2910 11744 2938
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11348 800 11376 2858
rect 11624 800 11652 2910
rect 11900 800 11928 3998
rect 12256 4014 12308 4020
rect 12070 3975 12126 3984
rect 12084 3641 12112 3975
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12070 3632 12126 3641
rect 12070 3567 12126 3576
rect 12176 800 12204 3878
rect 12360 3534 12388 4422
rect 12452 3584 12480 4712
rect 12544 4146 12572 4966
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12532 3596 12584 3602
rect 12452 3556 12532 3584
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12452 2938 12480 3556
rect 12532 3538 12584 3544
rect 12636 3058 12664 7142
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 4826 12756 5510
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12360 2910 12480 2938
rect 12360 2038 12388 2910
rect 12440 2848 12492 2854
rect 12438 2816 12440 2825
rect 12492 2816 12494 2825
rect 12438 2751 12494 2760
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12348 2032 12400 2038
rect 12348 1974 12400 1980
rect 12544 1902 12572 2314
rect 12532 1896 12584 1902
rect 12532 1838 12584 1844
rect 12440 1828 12492 1834
rect 12440 1770 12492 1776
rect 12452 800 12480 1770
rect 12728 800 12756 4558
rect 13004 4146 13032 10406
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 2310 12848 3334
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 13004 800 13032 3946
rect 13188 3738 13216 12786
rect 13280 5302 13308 13126
rect 13464 12434 13492 35430
rect 13648 31754 13676 36586
rect 13912 36168 13964 36174
rect 13912 36110 13964 36116
rect 13924 34610 13952 36110
rect 14292 35834 14320 36722
rect 14476 36378 14504 39200
rect 14556 37460 14608 37466
rect 14556 37402 14608 37408
rect 14568 37262 14596 37402
rect 14844 37262 14872 39200
rect 14924 37324 14976 37330
rect 14924 37266 14976 37272
rect 14556 37256 14608 37262
rect 14556 37198 14608 37204
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 14832 36712 14884 36718
rect 14832 36654 14884 36660
rect 14464 36372 14516 36378
rect 14464 36314 14516 36320
rect 14556 36168 14608 36174
rect 14556 36110 14608 36116
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14200 34950 14228 35634
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 13728 34536 13780 34542
rect 13728 34478 13780 34484
rect 13740 33862 13768 34478
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13740 32434 13768 33798
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13648 31726 13768 31754
rect 13740 14618 13768 31726
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13740 13802 13768 14554
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13924 12918 13952 34546
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24818 14136 25094
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14108 24206 14136 24754
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13372 12406 13492 12434
rect 13372 8022 13400 12406
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13464 9586 13492 9862
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4622 13400 4966
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13280 800 13308 3062
rect 13464 800 13492 4558
rect 13648 3194 13676 11018
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 4146 13768 9318
rect 13832 5778 13860 9522
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 2038 13584 2246
rect 13544 2032 13596 2038
rect 13544 1974 13596 1980
rect 13740 800 13768 3878
rect 13832 2378 13860 5714
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 3058 13952 4422
rect 14016 3738 14044 13874
rect 14200 7478 14228 34886
rect 14568 34610 14596 36110
rect 14844 35834 14872 36654
rect 14832 35828 14884 35834
rect 14832 35770 14884 35776
rect 14740 35692 14792 35698
rect 14740 35634 14792 35640
rect 14752 34610 14780 35634
rect 14280 34604 14332 34610
rect 14280 34546 14332 34552
rect 14556 34604 14608 34610
rect 14556 34546 14608 34552
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14292 14006 14320 34546
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14384 30326 14412 32370
rect 14372 30320 14424 30326
rect 14372 30262 14424 30268
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 25430 14504 25638
rect 14464 25424 14516 25430
rect 14464 25366 14516 25372
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14660 14346 14688 14758
rect 14752 14618 14780 34546
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14660 13870 14688 14282
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14660 13190 14688 13806
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11150 14596 12038
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9586 14320 9930
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13924 1834 13952 2994
rect 14108 2446 14136 4966
rect 14200 4622 14228 5510
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14188 3596 14240 3602
rect 14292 3584 14320 7278
rect 14936 7274 14964 37266
rect 15212 36922 15240 39200
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15304 36242 15332 37198
rect 15384 36712 15436 36718
rect 15384 36654 15436 36660
rect 15292 36236 15344 36242
rect 15292 36178 15344 36184
rect 15396 35290 15424 36654
rect 15488 35834 15516 39200
rect 15856 37194 15884 39200
rect 16028 37664 16080 37670
rect 16028 37606 16080 37612
rect 16040 37466 16068 37606
rect 16028 37460 16080 37466
rect 16028 37402 16080 37408
rect 16028 37324 16080 37330
rect 16028 37266 16080 37272
rect 15844 37188 15896 37194
rect 15844 37130 15896 37136
rect 15476 35828 15528 35834
rect 15476 35770 15528 35776
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15384 35284 15436 35290
rect 15384 35226 15436 35232
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 15752 35080 15804 35086
rect 15752 35022 15804 35028
rect 15120 34746 15148 35022
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14936 7002 14964 7210
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14240 3556 14320 3584
rect 14188 3538 14240 3544
rect 14096 2440 14148 2446
rect 14016 2400 14096 2428
rect 13912 1828 13964 1834
rect 13912 1770 13964 1776
rect 14016 800 14044 2400
rect 14096 2382 14148 2388
rect 14200 1970 14228 3538
rect 14476 3466 14504 4422
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 14292 1737 14320 2246
rect 14278 1728 14334 1737
rect 14278 1663 14334 1672
rect 14384 1578 14412 2994
rect 14476 2514 14504 3402
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14568 3097 14596 3130
rect 14554 3088 14610 3097
rect 14660 3058 14688 5510
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14554 3023 14610 3032
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14752 1986 14780 3878
rect 14844 2446 14872 4966
rect 15028 2774 15056 11562
rect 15120 11354 15148 34682
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15212 30258 15240 32166
rect 15384 30388 15436 30394
rect 15384 30330 15436 30336
rect 15396 30258 15424 30330
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15384 30252 15436 30258
rect 15384 30194 15436 30200
rect 15396 29850 15424 30194
rect 15476 30184 15528 30190
rect 15476 30126 15528 30132
rect 15488 30054 15516 30126
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 15396 29170 15424 29786
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15488 25770 15516 27270
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 15488 25362 15516 25706
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15212 17882 15240 20402
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15580 6458 15608 13806
rect 15764 9382 15792 35022
rect 15948 33862 15976 35634
rect 15936 33856 15988 33862
rect 15936 33798 15988 33804
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15856 26790 15884 26930
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15856 26586 15884 26726
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15856 20466 15884 26522
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15856 14074 15884 14418
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15948 14006 15976 33798
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 3058 15148 6054
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15382 3224 15438 3233
rect 15382 3159 15384 3168
rect 15436 3159 15438 3168
rect 15384 3130 15436 3136
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 14936 2746 15056 2774
rect 14936 2582 14964 2746
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14292 1550 14412 1578
rect 14568 1958 14780 1986
rect 14292 800 14320 1550
rect 14568 800 14596 1958
rect 14844 800 14872 2382
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15028 1873 15056 2246
rect 15014 1864 15070 1873
rect 15014 1799 15070 1808
rect 15120 800 15148 2994
rect 15488 2258 15516 4422
rect 15580 4078 15608 6394
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15672 2446 15700 5510
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15764 3126 15792 4966
rect 15856 4010 15884 6258
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15856 3602 15884 3946
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15948 3194 15976 9522
rect 16040 6866 16068 37266
rect 16224 36378 16252 39200
rect 16592 36378 16620 39200
rect 16960 36854 16988 39200
rect 17236 36922 17264 39200
rect 17408 37324 17460 37330
rect 17408 37266 17460 37272
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 16948 36848 17000 36854
rect 16948 36790 17000 36796
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 16212 36372 16264 36378
rect 16212 36314 16264 36320
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16684 35834 16712 36722
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16868 35834 16896 36110
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16132 5914 16160 14010
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16316 11354 16344 12242
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16224 7206 16252 7346
rect 16500 7206 16528 8502
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16224 7018 16252 7142
rect 16224 6990 16344 7018
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16132 4146 16160 5850
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3534 16160 3878
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15396 2230 15516 2258
rect 15396 800 15424 2230
rect 15672 800 15700 2382
rect 15948 800 15976 2926
rect 16132 1766 16160 3470
rect 16120 1760 16172 1766
rect 16120 1702 16172 1708
rect 16224 800 16252 4422
rect 16316 3602 16344 6990
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16500 6322 16528 6666
rect 16592 6390 16620 26862
rect 16684 11898 16712 35566
rect 16776 34950 16804 35634
rect 16764 34944 16816 34950
rect 16764 34886 16816 34892
rect 16776 26926 16804 34886
rect 16960 34746 16988 36790
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 17132 36168 17184 36174
rect 17132 36110 17184 36116
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 17144 33862 17172 36110
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16776 19854 16804 23462
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 17144 15162 17172 33798
rect 17236 22506 17264 36518
rect 17224 22500 17276 22506
rect 17224 22442 17276 22448
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16684 11082 16712 11154
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16408 4622 16436 5034
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16500 2446 16528 4966
rect 16960 3738 16988 14962
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16854 3632 16910 3641
rect 16854 3567 16910 3576
rect 16868 3194 16896 3567
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16500 800 16528 2382
rect 16776 800 16804 2926
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 1834 16896 2246
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 17052 800 17080 3878
rect 17144 3670 17172 13874
rect 17420 10198 17448 37266
rect 17500 37188 17552 37194
rect 17500 37130 17552 37136
rect 17512 35290 17540 37130
rect 17604 36378 17632 39200
rect 17972 37262 18000 39200
rect 17960 37256 18012 37262
rect 17960 37198 18012 37204
rect 17592 36372 17644 36378
rect 17592 36314 17644 36320
rect 17868 35692 17920 35698
rect 17868 35634 17920 35640
rect 17880 35494 17908 35634
rect 17868 35488 17920 35494
rect 17868 35430 17920 35436
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17512 29850 17540 30126
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17604 26858 17632 28358
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17604 23322 17632 26794
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17696 19718 17724 23122
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17696 17270 17724 18226
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17696 16590 17724 17206
rect 17788 17202 17816 19314
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 16658 17816 17138
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17420 9722 17448 10134
rect 17512 9926 17540 10406
rect 17880 10266 17908 35430
rect 17972 35290 18000 37198
rect 18340 36922 18368 39200
rect 18328 36916 18380 36922
rect 18328 36858 18380 36864
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 18064 36650 18092 36722
rect 18052 36644 18104 36650
rect 18052 36586 18104 36592
rect 18604 36644 18656 36650
rect 18604 36586 18656 36592
rect 18052 36168 18104 36174
rect 18052 36110 18104 36116
rect 18064 36038 18092 36110
rect 18052 36032 18104 36038
rect 18052 35974 18104 35980
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18064 34202 18092 35974
rect 18616 35290 18644 36586
rect 18708 35834 18736 39200
rect 18880 37324 18932 37330
rect 18880 37266 18932 37272
rect 18892 35894 18920 37266
rect 19076 37262 19104 39200
rect 19064 37256 19116 37262
rect 19064 37198 19116 37204
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 18892 35866 19012 35894
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18604 35284 18656 35290
rect 18604 35226 18656 35232
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 18340 33658 18368 34546
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18788 32292 18840 32298
rect 18788 32234 18840 32240
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 18328 30116 18380 30122
rect 18328 30058 18380 30064
rect 18340 28694 18368 30058
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 18432 28558 18460 29990
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 27470 18460 28358
rect 18708 27606 18736 30194
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18064 23322 18092 23666
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17972 22098 18000 23054
rect 17960 22092 18012 22098
rect 18800 22094 18828 32234
rect 17960 22034 18012 22040
rect 18616 22066 18828 22094
rect 17972 20058 18000 22034
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17972 18426 18000 19790
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18064 18290 18092 18566
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15570 18552 15846
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18420 14340 18472 14346
rect 18420 14282 18472 14288
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 7002 17264 7278
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17236 3058 17264 4966
rect 17512 4554 17540 9862
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17696 6118 17724 6258
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17500 4548 17552 4554
rect 17500 4490 17552 4496
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17328 3534 17356 3946
rect 17512 3602 17540 4490
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17512 3369 17540 3538
rect 17498 3360 17554 3369
rect 17498 3295 17554 3304
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17604 2446 17632 4422
rect 17696 3194 17724 6054
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17328 800 17356 2382
rect 17696 2258 17724 2994
rect 17604 2230 17724 2258
rect 17604 800 17632 2230
rect 17880 800 17908 3334
rect 17972 3126 18000 13942
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18064 3058 18092 4422
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18156 2378 18184 3878
rect 18248 2922 18276 12038
rect 18432 5914 18460 14282
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18340 3058 18368 4966
rect 18432 3534 18460 5850
rect 18524 4593 18552 9862
rect 18510 4584 18566 4593
rect 18510 4519 18566 4528
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18616 3194 18644 22066
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18708 16114 18736 16662
rect 18892 16114 18920 18566
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 18156 800 18184 2314
rect 18432 800 18460 2314
rect 18708 800 18736 2790
rect 18800 2582 18828 15370
rect 18984 10674 19012 35866
rect 19260 35290 19288 37198
rect 19352 36922 19380 39200
rect 19720 39114 19748 39200
rect 19812 39114 19840 39222
rect 19720 39086 19840 39114
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36922 20024 39222
rect 20074 39200 20130 40000
rect 20442 39200 20498 40000
rect 20810 39200 20866 40000
rect 21086 39200 21142 40000
rect 21454 39200 21510 40000
rect 21822 39200 21878 40000
rect 22190 39200 22246 40000
rect 22558 39200 22614 40000
rect 22926 39200 22982 40000
rect 23202 39200 23258 40000
rect 23570 39200 23626 40000
rect 23938 39200 23994 40000
rect 24306 39200 24362 40000
rect 24674 39200 24730 40000
rect 24950 39200 25006 40000
rect 25318 39200 25374 40000
rect 25686 39200 25742 40000
rect 26054 39200 26110 40000
rect 26422 39200 26478 40000
rect 26790 39200 26846 40000
rect 27066 39200 27122 40000
rect 27172 39222 27384 39250
rect 20088 37262 20116 39200
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19340 36372 19392 36378
rect 19340 36314 19392 36320
rect 19352 35834 19380 36314
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19444 34950 19472 36722
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19996 35494 20024 36110
rect 19984 35488 20036 35494
rect 19984 35430 20036 35436
rect 19432 34944 19484 34950
rect 19432 34886 19484 34892
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34678 20024 35430
rect 20088 35290 20116 37198
rect 20456 37126 20484 39200
rect 20168 37120 20220 37126
rect 20168 37062 20220 37068
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 20444 37120 20496 37126
rect 20444 37062 20496 37068
rect 20180 36961 20208 37062
rect 20166 36952 20222 36961
rect 20166 36887 20222 36896
rect 20168 36780 20220 36786
rect 20168 36722 20220 36728
rect 20076 35284 20128 35290
rect 20076 35226 20128 35232
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 20180 34626 20208 36722
rect 20260 36100 20312 36106
rect 20260 36042 20312 36048
rect 20272 34746 20300 36042
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 19076 11898 19104 34614
rect 20180 34598 20300 34626
rect 20272 34542 20300 34598
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19444 33454 19472 34342
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19340 33380 19392 33386
rect 19340 33322 19392 33328
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 19260 32910 19288 33254
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19260 30326 19288 32846
rect 19352 32774 19380 33322
rect 19444 32910 19472 33390
rect 19536 33114 19564 33458
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19444 30326 19472 32846
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19444 30190 19472 30262
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19444 30054 19472 30126
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 25158 20024 32710
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20180 29850 20208 30194
rect 20168 29844 20220 29850
rect 20168 29786 20220 29792
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19444 23526 19472 24074
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19168 11558 19196 11834
rect 19352 11694 19380 12106
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19352 11286 19380 11630
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 18984 3534 19012 4966
rect 19064 4072 19116 4078
rect 19062 4040 19064 4049
rect 19116 4040 19118 4049
rect 19062 3975 19118 3984
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18984 800 19012 2926
rect 19168 2378 19196 4966
rect 19352 4758 19380 11018
rect 19444 11014 19472 23462
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19514 20024 19858
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19812 18698 19840 19314
rect 19904 18970 19932 19382
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19996 18698 20024 19450
rect 20168 19236 20220 19242
rect 20168 19178 20220 19184
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 20180 16114 20208 19178
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20180 15706 20208 16050
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 20272 14822 20300 34478
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19812 12170 19840 12582
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20364 11150 20392 37062
rect 20824 36922 20852 39200
rect 21100 37262 21128 39200
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 21088 37256 21140 37262
rect 21088 37198 21140 37204
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20444 36780 20496 36786
rect 20444 36722 20496 36728
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20456 35018 20484 36722
rect 20548 36378 20576 36722
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20732 35494 20760 36110
rect 20916 35834 20944 37198
rect 21468 36922 21496 39200
rect 21456 36916 21508 36922
rect 21456 36858 21508 36864
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21008 36378 21036 36722
rect 21836 36378 21864 39200
rect 22204 37194 22232 39200
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 20996 36372 21048 36378
rect 20996 36314 21048 36320
rect 21824 36372 21876 36378
rect 21824 36314 21876 36320
rect 21916 36168 21968 36174
rect 21916 36110 21968 36116
rect 20904 35828 20956 35834
rect 20904 35770 20956 35776
rect 21928 35494 21956 36110
rect 22204 35834 22232 37130
rect 22572 36922 22600 39200
rect 22652 37324 22704 37330
rect 22652 37266 22704 37272
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22560 36780 22612 36786
rect 22560 36722 22612 36728
rect 22192 35828 22244 35834
rect 22192 35770 22244 35776
rect 22572 35562 22600 36722
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 21916 35488 21968 35494
rect 21916 35430 21968 35436
rect 20444 35012 20496 35018
rect 20444 34954 20496 34960
rect 20536 34944 20588 34950
rect 20536 34886 20588 34892
rect 20548 22778 20576 34886
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20640 23050 20668 23530
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20640 22710 20668 22986
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20640 19378 20668 21966
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11762 20484 12038
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20180 8498 20208 8774
rect 20364 8566 20392 8910
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19352 3738 19380 4082
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 19260 800 19288 3470
rect 19444 3058 19472 6598
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19904 3913 19932 4014
rect 19890 3904 19946 3913
rect 19890 3839 19946 3848
rect 19904 3738 19932 3839
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3194 20024 6666
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20088 4622 20116 5510
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19352 1698 19380 2246
rect 19340 1692 19392 1698
rect 19340 1634 19392 1640
rect 19444 1170 19472 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 1986 20024 2926
rect 19812 1958 20024 1986
rect 19444 1142 19564 1170
rect 19536 800 19564 1142
rect 19812 800 19840 1958
rect 20088 800 20116 4558
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 3058 20208 4422
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20272 2446 20300 8298
rect 20364 7750 20392 8502
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20364 6474 20392 7686
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20456 6662 20484 7278
rect 20548 7274 20576 12922
rect 20732 12442 20760 35430
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 20916 24410 20944 24754
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 21008 22030 21036 22374
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 21100 10538 21128 34886
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21284 22098 21312 23054
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21928 15094 21956 35430
rect 22192 34944 22244 34950
rect 22192 34886 22244 34892
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22112 25498 22140 25842
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 22020 23050 22048 25162
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22020 22642 22048 22986
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 22020 11830 22048 12038
rect 22204 11898 22232 34886
rect 22376 34400 22428 34406
rect 22374 34368 22376 34377
rect 22428 34368 22430 34377
rect 22374 34303 22430 34312
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22296 30190 22324 30534
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22296 29646 22324 29990
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22388 17882 22416 18702
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22282 13288 22338 13297
rect 22282 13223 22284 13232
rect 22336 13223 22338 13232
rect 22284 13194 22336 13200
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22296 11082 22324 11698
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21008 8906 21036 9046
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 8634 21220 8774
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20548 6934 20576 7210
rect 20536 6928 20588 6934
rect 20536 6870 20588 6876
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20364 6446 20484 6474
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 3534 20392 4966
rect 20456 4162 20484 6446
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4282 20576 4422
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20456 4134 20576 4162
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20364 2990 20392 3470
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20364 800 20392 2790
rect 20456 1601 20484 4014
rect 20548 3738 20576 4134
rect 20640 4049 20668 6598
rect 20626 4040 20682 4049
rect 20626 3975 20682 3984
rect 20732 3738 20760 8298
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6798 20852 7142
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 20916 4622 20944 5510
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20810 4448 20866 4457
rect 20810 4383 20866 4392
rect 20824 4010 20852 4383
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 2774 20668 3470
rect 20548 2746 20668 2774
rect 20548 2122 20576 2746
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 2281 20668 2314
rect 20626 2272 20682 2281
rect 20626 2207 20682 2216
rect 20548 2094 20668 2122
rect 20442 1592 20498 1601
rect 20442 1527 20498 1536
rect 20640 800 20668 2094
rect 20916 800 20944 4558
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21008 4282 21036 4490
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21008 3058 21036 3946
rect 21192 3534 21220 4966
rect 21468 4622 21496 4966
rect 22112 4622 22140 5510
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21192 800 21220 2790
rect 21468 800 21496 4558
rect 21744 800 21772 4558
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21928 3602 21956 4218
rect 22098 4176 22154 4185
rect 22098 4111 22154 4120
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21928 2650 21956 3538
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 22020 800 22048 3878
rect 22112 3602 22140 4111
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22204 3534 22232 4694
rect 22296 4146 22324 5714
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22112 1970 22140 2994
rect 22388 2774 22416 4966
rect 22480 4690 22508 14350
rect 22572 13530 22600 14962
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22664 12442 22692 37266
rect 22836 36848 22888 36854
rect 22836 36790 22888 36796
rect 22848 36310 22876 36790
rect 22836 36304 22888 36310
rect 22836 36246 22888 36252
rect 22940 35834 22968 39200
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 22928 35828 22980 35834
rect 22928 35770 22980 35776
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22848 34950 22876 35634
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22744 30660 22796 30666
rect 22744 30602 22796 30608
rect 22756 30394 22784 30602
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22940 29306 22968 30194
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 23032 26234 23060 37062
rect 23216 36786 23244 39200
rect 23584 36922 23612 39200
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23112 36100 23164 36106
rect 23112 36042 23164 36048
rect 23124 34678 23152 36042
rect 23204 36032 23256 36038
rect 23204 35974 23256 35980
rect 23112 34672 23164 34678
rect 23112 34614 23164 34620
rect 22940 26206 23060 26234
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22848 19310 22876 19654
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22848 18766 22876 19246
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22940 9518 22968 26206
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23124 25294 23152 25638
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23124 19378 23152 19790
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23124 18970 23152 19314
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23216 15162 23244 35974
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23308 24206 23336 25230
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23308 22098 23336 24142
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23308 21622 23336 22034
rect 23296 21616 23348 21622
rect 23296 21558 23348 21564
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 23308 18766 23336 19926
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23216 14482 23244 15098
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23202 13288 23258 13297
rect 23202 13223 23204 13232
rect 23256 13223 23258 13232
rect 23204 13194 23256 13200
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23124 11286 23152 13126
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 23400 8838 23428 36518
rect 23492 35834 23520 36722
rect 23768 36378 23796 36722
rect 23952 36378 23980 39200
rect 24320 37262 24348 39200
rect 24308 37256 24360 37262
rect 24308 37198 24360 37204
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23848 36032 23900 36038
rect 23848 35974 23900 35980
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23676 22094 23704 35974
rect 23860 34746 23888 35974
rect 24320 35834 24348 37198
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24308 35828 24360 35834
rect 24308 35770 24360 35776
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 23940 34468 23992 34474
rect 23940 34410 23992 34416
rect 23952 33862 23980 34410
rect 23940 33856 23992 33862
rect 23940 33798 23992 33804
rect 23952 22094 23980 33798
rect 23584 22066 23704 22094
rect 23768 22066 23980 22094
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 17678 23520 18566
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23584 13938 23612 22066
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23676 20058 23704 21490
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23676 19446 23704 19994
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23662 14920 23718 14929
rect 23662 14855 23664 14864
rect 23716 14855 23718 14864
rect 23664 14826 23716 14832
rect 23676 14414 23704 14826
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23584 13530 23612 13874
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23584 13002 23612 13262
rect 23492 12986 23612 13002
rect 23676 12986 23704 13330
rect 23480 12980 23612 12986
rect 23532 12974 23612 12980
rect 23664 12980 23716 12986
rect 23480 12922 23532 12928
rect 23664 12922 23716 12928
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23478 8392 23534 8401
rect 23478 8327 23480 8336
rect 23532 8327 23534 8336
rect 23480 8298 23532 8304
rect 23204 6928 23256 6934
rect 23768 6914 23796 22066
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24136 14006 24164 14350
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24320 14006 24348 14214
rect 24124 14000 24176 14006
rect 24308 14000 24360 14006
rect 24124 13942 24176 13948
rect 24306 13968 24308 13977
rect 24360 13968 24362 13977
rect 24306 13903 24362 13912
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 23860 12170 23888 12922
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 24596 11830 24624 37062
rect 24688 36938 24716 39200
rect 24964 36938 24992 39200
rect 25332 37262 25360 39200
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25504 37256 25556 37262
rect 25504 37198 25556 37204
rect 24688 36922 24900 36938
rect 24964 36922 25084 36938
rect 24688 36916 24912 36922
rect 24688 36910 24860 36916
rect 24964 36916 25096 36922
rect 24964 36910 25044 36916
rect 24860 36858 24912 36864
rect 25044 36858 25096 36864
rect 25332 36378 25360 37198
rect 25412 36780 25464 36786
rect 25412 36722 25464 36728
rect 25320 36372 25372 36378
rect 25320 36314 25372 36320
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24872 35494 24900 36110
rect 24952 35556 25004 35562
rect 24952 35498 25004 35504
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24872 14550 24900 35430
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24412 9518 24440 10678
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24676 9444 24728 9450
rect 24676 9386 24728 9392
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23204 6870 23256 6876
rect 23584 6886 23796 6914
rect 22650 5400 22706 5409
rect 22650 5335 22706 5344
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22572 2990 22600 4966
rect 22664 4078 22692 5335
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22756 3534 22784 4422
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22296 2746 22416 2774
rect 22296 2446 22324 2746
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 22296 800 22324 2382
rect 22572 800 22600 2926
rect 22848 800 22876 3878
rect 22940 3584 22968 4422
rect 23216 4146 23244 6870
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23032 3913 23060 4082
rect 23018 3904 23074 3913
rect 23018 3839 23074 3848
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23400 3641 23428 3674
rect 23386 3632 23442 3641
rect 23020 3596 23072 3602
rect 22940 3556 23020 3584
rect 23386 3567 23442 3576
rect 23020 3538 23072 3544
rect 23032 1902 23060 3538
rect 23294 3496 23350 3505
rect 23294 3431 23350 3440
rect 23308 3398 23336 3431
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23020 1896 23072 1902
rect 23020 1838 23072 1844
rect 23124 800 23152 2994
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23400 800 23428 2926
rect 23584 2650 23612 6886
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23676 800 23704 3878
rect 23768 3058 23796 4422
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23860 2650 23888 8910
rect 24688 8838 24716 9386
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24872 7886 24900 8570
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24964 6866 24992 35498
rect 25424 35494 25452 36722
rect 25412 35488 25464 35494
rect 25412 35430 25464 35436
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25332 32230 25360 32370
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25240 29170 25268 29514
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25240 28082 25268 29106
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25332 26234 25360 32166
rect 25240 26206 25360 26234
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 22642 25176 24006
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25240 22094 25268 26206
rect 25240 22066 25360 22094
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25056 8974 25084 9454
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 25056 6730 25084 7482
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24032 5840 24084 5846
rect 24032 5782 24084 5788
rect 23938 4312 23994 4321
rect 23938 4247 23994 4256
rect 23952 3738 23980 4247
rect 24044 4146 24072 5782
rect 24872 5642 24900 6666
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24044 3194 24072 3674
rect 24228 3466 24256 4966
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23940 1828 23992 1834
rect 23940 1770 23992 1776
rect 23952 800 23980 1770
rect 24228 800 24256 3402
rect 24412 2446 24440 4966
rect 24504 3058 24532 5510
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 25056 4622 25084 4966
rect 25148 4826 25176 9522
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25240 8634 25268 8842
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25240 5574 25268 8434
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24596 4282 24624 4422
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 24596 4078 24624 4218
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24766 3496 24822 3505
rect 24766 3431 24768 3440
rect 24820 3431 24822 3440
rect 24768 3402 24820 3408
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24492 2916 24544 2922
rect 24492 2858 24544 2864
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24412 1834 24440 2382
rect 24400 1828 24452 1834
rect 24400 1770 24452 1776
rect 24504 800 24532 2858
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24780 800 24808 2314
rect 24872 2009 24900 2314
rect 24858 2000 24914 2009
rect 24858 1935 24914 1944
rect 25056 800 25084 4558
rect 25332 4162 25360 22066
rect 25424 14006 25452 35430
rect 25516 35154 25544 37198
rect 25700 37126 25728 39200
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 25688 37120 25740 37126
rect 25688 37062 25740 37068
rect 25504 35148 25556 35154
rect 25504 35090 25556 35096
rect 25504 34536 25556 34542
rect 25504 34478 25556 34484
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25516 12434 25544 34478
rect 25608 22094 25636 37062
rect 26068 36666 26096 39200
rect 26240 36916 26292 36922
rect 26240 36858 26292 36864
rect 26252 36666 26280 36858
rect 26436 36786 26464 39200
rect 26804 37126 26832 39200
rect 27080 39114 27108 39200
rect 27172 39114 27200 39222
rect 27080 39086 27200 39114
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 26792 37120 26844 37126
rect 26792 37062 26844 37068
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 26884 36780 26936 36786
rect 26884 36722 26936 36728
rect 26068 36638 26280 36666
rect 26240 36576 26292 36582
rect 26240 36518 26292 36524
rect 26252 36310 26280 36518
rect 26436 36378 26464 36722
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26240 36304 26292 36310
rect 26240 36246 26292 36252
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26160 32570 26188 35634
rect 26240 35012 26292 35018
rect 26240 34954 26292 34960
rect 26252 34678 26280 34954
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 26240 34672 26292 34678
rect 26240 34614 26292 34620
rect 26148 32564 26200 32570
rect 26148 32506 26200 32512
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 26252 31890 26280 32370
rect 26240 31884 26292 31890
rect 26240 31826 26292 31832
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25700 24410 25728 25094
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25700 24206 25728 24346
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25608 22066 25728 22094
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25608 19922 25636 20266
rect 25596 19916 25648 19922
rect 25596 19858 25648 19864
rect 25608 18970 25636 19858
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25424 12406 25544 12434
rect 25424 9450 25452 12406
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25608 8498 25636 11154
rect 25700 10062 25728 22066
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25792 15502 25820 17478
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25884 8378 25912 31758
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 26160 27606 26188 28018
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26252 27470 26280 28018
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 26068 22778 26096 22986
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26252 19378 26280 19654
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26252 18766 26280 19110
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 26068 15434 26096 18566
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26344 14074 26372 34886
rect 26620 32026 26648 36110
rect 26896 35698 26924 36722
rect 26988 35834 27016 37198
rect 27080 36378 27108 37198
rect 27356 36922 27384 39222
rect 27434 39200 27490 40000
rect 27802 39200 27858 40000
rect 28170 39200 28226 40000
rect 28538 39200 28594 40000
rect 28814 39200 28870 40000
rect 29182 39200 29238 40000
rect 29550 39200 29606 40000
rect 29918 39200 29974 40000
rect 30286 39200 30342 40000
rect 30562 39200 30618 40000
rect 30930 39200 30986 40000
rect 31298 39200 31354 40000
rect 31666 39200 31722 40000
rect 32034 39200 32090 40000
rect 32402 39200 32458 40000
rect 32678 39200 32734 40000
rect 33046 39200 33102 40000
rect 33414 39200 33470 40000
rect 33782 39200 33838 40000
rect 34150 39200 34206 40000
rect 34426 39200 34482 40000
rect 34794 39200 34850 40000
rect 35162 39200 35218 40000
rect 35530 39200 35586 40000
rect 35898 39200 35954 40000
rect 36266 39200 36322 40000
rect 36542 39200 36598 40000
rect 36910 39200 36966 40000
rect 37016 39222 37228 39250
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27264 36378 27292 36722
rect 27068 36372 27120 36378
rect 27068 36314 27120 36320
rect 27252 36372 27304 36378
rect 27252 36314 27304 36320
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 26976 35828 27028 35834
rect 26976 35770 27028 35776
rect 26884 35692 26936 35698
rect 26884 35634 26936 35640
rect 26608 32020 26660 32026
rect 26608 31962 26660 31968
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 26436 28082 26464 28358
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26436 26042 26464 28018
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 26436 25158 26464 25978
rect 26424 25152 26476 25158
rect 26424 25094 26476 25100
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26436 19514 26464 22374
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26436 18902 26464 19450
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 25516 8350 25912 8378
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25240 4134 25360 4162
rect 25240 1737 25268 4134
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 25332 3534 25360 4014
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25424 3058 25452 5510
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25226 1728 25282 1737
rect 25226 1663 25282 1672
rect 25332 800 25360 2790
rect 25516 1873 25544 8350
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25700 5710 25728 6190
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 25596 3392 25648 3398
rect 25594 3360 25596 3369
rect 25648 3360 25650 3369
rect 25594 3295 25650 3304
rect 25792 2854 25820 3878
rect 25884 3058 25912 7686
rect 25976 4690 26004 10542
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26344 8362 26372 8774
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 25964 4276 26016 4282
rect 25964 4218 26016 4224
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25780 2848 25832 2854
rect 25608 2796 25780 2802
rect 25608 2790 25832 2796
rect 25608 2774 25820 2790
rect 25976 2774 26004 4218
rect 26068 4010 26096 5306
rect 26344 4622 26372 8298
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26344 4486 26372 4558
rect 26332 4480 26384 4486
rect 26332 4422 26384 4428
rect 26056 4004 26108 4010
rect 26056 3946 26108 3952
rect 26240 3664 26292 3670
rect 26240 3606 26292 3612
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 25502 1864 25558 1873
rect 25502 1799 25558 1808
rect 25608 800 25636 2774
rect 25884 2746 26004 2774
rect 26068 2774 26096 3334
rect 26252 2938 26280 3606
rect 26436 3602 26464 5510
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26528 3534 26556 5510
rect 26620 5370 26648 17274
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26712 5114 26740 31758
rect 27080 30938 27108 36110
rect 27448 35766 27476 39200
rect 27816 37126 27844 39200
rect 27804 37120 27856 37126
rect 27804 37062 27856 37068
rect 28184 36922 28212 39200
rect 28448 37392 28500 37398
rect 28448 37334 28500 37340
rect 28172 36916 28224 36922
rect 28172 36858 28224 36864
rect 28172 36712 28224 36718
rect 28172 36654 28224 36660
rect 28184 36378 28212 36654
rect 28172 36372 28224 36378
rect 28172 36314 28224 36320
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 27908 36106 27936 36246
rect 27896 36100 27948 36106
rect 27896 36042 27948 36048
rect 28460 36038 28488 37334
rect 28552 37262 28580 39200
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28644 36378 28672 36722
rect 28632 36372 28684 36378
rect 28632 36314 28684 36320
rect 28448 36032 28500 36038
rect 28448 35974 28500 35980
rect 28736 35894 28764 37062
rect 28644 35866 28764 35894
rect 27436 35760 27488 35766
rect 27436 35702 27488 35708
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 27172 34746 27200 35634
rect 28172 35488 28224 35494
rect 28172 35430 28224 35436
rect 28184 35222 28212 35430
rect 28172 35216 28224 35222
rect 28172 35158 28224 35164
rect 28448 35148 28500 35154
rect 28448 35090 28500 35096
rect 27160 34740 27212 34746
rect 27160 34682 27212 34688
rect 27528 34672 27580 34678
rect 27528 34614 27580 34620
rect 27540 33522 27568 34614
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27816 32910 27844 33390
rect 28460 33046 28488 35090
rect 28448 33040 28500 33046
rect 28448 32982 28500 32988
rect 27804 32904 27856 32910
rect 27804 32846 27856 32852
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27068 30932 27120 30938
rect 27068 30874 27120 30880
rect 27540 30870 27568 31826
rect 28460 31822 28488 32982
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 27528 30864 27580 30870
rect 27528 30806 27580 30812
rect 27160 30660 27212 30666
rect 27160 30602 27212 30608
rect 27172 28082 27200 30602
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 27080 27470 27108 27814
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27172 25974 27200 28018
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27264 22574 27292 22918
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27264 19990 27292 22510
rect 27252 19984 27304 19990
rect 27252 19926 27304 19932
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27172 19446 27200 19790
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27264 19446 27292 19654
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27252 19440 27304 19446
rect 27252 19382 27304 19388
rect 27264 15706 27292 19382
rect 27252 15700 27304 15706
rect 27252 15642 27304 15648
rect 27068 11620 27120 11626
rect 27068 11562 27120 11568
rect 27080 11354 27108 11562
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26896 5574 26924 9590
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26620 5086 26740 5114
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26252 2922 26464 2938
rect 26252 2916 26476 2922
rect 26252 2910 26424 2916
rect 26424 2858 26476 2864
rect 26068 2746 26188 2774
rect 25780 2576 25832 2582
rect 25780 2518 25832 2524
rect 25792 2310 25820 2518
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25884 800 25912 2746
rect 26160 800 26188 2746
rect 26620 1902 26648 5086
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26712 2378 26740 4966
rect 26792 4548 26844 4554
rect 26792 4490 26844 4496
rect 26804 3466 26832 4490
rect 26988 4010 27016 8842
rect 27252 4752 27304 4758
rect 27252 4694 27304 4700
rect 27068 4684 27120 4690
rect 27068 4626 27120 4632
rect 27080 4214 27108 4626
rect 27160 4548 27212 4554
rect 27160 4490 27212 4496
rect 27068 4208 27120 4214
rect 27068 4150 27120 4156
rect 26976 4004 27028 4010
rect 26976 3946 27028 3952
rect 26792 3460 26844 3466
rect 26792 3402 26844 3408
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26700 2372 26752 2378
rect 26700 2314 26752 2320
rect 26608 1896 26660 1902
rect 26608 1838 26660 1844
rect 26424 1692 26476 1698
rect 26424 1634 26476 1640
rect 26436 800 26464 1634
rect 26712 800 26740 2314
rect 26896 800 26924 3334
rect 27172 2310 27200 4490
rect 27264 2446 27292 4694
rect 27356 3097 27384 30534
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 27448 27674 27476 28018
rect 27436 27668 27488 27674
rect 27436 27610 27488 27616
rect 28172 25152 28224 25158
rect 28172 25094 28224 25100
rect 28184 24818 28212 25094
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 20330 28304 23054
rect 28264 20324 28316 20330
rect 28264 20266 28316 20272
rect 28276 19174 28304 20266
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28276 15502 28304 19110
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28540 14884 28592 14890
rect 28540 14826 28592 14832
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 27540 11898 27568 12786
rect 28356 12096 28408 12102
rect 28356 12038 28408 12044
rect 27528 11892 27580 11898
rect 27528 11834 27580 11840
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 27816 10810 27844 11222
rect 28000 11218 28028 11766
rect 28368 11626 28396 12038
rect 28356 11620 28408 11626
rect 28356 11562 28408 11568
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 28460 10062 28488 11494
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 27436 5160 27488 5166
rect 27436 5102 27488 5108
rect 27448 4486 27476 5102
rect 27632 5098 27660 7210
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27620 5092 27672 5098
rect 27620 5034 27672 5040
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27436 4480 27488 4486
rect 27436 4422 27488 4428
rect 27540 4146 27568 4966
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27632 4282 27660 4558
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27816 3534 27844 7142
rect 28552 6914 28580 14826
rect 28644 7546 28672 35866
rect 28828 35834 28856 39200
rect 29092 37460 29144 37466
rect 29092 37402 29144 37408
rect 28908 37256 28960 37262
rect 28908 37198 28960 37204
rect 28920 36378 28948 37198
rect 28908 36372 28960 36378
rect 28908 36314 28960 36320
rect 29000 36236 29052 36242
rect 29000 36178 29052 36184
rect 29012 36145 29040 36178
rect 28998 36136 29054 36145
rect 28998 36071 29054 36080
rect 28908 36032 28960 36038
rect 28908 35974 28960 35980
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 28920 26234 28948 35974
rect 29104 35894 29132 37402
rect 29196 36922 29224 39200
rect 29460 37256 29512 37262
rect 29460 37198 29512 37204
rect 29564 37210 29592 39200
rect 29184 36916 29236 36922
rect 29184 36858 29236 36864
rect 29368 36780 29420 36786
rect 29368 36722 29420 36728
rect 29104 35866 29316 35894
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 29196 32026 29224 33458
rect 29184 32020 29236 32026
rect 29184 31962 29236 31968
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 28736 26206 28948 26234
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28460 6886 28580 6914
rect 27988 5024 28040 5030
rect 27988 4966 28040 4972
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27342 3088 27398 3097
rect 27342 3023 27398 3032
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 27342 2408 27398 2417
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 27172 800 27200 2246
rect 27264 1698 27292 2382
rect 27342 2343 27344 2352
rect 27396 2343 27398 2352
rect 27344 2314 27396 2320
rect 27252 1692 27304 1698
rect 27252 1634 27304 1640
rect 27448 800 27476 2994
rect 27526 2952 27582 2961
rect 27526 2887 27528 2896
rect 27580 2887 27582 2896
rect 27528 2858 27580 2864
rect 27724 800 27752 3334
rect 28000 3058 28028 4966
rect 28092 3058 28120 4966
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28172 3392 28224 3398
rect 28172 3334 28224 3340
rect 28184 3126 28212 3334
rect 28172 3120 28224 3126
rect 28172 3062 28224 3068
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28092 2938 28120 2994
rect 28000 2910 28120 2938
rect 28000 800 28028 2910
rect 28078 2544 28134 2553
rect 28078 2479 28134 2488
rect 28092 2446 28120 2479
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28276 800 28304 4218
rect 28356 3664 28408 3670
rect 28356 3606 28408 3612
rect 28368 3126 28396 3606
rect 28356 3120 28408 3126
rect 28356 3062 28408 3068
rect 28460 1630 28488 6886
rect 28736 6866 28764 26206
rect 29012 25226 29040 28426
rect 29000 25220 29052 25226
rect 29000 25162 29052 25168
rect 29012 20534 29040 25162
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29012 15162 29040 16050
rect 29184 15496 29236 15502
rect 29184 15438 29236 15444
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 29196 15094 29224 15438
rect 29184 15088 29236 15094
rect 29184 15030 29236 15036
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 29012 12918 29040 14418
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 29012 9586 29040 11494
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 28814 7848 28870 7857
rect 28814 7783 28870 7792
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28644 4146 28672 6598
rect 28724 4548 28776 4554
rect 28724 4490 28776 4496
rect 28736 4457 28764 4490
rect 28722 4448 28778 4457
rect 28722 4383 28778 4392
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 28448 1624 28500 1630
rect 28448 1566 28500 1572
rect 28552 800 28580 3878
rect 28828 3126 28856 7783
rect 28908 6996 28960 7002
rect 28908 6938 28960 6944
rect 28920 3126 28948 6938
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28920 2774 28948 2926
rect 28828 2746 28948 2774
rect 28724 2304 28776 2310
rect 28724 2246 28776 2252
rect 28736 1970 28764 2246
rect 28724 1964 28776 1970
rect 28724 1906 28776 1912
rect 28828 800 28856 2746
rect 29012 2446 29040 3878
rect 29104 2990 29132 5510
rect 29288 5370 29316 35866
rect 29380 33658 29408 36722
rect 29472 35562 29500 37198
rect 29564 37194 29684 37210
rect 29564 37188 29696 37194
rect 29564 37182 29644 37188
rect 29644 37130 29696 37136
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 29552 36168 29604 36174
rect 29552 36110 29604 36116
rect 29460 35556 29512 35562
rect 29460 35498 29512 35504
rect 29564 35290 29592 36110
rect 29748 35834 29776 37062
rect 29932 36922 29960 39200
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 30102 36408 30158 36417
rect 30102 36343 30158 36352
rect 30116 36038 30144 36343
rect 30194 36272 30250 36281
rect 30194 36207 30250 36216
rect 30208 36174 30236 36207
rect 30196 36168 30248 36174
rect 30196 36110 30248 36116
rect 30104 36032 30156 36038
rect 30104 35974 30156 35980
rect 30300 35834 30328 39200
rect 30576 37262 30604 39200
rect 30656 37324 30708 37330
rect 30656 37266 30708 37272
rect 30564 37256 30616 37262
rect 30564 37198 30616 37204
rect 30472 36100 30524 36106
rect 30472 36042 30524 36048
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 30288 35828 30340 35834
rect 30288 35770 30340 35776
rect 29644 35488 29696 35494
rect 29644 35430 29696 35436
rect 29552 35284 29604 35290
rect 29552 35226 29604 35232
rect 29656 35086 29684 35430
rect 29644 35080 29696 35086
rect 29644 35022 29696 35028
rect 29920 34944 29972 34950
rect 29920 34886 29972 34892
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 29368 33652 29420 33658
rect 29368 33594 29420 33600
rect 29932 21321 29960 34886
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30300 29170 30328 30194
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30300 28218 30328 29106
rect 30288 28212 30340 28218
rect 30288 28154 30340 28160
rect 30104 24132 30156 24138
rect 30104 24074 30156 24080
rect 30116 23526 30144 24074
rect 30104 23520 30156 23526
rect 30104 23462 30156 23468
rect 29918 21312 29974 21321
rect 29918 21247 29974 21256
rect 29460 14884 29512 14890
rect 29460 14826 29512 14832
rect 29472 14414 29500 14826
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 30012 11212 30064 11218
rect 30012 11154 30064 11160
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29276 5364 29328 5370
rect 29276 5306 29328 5312
rect 29368 4140 29420 4146
rect 29368 4082 29420 4088
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29092 1692 29144 1698
rect 29092 1634 29144 1640
rect 29104 800 29132 1634
rect 29380 800 29408 4082
rect 29552 4004 29604 4010
rect 29552 3946 29604 3952
rect 29564 3777 29592 3946
rect 29550 3768 29606 3777
rect 29550 3703 29606 3712
rect 29656 2446 29684 6054
rect 29748 4185 29776 9862
rect 30024 9586 30052 11154
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 30012 7812 30064 7818
rect 30012 7754 30064 7760
rect 30024 6730 30052 7754
rect 30012 6724 30064 6730
rect 30012 6666 30064 6672
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 29828 4480 29880 4486
rect 29828 4422 29880 4428
rect 29734 4176 29790 4185
rect 29734 4111 29790 4120
rect 29840 4078 29868 4422
rect 29828 4072 29880 4078
rect 29828 4014 29880 4020
rect 29840 3670 29868 4014
rect 29828 3664 29880 3670
rect 29828 3606 29880 3612
rect 29932 3534 29960 6598
rect 30012 6180 30064 6186
rect 30012 6122 30064 6128
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29656 800 29684 2382
rect 29932 800 29960 3470
rect 30024 2378 30052 6122
rect 30116 2514 30144 23462
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30196 19780 30248 19786
rect 30196 19722 30248 19728
rect 30208 19514 30236 19722
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 30196 4480 30248 4486
rect 30196 4422 30248 4428
rect 30104 2508 30156 2514
rect 30104 2450 30156 2456
rect 30012 2372 30064 2378
rect 30012 2314 30064 2320
rect 30024 1698 30052 2314
rect 30012 1692 30064 1698
rect 30012 1634 30064 1640
rect 30208 800 30236 4422
rect 30300 3602 30328 21830
rect 30392 16182 30420 34886
rect 30484 21894 30512 36042
rect 30576 35766 30604 37198
rect 30564 35760 30616 35766
rect 30564 35702 30616 35708
rect 30564 35012 30616 35018
rect 30564 34954 30616 34960
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30576 16250 30604 34954
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30576 15162 30604 16050
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30564 11620 30616 11626
rect 30564 11562 30616 11568
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30392 8566 30420 11018
rect 30380 8560 30432 8566
rect 30380 8502 30432 8508
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30392 4622 30420 6598
rect 30472 6112 30524 6118
rect 30472 6054 30524 6060
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30392 4282 30420 4558
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30484 3058 30512 6054
rect 30576 4826 30604 11562
rect 30668 5914 30696 37266
rect 30944 36922 30972 39200
rect 31208 37188 31260 37194
rect 31208 37130 31260 37136
rect 30932 36916 30984 36922
rect 30932 36858 30984 36864
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 30932 36100 30984 36106
rect 30932 36042 30984 36048
rect 30840 30048 30892 30054
rect 30840 29990 30892 29996
rect 30748 28416 30800 28422
rect 30748 28358 30800 28364
rect 30760 28150 30788 28358
rect 30748 28144 30800 28150
rect 30748 28086 30800 28092
rect 30852 27962 30880 29990
rect 30760 27934 30880 27962
rect 30760 25974 30788 27934
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30852 27334 30880 27406
rect 30840 27328 30892 27334
rect 30840 27270 30892 27276
rect 30852 26586 30880 27270
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 30852 26042 30880 26522
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 30748 25968 30800 25974
rect 30748 25910 30800 25916
rect 30944 25498 30972 36042
rect 31036 34950 31064 36722
rect 31220 35834 31248 37130
rect 31312 36378 31340 39200
rect 31680 37244 31708 39200
rect 31760 37256 31812 37262
rect 31680 37216 31760 37244
rect 31760 37198 31812 37204
rect 31392 37120 31444 37126
rect 31392 37062 31444 37068
rect 31404 36854 31432 37062
rect 32048 36922 32076 39200
rect 32312 37324 32364 37330
rect 32312 37266 32364 37272
rect 32036 36916 32088 36922
rect 32036 36858 32088 36864
rect 31392 36848 31444 36854
rect 31392 36790 31444 36796
rect 31944 36780 31996 36786
rect 31944 36722 31996 36728
rect 31300 36372 31352 36378
rect 31300 36314 31352 36320
rect 31668 36168 31720 36174
rect 31668 36110 31720 36116
rect 31208 35828 31260 35834
rect 31208 35770 31260 35776
rect 31300 35692 31352 35698
rect 31300 35634 31352 35640
rect 31024 34944 31076 34950
rect 31024 34886 31076 34892
rect 31312 34202 31340 35634
rect 31680 35018 31708 36110
rect 31668 35012 31720 35018
rect 31668 34954 31720 34960
rect 31956 34950 31984 36722
rect 31944 34944 31996 34950
rect 31944 34886 31996 34892
rect 31300 34196 31352 34202
rect 31300 34138 31352 34144
rect 31576 29640 31628 29646
rect 31576 29582 31628 29588
rect 31588 29034 31616 29582
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31588 28218 31616 28970
rect 31576 28212 31628 28218
rect 31576 28154 31628 28160
rect 31588 27470 31616 28154
rect 31760 28076 31812 28082
rect 31760 28018 31812 28024
rect 31772 27674 31800 28018
rect 31760 27668 31812 27674
rect 31760 27610 31812 27616
rect 31772 27538 31800 27610
rect 31760 27532 31812 27538
rect 31760 27474 31812 27480
rect 31576 27464 31628 27470
rect 31576 27406 31628 27412
rect 30932 25492 30984 25498
rect 30932 25434 30984 25440
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31404 24206 31432 25298
rect 31576 25220 31628 25226
rect 31576 25162 31628 25168
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30668 5710 30696 5850
rect 30656 5704 30708 5710
rect 30656 5646 30708 5652
rect 30654 5264 30710 5273
rect 30654 5199 30656 5208
rect 30708 5199 30710 5208
rect 30656 5170 30708 5176
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30668 3942 30696 5170
rect 30746 4176 30802 4185
rect 30746 4111 30748 4120
rect 30800 4111 30802 4120
rect 30748 4082 30800 4088
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30484 800 30512 2994
rect 30760 800 30788 3470
rect 30852 3058 30880 24074
rect 31404 23798 31432 24142
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 31404 23186 31432 23734
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31404 22166 31432 23122
rect 31392 22160 31444 22166
rect 31392 22102 31444 22108
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30944 19378 30972 19654
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 31392 16584 31444 16590
rect 31392 16526 31444 16532
rect 31404 15706 31432 16526
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31392 14340 31444 14346
rect 31392 14282 31444 14288
rect 31404 14074 31432 14282
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31496 14006 31524 15302
rect 31484 14000 31536 14006
rect 31484 13942 31536 13948
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31404 11898 31432 12106
rect 31392 11892 31444 11898
rect 31392 11834 31444 11840
rect 31024 9444 31076 9450
rect 31024 9386 31076 9392
rect 30932 7268 30984 7274
rect 30932 7210 30984 7216
rect 30944 6934 30972 7210
rect 30932 6928 30984 6934
rect 30932 6870 30984 6876
rect 30932 6112 30984 6118
rect 30932 6054 30984 6060
rect 30944 4214 30972 6054
rect 31036 4622 31064 9386
rect 31206 6216 31262 6225
rect 31206 6151 31262 6160
rect 31220 5914 31248 6151
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31220 5234 31248 5850
rect 31300 5568 31352 5574
rect 31300 5510 31352 5516
rect 31312 5302 31340 5510
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 30932 4208 30984 4214
rect 30932 4150 30984 4156
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 31036 800 31064 3334
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 2106 31156 2246
rect 31116 2100 31168 2106
rect 31116 2042 31168 2048
rect 31312 800 31340 5238
rect 31484 4276 31536 4282
rect 31484 4218 31536 4224
rect 31496 3482 31524 4218
rect 31588 3670 31616 25162
rect 31956 16658 31984 34886
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 32140 32570 32168 33934
rect 32128 32564 32180 32570
rect 32128 32506 32180 32512
rect 32324 31754 32352 37266
rect 32416 35834 32444 39200
rect 32692 37244 32720 39200
rect 32772 37256 32824 37262
rect 32692 37216 32772 37244
rect 32772 37198 32824 37204
rect 33060 36938 33088 39200
rect 33060 36922 33180 36938
rect 33060 36916 33192 36922
rect 33060 36910 33140 36916
rect 33140 36858 33192 36864
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 32680 36100 32732 36106
rect 32680 36042 32732 36048
rect 32404 35828 32456 35834
rect 32404 35770 32456 35776
rect 32232 31726 32352 31754
rect 32036 30320 32088 30326
rect 32036 30262 32088 30268
rect 32048 29646 32076 30262
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 32036 29640 32088 29646
rect 32036 29582 32088 29588
rect 32140 29578 32168 30126
rect 32128 29572 32180 29578
rect 32128 29514 32180 29520
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 31944 16652 31996 16658
rect 31944 16594 31996 16600
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 31956 15570 31984 15982
rect 31944 15564 31996 15570
rect 31944 15506 31996 15512
rect 31852 13252 31904 13258
rect 31852 13194 31904 13200
rect 31864 7954 31892 13194
rect 32048 12434 32076 22374
rect 32140 12850 32168 22510
rect 32232 15706 32260 31726
rect 32588 30660 32640 30666
rect 32588 30602 32640 30608
rect 32600 30394 32628 30602
rect 32404 30388 32456 30394
rect 32404 30330 32456 30336
rect 32588 30388 32640 30394
rect 32588 30330 32640 30336
rect 32416 29714 32444 30330
rect 32404 29708 32456 29714
rect 32404 29650 32456 29656
rect 32588 29708 32640 29714
rect 32588 29650 32640 29656
rect 32600 28082 32628 29650
rect 32588 28076 32640 28082
rect 32588 28018 32640 28024
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32416 27470 32444 27814
rect 32600 27606 32628 28018
rect 32588 27600 32640 27606
rect 32588 27542 32640 27548
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32496 27328 32548 27334
rect 32496 27270 32548 27276
rect 32508 27062 32536 27270
rect 32496 27056 32548 27062
rect 32496 26998 32548 27004
rect 32600 26858 32628 27542
rect 32588 26852 32640 26858
rect 32588 26794 32640 26800
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 32324 16574 32352 23462
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32416 22574 32444 23054
rect 32692 22778 32720 36042
rect 33152 35894 33180 36722
rect 32968 35866 33180 35894
rect 32772 35692 32824 35698
rect 32772 35634 32824 35640
rect 32784 34950 32812 35634
rect 32772 34944 32824 34950
rect 32772 34886 32824 34892
rect 32680 22772 32732 22778
rect 32680 22714 32732 22720
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32692 22438 32720 22578
rect 32680 22432 32732 22438
rect 32680 22374 32732 22380
rect 32324 16546 32536 16574
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32404 12776 32456 12782
rect 32404 12718 32456 12724
rect 32048 12406 32168 12434
rect 31944 11552 31996 11558
rect 31944 11494 31996 11500
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 31852 6248 31904 6254
rect 31852 6190 31904 6196
rect 31760 6112 31812 6118
rect 31760 6054 31812 6060
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 31576 3664 31628 3670
rect 31576 3606 31628 3612
rect 31496 3454 31616 3482
rect 31680 3466 31708 4218
rect 31772 3534 31800 6054
rect 31864 4758 31892 6190
rect 31956 5370 31984 11494
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 32036 5092 32088 5098
rect 32036 5034 32088 5040
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 31392 2644 31444 2650
rect 31392 2586 31444 2592
rect 31404 2378 31432 2586
rect 31392 2372 31444 2378
rect 31392 2314 31444 2320
rect 31588 800 31616 3454
rect 31668 3460 31720 3466
rect 31668 3402 31720 3408
rect 31864 800 31892 3878
rect 31956 3466 31984 4966
rect 32048 3534 32076 5034
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 31944 3460 31996 3466
rect 31944 3402 31996 3408
rect 32140 2990 32168 12406
rect 32416 11830 32444 12718
rect 32404 11824 32456 11830
rect 32404 11766 32456 11772
rect 32220 9376 32272 9382
rect 32220 9318 32272 9324
rect 32232 4146 32260 9318
rect 32312 9036 32364 9042
rect 32312 8978 32364 8984
rect 32324 8566 32352 8978
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 32312 8424 32364 8430
rect 32312 8366 32364 8372
rect 32324 7818 32352 8366
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32312 7812 32364 7818
rect 32312 7754 32364 7760
rect 32324 6866 32352 7754
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 32312 6656 32364 6662
rect 32312 6598 32364 6604
rect 32324 4146 32352 6598
rect 32416 5370 32444 7822
rect 32404 5364 32456 5370
rect 32404 5306 32456 5312
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32220 4004 32272 4010
rect 32220 3946 32272 3952
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 32232 2514 32260 3946
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32220 2508 32272 2514
rect 32140 2468 32220 2496
rect 32140 800 32168 2468
rect 32220 2450 32272 2456
rect 32416 800 32444 2994
rect 32508 2514 32536 16546
rect 32784 8566 32812 34886
rect 32968 34542 32996 35866
rect 33428 35562 33456 39200
rect 33796 37262 33824 39200
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 33416 35556 33468 35562
rect 33416 35498 33468 35504
rect 33520 35290 33548 37198
rect 33692 37120 33744 37126
rect 33692 37062 33744 37068
rect 33508 35284 33560 35290
rect 33508 35226 33560 35232
rect 33232 34944 33284 34950
rect 33232 34886 33284 34892
rect 32956 34536 33008 34542
rect 32956 34478 33008 34484
rect 32864 32904 32916 32910
rect 32864 32846 32916 32852
rect 32876 32366 32904 32846
rect 32864 32360 32916 32366
rect 32864 32302 32916 32308
rect 32864 30864 32916 30870
rect 32864 30806 32916 30812
rect 32876 29850 32904 30806
rect 32864 29844 32916 29850
rect 32864 29786 32916 29792
rect 32772 8560 32824 8566
rect 32772 8502 32824 8508
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32600 3058 32628 6598
rect 32692 5914 32720 8434
rect 32968 8022 32996 34478
rect 33048 31340 33100 31346
rect 33048 31282 33100 31288
rect 33060 30938 33088 31282
rect 33140 31136 33192 31142
rect 33140 31078 33192 31084
rect 33048 30932 33100 30938
rect 33048 30874 33100 30880
rect 33152 30326 33180 31078
rect 33140 30320 33192 30326
rect 33140 30262 33192 30268
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 33060 20602 33088 21830
rect 33140 21344 33192 21350
rect 33140 21286 33192 21292
rect 33048 20596 33100 20602
rect 33048 20538 33100 20544
rect 32956 8016 33008 8022
rect 32956 7958 33008 7964
rect 32956 6112 33008 6118
rect 32956 6054 33008 6060
rect 32680 5908 32732 5914
rect 32680 5850 32732 5856
rect 32864 5296 32916 5302
rect 32864 5238 32916 5244
rect 32876 4321 32904 5238
rect 32968 5234 32996 6054
rect 32956 5228 33008 5234
rect 32956 5170 33008 5176
rect 32862 4312 32918 4321
rect 32862 4247 32918 4256
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 32692 800 32720 3334
rect 32968 800 32996 5170
rect 33152 4078 33180 21286
rect 33244 11354 33272 34886
rect 33600 33856 33652 33862
rect 33600 33798 33652 33804
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33428 19514 33456 19790
rect 33416 19508 33468 19514
rect 33416 19450 33468 19456
rect 33428 19378 33456 19450
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 33612 16574 33640 33798
rect 33520 16546 33640 16574
rect 33416 16108 33468 16114
rect 33416 16050 33468 16056
rect 33428 15910 33456 16050
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 33232 11348 33284 11354
rect 33232 11290 33284 11296
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 33244 800 33272 5510
rect 33428 2281 33456 15846
rect 33520 4978 33548 16546
rect 33704 13326 33732 37062
rect 34164 36922 34192 39200
rect 34152 36916 34204 36922
rect 34152 36858 34204 36864
rect 34336 36848 34388 36854
rect 34336 36790 34388 36796
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 34152 36100 34204 36106
rect 34152 36042 34204 36048
rect 33968 35692 34020 35698
rect 33968 35634 34020 35640
rect 34060 35692 34112 35698
rect 34060 35634 34112 35640
rect 33980 34542 34008 35634
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 33980 17202 34008 34478
rect 34072 33862 34100 35634
rect 34060 33856 34112 33862
rect 34060 33798 34112 33804
rect 34164 22094 34192 36042
rect 34256 34950 34284 36722
rect 34244 34944 34296 34950
rect 34244 34886 34296 34892
rect 34244 32428 34296 32434
rect 34244 32370 34296 32376
rect 34256 31210 34284 32370
rect 34244 31204 34296 31210
rect 34244 31146 34296 31152
rect 34072 22066 34192 22094
rect 33968 17196 34020 17202
rect 33968 17138 34020 17144
rect 33692 13320 33744 13326
rect 33692 13262 33744 13268
rect 33692 12640 33744 12646
rect 33692 12582 33744 12588
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33612 5370 33640 8434
rect 33600 5364 33652 5370
rect 33600 5306 33652 5312
rect 33520 4950 33640 4978
rect 33506 4856 33562 4865
rect 33506 4791 33508 4800
rect 33560 4791 33562 4800
rect 33508 4762 33560 4768
rect 33612 4758 33640 4950
rect 33600 4752 33652 4758
rect 33600 4694 33652 4700
rect 33508 4548 33560 4554
rect 33508 4490 33560 4496
rect 33520 3641 33548 4490
rect 33506 3632 33562 3641
rect 33506 3567 33562 3576
rect 33704 3534 33732 12582
rect 34072 9178 34100 22066
rect 34348 17338 34376 36790
rect 34440 36394 34468 39200
rect 34612 37120 34664 37126
rect 34612 37062 34664 37068
rect 34440 36378 34560 36394
rect 34440 36372 34572 36378
rect 34440 36366 34520 36372
rect 34520 36314 34572 36320
rect 34624 35894 34652 37062
rect 34808 36922 34836 39200
rect 35176 37754 35204 39200
rect 35176 37726 35388 37754
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34888 37120 34940 37126
rect 34888 37062 34940 37068
rect 34796 36916 34848 36922
rect 34796 36858 34848 36864
rect 34900 36854 34928 37062
rect 35360 36922 35388 37726
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 35348 36916 35400 36922
rect 35348 36858 35400 36864
rect 34888 36848 34940 36854
rect 34888 36790 34940 36796
rect 34796 36780 34848 36786
rect 34796 36722 34848 36728
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 34532 35866 34652 35894
rect 34428 30932 34480 30938
rect 34428 30874 34480 30880
rect 34440 28150 34468 30874
rect 34428 28144 34480 28150
rect 34428 28086 34480 28092
rect 34440 27606 34468 28086
rect 34428 27600 34480 27606
rect 34428 27542 34480 27548
rect 34440 27130 34468 27542
rect 34428 27124 34480 27130
rect 34428 27066 34480 27072
rect 34428 18692 34480 18698
rect 34428 18634 34480 18640
rect 34336 17332 34388 17338
rect 34336 17274 34388 17280
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34164 16250 34192 17070
rect 34440 16250 34468 18634
rect 34532 16574 34560 35866
rect 34716 35170 34744 36110
rect 34624 35142 34744 35170
rect 34624 33862 34652 35142
rect 34808 35034 34836 36722
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35452 36378 35480 37198
rect 35440 36372 35492 36378
rect 35440 36314 35492 36320
rect 35544 35834 35572 39200
rect 35622 39128 35678 39137
rect 35622 39063 35678 39072
rect 35532 35828 35584 35834
rect 35532 35770 35584 35776
rect 35440 35692 35492 35698
rect 35440 35634 35492 35640
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34716 35006 34836 35034
rect 34716 34950 34744 35006
rect 34704 34944 34756 34950
rect 34704 34886 34756 34892
rect 34612 33856 34664 33862
rect 34610 33824 34612 33833
rect 34664 33824 34666 33833
rect 34610 33759 34666 33768
rect 34716 21350 34744 34886
rect 35254 34640 35310 34649
rect 35254 34575 35256 34584
rect 35308 34575 35310 34584
rect 35256 34546 35308 34552
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35452 33862 35480 35634
rect 35532 35624 35584 35630
rect 35532 35566 35584 35572
rect 35440 33856 35492 33862
rect 35440 33798 35492 33804
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 27872 34848 27878
rect 34796 27814 34848 27820
rect 34808 25294 34836 27814
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34796 22636 34848 22642
rect 34796 22578 34848 22584
rect 34808 21962 34836 22578
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34796 21956 34848 21962
rect 34796 21898 34848 21904
rect 34704 21344 34756 21350
rect 34704 21286 34756 21292
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34704 19440 34756 19446
rect 34704 19382 34756 19388
rect 34716 18970 34744 19382
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34532 16546 34652 16574
rect 34152 16244 34204 16250
rect 34152 16186 34204 16192
rect 34428 16244 34480 16250
rect 34428 16186 34480 16192
rect 34060 9172 34112 9178
rect 34060 9114 34112 9120
rect 34624 8634 34652 16546
rect 34808 15706 34836 19314
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34716 14618 34744 15438
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34704 14612 34756 14618
rect 34704 14554 34756 14560
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 33876 6656 33928 6662
rect 33876 6598 33928 6604
rect 33888 5234 33916 6598
rect 33980 5914 34008 7346
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 34520 6724 34572 6730
rect 34520 6666 34572 6672
rect 34532 6338 34560 6666
rect 34440 6310 34560 6338
rect 34060 6112 34112 6118
rect 34060 6054 34112 6060
rect 33968 5908 34020 5914
rect 33968 5850 34020 5856
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33692 3528 33744 3534
rect 33692 3470 33744 3476
rect 33796 3058 33824 3878
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33414 2272 33470 2281
rect 33414 2207 33470 2216
rect 33520 800 33548 2790
rect 33888 2774 33916 5170
rect 33980 4622 34008 5850
rect 34072 5710 34100 6054
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 33968 4140 34020 4146
rect 33968 4082 34020 4088
rect 33980 3369 34008 4082
rect 33966 3360 34022 3369
rect 33966 3295 34022 3304
rect 33796 2746 33916 2774
rect 33796 800 33824 2746
rect 34072 800 34100 5646
rect 34244 5228 34296 5234
rect 34244 5170 34296 5176
rect 34152 4480 34204 4486
rect 34152 4422 34204 4428
rect 34164 4146 34192 4422
rect 34256 4282 34284 5170
rect 34244 4276 34296 4282
rect 34244 4218 34296 4224
rect 34152 4140 34204 4146
rect 34152 4082 34204 4088
rect 34440 3942 34468 6310
rect 34520 6180 34572 6186
rect 34520 6122 34572 6128
rect 34428 3936 34480 3942
rect 34150 3904 34206 3913
rect 34428 3878 34480 3884
rect 34150 3839 34206 3848
rect 34164 3670 34192 3839
rect 34152 3664 34204 3670
rect 34532 3618 34560 6122
rect 34152 3606 34204 3612
rect 34256 3590 34560 3618
rect 34256 2446 34284 3590
rect 34520 3460 34572 3466
rect 34520 3402 34572 3408
rect 34336 3392 34388 3398
rect 34336 3334 34388 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34244 2440 34296 2446
rect 34244 2382 34296 2388
rect 34348 800 34376 3334
rect 34440 3126 34468 3334
rect 34428 3120 34480 3126
rect 34428 3062 34480 3068
rect 34532 1902 34560 3402
rect 34624 2446 34652 7142
rect 34716 2650 34744 14554
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34796 8900 34848 8906
rect 34796 8842 34848 8848
rect 34808 5914 34836 8842
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35348 7744 35400 7750
rect 35348 7686 35400 7692
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35360 6984 35388 7686
rect 35268 6956 35388 6984
rect 35268 6322 35296 6956
rect 35348 6724 35400 6730
rect 35348 6666 35400 6672
rect 35256 6316 35308 6322
rect 35256 6258 35308 6264
rect 35268 6225 35296 6258
rect 35254 6216 35310 6225
rect 35254 6151 35310 6160
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34796 5908 34848 5914
rect 34796 5850 34848 5856
rect 34886 5536 34942 5545
rect 34886 5471 34942 5480
rect 34900 5370 34928 5471
rect 34888 5364 34940 5370
rect 34888 5306 34940 5312
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35360 4026 35388 6666
rect 35452 4758 35480 33798
rect 35544 33318 35572 35566
rect 35636 35290 35664 39063
rect 35806 37496 35862 37505
rect 35806 37431 35862 37440
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35728 36854 35756 37198
rect 35716 36848 35768 36854
rect 35716 36790 35768 36796
rect 35624 35284 35676 35290
rect 35624 35226 35676 35232
rect 35820 34746 35848 37431
rect 35912 37262 35940 39200
rect 35900 37256 35952 37262
rect 36280 37244 36308 39200
rect 36280 37216 36400 37244
rect 35900 37198 35952 37204
rect 36268 37120 36320 37126
rect 36268 37062 36320 37068
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 35992 35080 36044 35086
rect 35992 35022 36044 35028
rect 36084 35080 36136 35086
rect 36084 35022 36136 35028
rect 35808 34740 35860 34746
rect 35808 34682 35860 34688
rect 35808 34400 35860 34406
rect 35808 34342 35860 34348
rect 35820 34241 35848 34342
rect 35806 34232 35862 34241
rect 36004 34202 36032 35022
rect 36096 34202 36124 35022
rect 36188 34610 36216 36722
rect 36280 36553 36308 37062
rect 36372 36922 36400 37216
rect 36360 36916 36412 36922
rect 36360 36858 36412 36864
rect 36266 36544 36322 36553
rect 36266 36479 36322 36488
rect 36360 35692 36412 35698
rect 36360 35634 36412 35640
rect 36176 34604 36228 34610
rect 36176 34546 36228 34552
rect 35806 34167 35862 34176
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 36084 34196 36136 34202
rect 36084 34138 36136 34144
rect 35532 33312 35584 33318
rect 35532 33254 35584 33260
rect 35544 5370 35572 33254
rect 36004 31414 36032 34138
rect 36372 33318 36400 35634
rect 36556 35562 36584 39200
rect 36924 39114 36952 39200
rect 37016 39114 37044 39222
rect 36924 39086 37044 39114
rect 37200 37244 37228 39222
rect 37278 39200 37334 40000
rect 37646 39200 37702 40000
rect 38014 39200 38070 40000
rect 38290 39200 38346 40000
rect 38658 39200 38714 40000
rect 39026 39200 39082 40000
rect 39394 39200 39450 40000
rect 39762 39200 39818 40000
rect 37292 37618 37320 39200
rect 37292 37590 37412 37618
rect 37280 37256 37332 37262
rect 37200 37216 37280 37244
rect 37280 37198 37332 37204
rect 36726 35864 36782 35873
rect 37292 35834 37320 37198
rect 36726 35799 36782 35808
rect 37280 35828 37332 35834
rect 36544 35556 36596 35562
rect 36544 35498 36596 35504
rect 36452 35012 36504 35018
rect 36452 34954 36504 34960
rect 36360 33312 36412 33318
rect 36360 33254 36412 33260
rect 35992 31408 36044 31414
rect 35992 31350 36044 31356
rect 36004 30938 36032 31350
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 35716 27532 35768 27538
rect 35716 27474 35768 27480
rect 35728 26994 35756 27474
rect 36268 27396 36320 27402
rect 36268 27338 36320 27344
rect 36280 27062 36308 27338
rect 36268 27056 36320 27062
rect 36268 26998 36320 27004
rect 35716 26988 35768 26994
rect 35716 26930 35768 26936
rect 35900 23656 35952 23662
rect 35900 23598 35952 23604
rect 35912 22710 35940 23598
rect 35900 22704 35952 22710
rect 35900 22646 35952 22652
rect 35912 22094 35940 22646
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 35912 22066 36032 22094
rect 36004 19514 36032 22066
rect 36096 21010 36124 22374
rect 36084 21004 36136 21010
rect 36084 20946 36136 20952
rect 35992 19508 36044 19514
rect 35992 19450 36044 19456
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 36004 14822 36032 14962
rect 35992 14816 36044 14822
rect 35992 14758 36044 14764
rect 35900 10600 35952 10606
rect 35900 10542 35952 10548
rect 35808 10124 35860 10130
rect 35808 10066 35860 10072
rect 35820 8974 35848 10066
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35716 7812 35768 7818
rect 35716 7754 35768 7760
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35636 5710 35664 6734
rect 35624 5704 35676 5710
rect 35624 5646 35676 5652
rect 35532 5364 35584 5370
rect 35532 5306 35584 5312
rect 35440 4752 35492 4758
rect 35440 4694 35492 4700
rect 35360 3998 35480 4026
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34808 3652 34836 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34808 3624 34928 3652
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 34808 2530 34836 3470
rect 34900 3126 34928 3624
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35176 3194 35204 3402
rect 35164 3188 35216 3194
rect 35164 3130 35216 3136
rect 34888 3120 34940 3126
rect 34888 3062 34940 3068
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34808 2502 34928 2530
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34520 1896 34572 1902
rect 34520 1838 34572 1844
rect 34624 800 34652 2382
rect 34900 800 34928 2502
rect 35360 1986 35388 3878
rect 35452 3534 35480 3998
rect 35440 3528 35492 3534
rect 35440 3470 35492 3476
rect 35728 3126 35756 7754
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35820 5642 35848 6598
rect 35912 6458 35940 10542
rect 36004 7410 36032 14758
rect 36084 9036 36136 9042
rect 36084 8978 36136 8984
rect 36096 8566 36124 8978
rect 36084 8560 36136 8566
rect 36084 8502 36136 8508
rect 35992 7404 36044 7410
rect 35992 7346 36044 7352
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 36004 6390 36032 7142
rect 35992 6384 36044 6390
rect 35992 6326 36044 6332
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35808 5636 35860 5642
rect 35808 5578 35860 5584
rect 35912 5522 35940 6258
rect 36096 5778 36124 8502
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36176 7200 36228 7206
rect 36176 7142 36228 7148
rect 36084 5772 36136 5778
rect 36084 5714 36136 5720
rect 35820 5494 35940 5522
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 35820 4185 35848 5494
rect 36096 4622 36124 5510
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 35992 4480 36044 4486
rect 35992 4422 36044 4428
rect 35806 4176 35862 4185
rect 35806 4111 35862 4120
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 35716 3120 35768 3126
rect 35716 3062 35768 3068
rect 35176 1958 35388 1986
rect 35176 800 35204 1958
rect 35452 800 35480 3062
rect 35716 2372 35768 2378
rect 35716 2314 35768 2320
rect 35728 800 35756 2314
rect 36004 800 36032 4422
rect 36188 2530 36216 7142
rect 36280 4214 36308 8298
rect 36268 4208 36320 4214
rect 36268 4150 36320 4156
rect 36096 2514 36216 2530
rect 36084 2508 36216 2514
rect 36136 2502 36216 2508
rect 36084 2450 36136 2456
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 36188 1766 36216 2382
rect 36176 1760 36228 1766
rect 36176 1702 36228 1708
rect 36280 800 36308 4150
rect 36372 3194 36400 33254
rect 36464 31346 36492 34954
rect 36740 34066 36768 35799
rect 37280 35770 37332 35776
rect 37384 35562 37412 37590
rect 37556 36644 37608 36650
rect 37556 36586 37608 36592
rect 37568 36242 37596 36586
rect 37464 36236 37516 36242
rect 37464 36178 37516 36184
rect 37556 36236 37608 36242
rect 37556 36178 37608 36184
rect 37372 35556 37424 35562
rect 37372 35498 37424 35504
rect 37280 35080 37332 35086
rect 37280 35022 37332 35028
rect 37292 34746 37320 35022
rect 37280 34740 37332 34746
rect 37280 34682 37332 34688
rect 37188 34672 37240 34678
rect 37188 34614 37240 34620
rect 36912 34536 36964 34542
rect 36912 34478 36964 34484
rect 36728 34060 36780 34066
rect 36728 34002 36780 34008
rect 36636 33992 36688 33998
rect 36556 33940 36636 33946
rect 36556 33934 36688 33940
rect 36556 33918 36676 33934
rect 36556 32774 36584 33918
rect 36740 33658 36768 34002
rect 36728 33652 36780 33658
rect 36728 33594 36780 33600
rect 36924 32774 36952 34478
rect 37200 34202 37228 34614
rect 37188 34196 37240 34202
rect 37188 34138 37240 34144
rect 36544 32768 36596 32774
rect 36544 32710 36596 32716
rect 36912 32768 36964 32774
rect 36912 32710 36964 32716
rect 36452 31340 36504 31346
rect 36452 31282 36504 31288
rect 36450 15464 36506 15473
rect 36450 15399 36452 15408
rect 36504 15399 36506 15408
rect 36452 15370 36504 15376
rect 36556 15162 36584 32710
rect 36636 15360 36688 15366
rect 36636 15302 36688 15308
rect 36544 15156 36596 15162
rect 36544 15098 36596 15104
rect 36452 8832 36504 8838
rect 36452 8774 36504 8780
rect 36464 5234 36492 8774
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 36452 5228 36504 5234
rect 36452 5170 36504 5176
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36464 3738 36492 3878
rect 36452 3732 36504 3738
rect 36452 3674 36504 3680
rect 36556 3505 36584 7346
rect 36648 5710 36676 15302
rect 36728 14476 36780 14482
rect 36728 14418 36780 14424
rect 36740 13530 36768 14418
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36924 8090 36952 32710
rect 37188 30728 37240 30734
rect 37188 30670 37240 30676
rect 37200 29850 37228 30670
rect 37188 29844 37240 29850
rect 37188 29786 37240 29792
rect 37476 23866 37504 36178
rect 37556 34604 37608 34610
rect 37556 34546 37608 34552
rect 37568 27606 37596 34546
rect 37660 34202 37688 39200
rect 38028 36854 38056 39200
rect 38016 36848 38068 36854
rect 38016 36790 38068 36796
rect 37832 35692 37884 35698
rect 37832 35634 37884 35640
rect 37648 34196 37700 34202
rect 37648 34138 37700 34144
rect 37740 33992 37792 33998
rect 37740 33934 37792 33940
rect 37752 32230 37780 33934
rect 37844 33658 37872 35634
rect 37924 34740 37976 34746
rect 38028 34728 38056 36790
rect 38304 35290 38332 39200
rect 38384 37188 38436 37194
rect 38384 37130 38436 37136
rect 38292 35284 38344 35290
rect 38292 35226 38344 35232
rect 38292 35080 38344 35086
rect 38292 35022 38344 35028
rect 37976 34700 38056 34728
rect 37924 34682 37976 34688
rect 37832 33652 37884 33658
rect 37832 33594 37884 33600
rect 37832 33516 37884 33522
rect 37832 33458 37884 33464
rect 37740 32224 37792 32230
rect 37740 32166 37792 32172
rect 37556 27600 37608 27606
rect 37556 27542 37608 27548
rect 37568 23866 37596 27542
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37556 23860 37608 23866
rect 37556 23802 37608 23808
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 37660 22982 37688 23666
rect 37556 22976 37608 22982
rect 37556 22918 37608 22924
rect 37648 22976 37700 22982
rect 37648 22918 37700 22924
rect 37568 22710 37596 22918
rect 37556 22704 37608 22710
rect 37556 22646 37608 22652
rect 37096 20936 37148 20942
rect 37096 20878 37148 20884
rect 36912 8084 36964 8090
rect 36912 8026 36964 8032
rect 36728 7812 36780 7818
rect 36728 7754 36780 7760
rect 36636 5704 36688 5710
rect 36636 5646 36688 5652
rect 36542 3496 36598 3505
rect 36542 3431 36598 3440
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36464 2582 36492 2994
rect 36452 2576 36504 2582
rect 36452 2518 36504 2524
rect 36544 2508 36596 2514
rect 36544 2450 36596 2456
rect 36556 800 36584 2450
rect 36740 2310 36768 7754
rect 37108 5710 37136 20878
rect 37556 19372 37608 19378
rect 37556 19314 37608 19320
rect 37372 15020 37424 15026
rect 37372 14962 37424 14968
rect 37280 14408 37332 14414
rect 37280 14350 37332 14356
rect 37292 14249 37320 14350
rect 37278 14240 37334 14249
rect 37278 14175 37334 14184
rect 37280 10464 37332 10470
rect 37280 10406 37332 10412
rect 37292 6798 37320 10406
rect 37280 6792 37332 6798
rect 37280 6734 37332 6740
rect 37384 6662 37412 14962
rect 37464 8356 37516 8362
rect 37464 8298 37516 8304
rect 37372 6656 37424 6662
rect 37372 6598 37424 6604
rect 37372 6384 37424 6390
rect 37372 6326 37424 6332
rect 37096 5704 37148 5710
rect 37096 5646 37148 5652
rect 37278 5400 37334 5409
rect 37384 5370 37412 6326
rect 37278 5335 37334 5344
rect 37372 5364 37424 5370
rect 37292 5250 37320 5335
rect 37372 5306 37424 5312
rect 37292 5222 37412 5250
rect 36820 5024 36872 5030
rect 36820 4966 36872 4972
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36832 800 36860 4966
rect 37096 4616 37148 4622
rect 37096 4558 37148 4564
rect 37186 4584 37242 4593
rect 37108 2553 37136 4558
rect 37186 4519 37188 4528
rect 37240 4519 37242 4528
rect 37280 4548 37332 4554
rect 37188 4490 37240 4496
rect 37280 4490 37332 4496
rect 37292 4264 37320 4490
rect 37200 4236 37320 4264
rect 37094 2544 37150 2553
rect 37094 2479 37150 2488
rect 37200 2394 37228 4236
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 37292 3602 37320 4082
rect 37280 3596 37332 3602
rect 37280 3538 37332 3544
rect 37384 2990 37412 5222
rect 37476 3058 37504 8298
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 37476 2774 37504 2994
rect 37108 2366 37228 2394
rect 37384 2746 37504 2774
rect 37108 800 37136 2366
rect 37384 800 37412 2746
rect 37568 2514 37596 19314
rect 37660 3602 37688 22918
rect 37740 16448 37792 16454
rect 37740 16390 37792 16396
rect 37752 16114 37780 16390
rect 37844 16250 37872 33458
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38120 32502 38148 32846
rect 38108 32496 38160 32502
rect 38106 32464 38108 32473
rect 38160 32464 38162 32473
rect 38106 32399 38162 32408
rect 38108 31340 38160 31346
rect 38108 31282 38160 31288
rect 38120 30841 38148 31282
rect 38106 30832 38162 30841
rect 38106 30767 38162 30776
rect 38108 29640 38160 29646
rect 38108 29582 38160 29588
rect 38120 29209 38148 29582
rect 38106 29200 38162 29209
rect 38106 29135 38162 29144
rect 38108 28076 38160 28082
rect 38108 28018 38160 28024
rect 38120 27577 38148 28018
rect 38106 27568 38162 27577
rect 38106 27503 38162 27512
rect 38106 25800 38162 25809
rect 38106 25735 38108 25744
rect 38160 25735 38162 25744
rect 38108 25706 38160 25712
rect 38014 24168 38070 24177
rect 38014 24103 38016 24112
rect 38068 24103 38070 24112
rect 38016 24074 38068 24080
rect 37924 24064 37976 24070
rect 37924 24006 37976 24012
rect 37936 22574 37964 24006
rect 38200 22704 38252 22710
rect 38200 22646 38252 22652
rect 37924 22568 37976 22574
rect 37924 22510 37976 22516
rect 38106 22536 38162 22545
rect 38106 22471 38162 22480
rect 38120 22030 38148 22471
rect 38108 22024 38160 22030
rect 38108 21966 38160 21972
rect 38106 20904 38162 20913
rect 38106 20839 38162 20848
rect 38120 20466 38148 20839
rect 38108 20460 38160 20466
rect 38108 20402 38160 20408
rect 38106 19136 38162 19145
rect 38106 19071 38162 19080
rect 38120 18766 38148 19071
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 38120 17513 38148 17614
rect 38106 17504 38162 17513
rect 38106 17439 38162 17448
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37740 16108 37792 16114
rect 37740 16050 37792 16056
rect 37924 16040 37976 16046
rect 37924 15982 37976 15988
rect 37936 15706 37964 15982
rect 38014 15872 38070 15881
rect 38014 15807 38070 15816
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 38028 15502 38056 15807
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 38028 15162 38056 15438
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37752 13190 37780 13874
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 38108 12640 38160 12646
rect 38108 12582 38160 12588
rect 38120 12481 38148 12582
rect 38106 12472 38162 12481
rect 38106 12407 38162 12416
rect 38212 12434 38240 22646
rect 38304 14006 38332 35022
rect 38292 14000 38344 14006
rect 38292 13942 38344 13948
rect 38212 12406 38332 12434
rect 37924 12096 37976 12102
rect 37924 12038 37976 12044
rect 37936 11354 37964 12038
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 38108 11144 38160 11150
rect 38108 11086 38160 11092
rect 38120 10849 38148 11086
rect 38106 10840 38162 10849
rect 38106 10775 38162 10784
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 37752 6458 37780 9522
rect 38106 9208 38162 9217
rect 38106 9143 38162 9152
rect 38120 8974 38148 9143
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 37832 8628 37884 8634
rect 37832 8570 37884 8576
rect 37844 7478 37872 8570
rect 37924 8424 37976 8430
rect 37924 8366 37976 8372
rect 37832 7472 37884 7478
rect 37832 7414 37884 7420
rect 37832 7336 37884 7342
rect 37832 7278 37884 7284
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37740 6112 37792 6118
rect 37740 6054 37792 6060
rect 37752 5846 37780 6054
rect 37740 5840 37792 5846
rect 37740 5782 37792 5788
rect 37740 5568 37792 5574
rect 37740 5510 37792 5516
rect 37648 3596 37700 3602
rect 37648 3538 37700 3544
rect 37752 2774 37780 5510
rect 37660 2746 37780 2774
rect 37556 2508 37608 2514
rect 37556 2450 37608 2456
rect 37660 800 37688 2746
rect 37844 2446 37872 7278
rect 37936 4554 37964 8366
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 38120 7585 38148 7822
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38106 7576 38162 7585
rect 38106 7511 38162 7520
rect 38108 7200 38160 7206
rect 38108 7142 38160 7148
rect 38014 5808 38070 5817
rect 38014 5743 38070 5752
rect 38028 5642 38056 5743
rect 38016 5636 38068 5642
rect 38016 5578 38068 5584
rect 38120 5234 38148 7142
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 37832 2440 37884 2446
rect 37884 2388 37964 2394
rect 37832 2382 37964 2388
rect 37844 2366 37964 2382
rect 37936 800 37964 2366
rect 38120 921 38148 5170
rect 38212 3602 38240 7686
rect 38200 3596 38252 3602
rect 38200 3538 38252 3544
rect 38106 912 38162 921
rect 38106 847 38162 856
rect 38212 800 38240 3538
rect 38304 3126 38332 12406
rect 38396 4146 38424 37130
rect 38568 36644 38620 36650
rect 38568 36586 38620 36592
rect 38476 36168 38528 36174
rect 38476 36110 38528 36116
rect 38488 19310 38516 36110
rect 38476 19304 38528 19310
rect 38476 19246 38528 19252
rect 38476 13184 38528 13190
rect 38476 13126 38528 13132
rect 38488 6746 38516 13126
rect 38580 8634 38608 36586
rect 38672 33658 38700 39200
rect 39040 35698 39068 39200
rect 39028 35692 39080 35698
rect 39028 35634 39080 35640
rect 38752 35488 38804 35494
rect 38752 35430 38804 35436
rect 38660 33652 38712 33658
rect 38660 33594 38712 33600
rect 38660 32224 38712 32230
rect 38660 32166 38712 32172
rect 38568 8628 38620 8634
rect 38568 8570 38620 8576
rect 38488 6718 38608 6746
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 38396 3534 38424 4082
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 38292 3120 38344 3126
rect 38292 3062 38344 3068
rect 38488 800 38516 6598
rect 38580 3398 38608 6718
rect 38672 4010 38700 32166
rect 38764 6390 38792 35430
rect 39408 34746 39436 39200
rect 39396 34740 39448 34746
rect 39396 34682 39448 34688
rect 39776 34678 39804 39200
rect 39764 34672 39816 34678
rect 39764 34614 39816 34620
rect 38936 16108 38988 16114
rect 38936 16050 38988 16056
rect 38752 6384 38804 6390
rect 38752 6326 38804 6332
rect 38660 4004 38712 4010
rect 38660 3946 38712 3952
rect 38948 3466 38976 16050
rect 39580 6724 39632 6730
rect 39580 6666 39632 6672
rect 39028 6316 39080 6322
rect 39028 6258 39080 6264
rect 38936 3460 38988 3466
rect 38936 3402 38988 3408
rect 38568 3392 38620 3398
rect 38568 3334 38620 3340
rect 38752 2916 38804 2922
rect 38752 2858 38804 2864
rect 38764 800 38792 2858
rect 39040 800 39068 6258
rect 39304 5908 39356 5914
rect 39304 5850 39356 5856
rect 39316 800 39344 5850
rect 39592 800 39620 6666
rect 39854 6216 39910 6225
rect 39854 6151 39910 6160
rect 39868 800 39896 6151
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
<< via2 >>
rect 1582 29960 1638 30016
rect 1950 8336 2006 8392
rect 3422 9968 3478 10024
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4710 5636 4766 5672
rect 4710 5616 4712 5636
rect 4712 5616 4764 5636
rect 4764 5616 4766 5636
rect 3422 2352 3478 2408
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3882 4428 3884 4448
rect 3884 4428 3936 4448
rect 3936 4428 3938 4448
rect 3882 4392 3938 4428
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4158 3304 4214 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4894 3168 4950 3224
rect 5538 2896 5594 2952
rect 6090 3712 6146 3768
rect 7470 36216 7526 36272
rect 9218 36116 9220 36136
rect 9220 36116 9272 36136
rect 9272 36116 9274 36136
rect 9218 36080 9274 36116
rect 12254 36352 12310 36408
rect 8482 3848 8538 3904
rect 8298 3612 8300 3632
rect 8300 3612 8352 3632
rect 8352 3612 8354 3632
rect 8298 3576 8354 3612
rect 8206 3304 8262 3360
rect 8390 1536 8446 1592
rect 9218 4120 9274 4176
rect 9954 7792 10010 7848
rect 10598 4004 10654 4040
rect 10598 3984 10600 4004
rect 10600 3984 10652 4004
rect 10652 3984 10654 4004
rect 10506 2760 10562 2816
rect 10966 3440 11022 3496
rect 11058 3340 11060 3360
rect 11060 3340 11112 3360
rect 11112 3340 11114 3360
rect 11058 3304 11114 3340
rect 10782 2624 10838 2680
rect 11518 3984 11574 4040
rect 11334 3440 11390 3496
rect 12070 6160 12126 6216
rect 12070 3984 12126 4040
rect 12070 3576 12126 3632
rect 12438 2796 12440 2816
rect 12440 2796 12492 2816
rect 12492 2796 12494 2816
rect 12438 2760 12494 2796
rect 14278 1672 14334 1728
rect 14554 3032 14610 3088
rect 15382 3188 15438 3224
rect 15382 3168 15384 3188
rect 15384 3168 15436 3188
rect 15436 3168 15438 3188
rect 15014 1808 15070 1864
rect 16854 3576 16910 3632
rect 17498 3304 17554 3360
rect 18510 4528 18566 4584
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 20166 36896 20222 36952
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19062 4020 19064 4040
rect 19064 4020 19116 4040
rect 19116 4020 19118 4040
rect 19062 3984 19118 4020
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 3848 19946 3904
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22374 34348 22376 34368
rect 22376 34348 22428 34368
rect 22428 34348 22430 34368
rect 22374 34312 22430 34348
rect 22282 13252 22338 13288
rect 22282 13232 22284 13252
rect 22284 13232 22336 13252
rect 22336 13232 22338 13252
rect 20626 3984 20682 4040
rect 20810 4392 20866 4448
rect 20626 2216 20682 2272
rect 20442 1536 20498 1592
rect 22098 4120 22154 4176
rect 23202 13252 23258 13288
rect 23202 13232 23204 13252
rect 23204 13232 23256 13252
rect 23256 13232 23258 13252
rect 23662 14884 23718 14920
rect 23662 14864 23664 14884
rect 23664 14864 23716 14884
rect 23716 14864 23718 14884
rect 23478 8356 23534 8392
rect 23478 8336 23480 8356
rect 23480 8336 23532 8356
rect 23532 8336 23534 8356
rect 24306 13948 24308 13968
rect 24308 13948 24360 13968
rect 24360 13948 24362 13968
rect 24306 13912 24362 13948
rect 22650 5344 22706 5400
rect 23018 3848 23074 3904
rect 23386 3576 23442 3632
rect 23294 3440 23350 3496
rect 23938 4256 23994 4312
rect 24766 3460 24822 3496
rect 24766 3440 24768 3460
rect 24768 3440 24820 3460
rect 24820 3440 24822 3460
rect 24858 1944 24914 2000
rect 25226 1672 25282 1728
rect 25594 3340 25596 3360
rect 25596 3340 25648 3360
rect 25648 3340 25650 3360
rect 25594 3304 25650 3340
rect 25502 1808 25558 1864
rect 28998 36080 29054 36136
rect 27342 3032 27398 3088
rect 27342 2372 27398 2408
rect 27342 2352 27344 2372
rect 27344 2352 27396 2372
rect 27396 2352 27398 2372
rect 27526 2916 27582 2952
rect 27526 2896 27528 2916
rect 27528 2896 27580 2916
rect 27580 2896 27582 2916
rect 28078 2488 28134 2544
rect 28814 7792 28870 7848
rect 28722 4392 28778 4448
rect 30102 36352 30158 36408
rect 30194 36216 30250 36272
rect 29918 21256 29974 21312
rect 29550 3712 29606 3768
rect 29734 4120 29790 4176
rect 30654 5228 30710 5264
rect 30654 5208 30656 5228
rect 30656 5208 30708 5228
rect 30708 5208 30710 5228
rect 30746 4140 30802 4176
rect 30746 4120 30748 4140
rect 30748 4120 30800 4140
rect 30800 4120 30802 4140
rect 31206 6160 31262 6216
rect 32862 4256 32918 4312
rect 33506 4820 33562 4856
rect 33506 4800 33508 4820
rect 33508 4800 33560 4820
rect 33560 4800 33562 4820
rect 33506 3576 33562 3632
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35622 39072 35678 39128
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34610 33804 34612 33824
rect 34612 33804 34664 33824
rect 34664 33804 34666 33824
rect 34610 33768 34666 33804
rect 35254 34604 35310 34640
rect 35254 34584 35256 34604
rect 35256 34584 35308 34604
rect 35308 34584 35310 34604
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 33414 2216 33470 2272
rect 33966 3304 34022 3360
rect 34150 3848 34206 3904
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35254 6160 35310 6216
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34886 5480 34942 5536
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35806 37440 35862 37496
rect 35806 34176 35862 34232
rect 36266 36488 36322 36544
rect 36726 35808 36782 35864
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35806 4120 35862 4176
rect 36450 15428 36506 15464
rect 36450 15408 36452 15428
rect 36452 15408 36504 15428
rect 36504 15408 36506 15428
rect 36542 3440 36598 3496
rect 37278 14184 37334 14240
rect 37278 5344 37334 5400
rect 37186 4548 37242 4584
rect 37186 4528 37188 4548
rect 37188 4528 37240 4548
rect 37240 4528 37242 4548
rect 37094 2488 37150 2544
rect 38106 32444 38108 32464
rect 38108 32444 38160 32464
rect 38160 32444 38162 32464
rect 38106 32408 38162 32444
rect 38106 30776 38162 30832
rect 38106 29144 38162 29200
rect 38106 27512 38162 27568
rect 38106 25764 38162 25800
rect 38106 25744 38108 25764
rect 38108 25744 38160 25764
rect 38160 25744 38162 25764
rect 38014 24132 38070 24168
rect 38014 24112 38016 24132
rect 38016 24112 38068 24132
rect 38068 24112 38070 24132
rect 38106 22480 38162 22536
rect 38106 20848 38162 20904
rect 38106 19080 38162 19136
rect 38106 17448 38162 17504
rect 38014 15816 38070 15872
rect 38106 12416 38162 12472
rect 38106 10784 38162 10840
rect 38106 9152 38162 9208
rect 38106 7520 38162 7576
rect 38014 5752 38070 5808
rect 38106 856 38162 912
rect 39854 6160 39910 6216
<< metal3 >>
rect 35617 39130 35683 39133
rect 39200 39130 40000 39160
rect 35617 39128 40000 39130
rect 35617 39072 35622 39128
rect 35678 39072 40000 39128
rect 35617 39070 40000 39072
rect 35617 39067 35683 39070
rect 39200 39040 40000 39070
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 35801 37498 35867 37501
rect 39200 37498 40000 37528
rect 35801 37496 40000 37498
rect 35801 37440 35806 37496
rect 35862 37440 40000 37496
rect 35801 37438 40000 37440
rect 35801 37435 35867 37438
rect 39200 37408 40000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 20161 36956 20227 36957
rect 20110 36954 20116 36956
rect 20070 36894 20116 36954
rect 20180 36952 20227 36956
rect 20222 36896 20227 36952
rect 20110 36892 20116 36894
rect 20180 36892 20227 36896
rect 20161 36891 20227 36892
rect 36261 36548 36327 36549
rect 36261 36544 36308 36548
rect 36372 36546 36378 36548
rect 36261 36488 36266 36544
rect 36261 36484 36308 36488
rect 36372 36486 36418 36546
rect 36372 36484 36378 36486
rect 36261 36483 36327 36484
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 12249 36410 12315 36413
rect 30097 36410 30163 36413
rect 12249 36408 30163 36410
rect 12249 36352 12254 36408
rect 12310 36352 30102 36408
rect 30158 36352 30163 36408
rect 12249 36350 30163 36352
rect 12249 36347 12315 36350
rect 30097 36347 30163 36350
rect 7465 36274 7531 36277
rect 30189 36274 30255 36277
rect 7465 36272 30255 36274
rect 7465 36216 7470 36272
rect 7526 36216 30194 36272
rect 30250 36216 30255 36272
rect 7465 36214 30255 36216
rect 7465 36211 7531 36214
rect 30189 36211 30255 36214
rect 9213 36138 9279 36141
rect 28993 36138 29059 36141
rect 9213 36136 29059 36138
rect 9213 36080 9218 36136
rect 9274 36080 28998 36136
rect 29054 36080 29059 36136
rect 9213 36078 29059 36080
rect 9213 36075 9279 36078
rect 28993 36075 29059 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 36721 35866 36787 35869
rect 39200 35866 40000 35896
rect 36721 35864 40000 35866
rect 36721 35808 36726 35864
rect 36782 35808 40000 35864
rect 36721 35806 40000 35808
rect 36721 35803 36787 35806
rect 39200 35776 40000 35806
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 34646 34580 34652 34644
rect 34716 34642 34722 34644
rect 35249 34642 35315 34645
rect 34716 34640 35315 34642
rect 34716 34584 35254 34640
rect 35310 34584 35315 34640
rect 34716 34582 35315 34584
rect 34716 34580 34722 34582
rect 35249 34579 35315 34582
rect 22369 34372 22435 34373
rect 22318 34308 22324 34372
rect 22388 34370 22435 34372
rect 22388 34368 22480 34370
rect 22430 34312 22480 34368
rect 22388 34310 22480 34312
rect 22388 34308 22435 34310
rect 22369 34307 22435 34308
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 35801 34234 35867 34237
rect 39200 34234 40000 34264
rect 35801 34232 40000 34234
rect 35801 34176 35806 34232
rect 35862 34176 40000 34232
rect 35801 34174 40000 34176
rect 35801 34171 35867 34174
rect 39200 34144 40000 34174
rect 34462 33764 34468 33828
rect 34532 33826 34538 33828
rect 34605 33826 34671 33829
rect 34532 33824 34671 33826
rect 34532 33768 34610 33824
rect 34666 33768 34671 33824
rect 34532 33766 34671 33768
rect 34532 33764 34538 33766
rect 34605 33763 34671 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 38101 32466 38167 32469
rect 39200 32466 40000 32496
rect 38101 32464 40000 32466
rect 38101 32408 38106 32464
rect 38162 32408 40000 32464
rect 38101 32406 40000 32408
rect 38101 32403 38167 32406
rect 39200 32376 40000 32406
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 38101 30834 38167 30837
rect 39200 30834 40000 30864
rect 38101 30832 40000 30834
rect 38101 30776 38106 30832
rect 38162 30776 40000 30832
rect 38101 30774 40000 30776
rect 38101 30771 38167 30774
rect 39200 30744 40000 30774
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 38101 29202 38167 29205
rect 39200 29202 40000 29232
rect 38101 29200 40000 29202
rect 38101 29144 38106 29200
rect 38162 29144 40000 29200
rect 38101 29142 40000 29144
rect 38101 29139 38167 29142
rect 39200 29112 40000 29142
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 38101 27570 38167 27573
rect 39200 27570 40000 27600
rect 38101 27568 40000 27570
rect 38101 27512 38106 27568
rect 38162 27512 40000 27568
rect 38101 27510 40000 27512
rect 38101 27507 38167 27510
rect 39200 27480 40000 27510
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 38101 25802 38167 25805
rect 39200 25802 40000 25832
rect 38101 25800 40000 25802
rect 38101 25744 38106 25800
rect 38162 25744 40000 25800
rect 38101 25742 40000 25744
rect 38101 25739 38167 25742
rect 39200 25712 40000 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 38009 24170 38075 24173
rect 39200 24170 40000 24200
rect 38009 24168 40000 24170
rect 38009 24112 38014 24168
rect 38070 24112 40000 24168
rect 38009 24110 40000 24112
rect 38009 24107 38075 24110
rect 39200 24080 40000 24110
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 38101 22538 38167 22541
rect 39200 22538 40000 22568
rect 38101 22536 40000 22538
rect 38101 22480 38106 22536
rect 38162 22480 40000 22536
rect 38101 22478 40000 22480
rect 38101 22475 38167 22478
rect 39200 22448 40000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 15510 21252 15516 21316
rect 15580 21314 15586 21316
rect 29913 21314 29979 21317
rect 15580 21312 29979 21314
rect 15580 21256 29918 21312
rect 29974 21256 29979 21312
rect 15580 21254 29979 21256
rect 15580 21252 15586 21254
rect 29913 21251 29979 21254
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 38101 20906 38167 20909
rect 39200 20906 40000 20936
rect 38101 20904 40000 20906
rect 38101 20848 38106 20904
rect 38162 20848 40000 20904
rect 38101 20846 40000 20848
rect 38101 20843 38167 20846
rect 39200 20816 40000 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 38101 19138 38167 19141
rect 39200 19138 40000 19168
rect 38101 19136 40000 19138
rect 38101 19080 38106 19136
rect 38162 19080 40000 19136
rect 38101 19078 40000 19080
rect 38101 19075 38167 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 39200 19048 40000 19078
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 38101 17506 38167 17509
rect 39200 17506 40000 17536
rect 38101 17504 40000 17506
rect 38101 17448 38106 17504
rect 38162 17448 40000 17504
rect 38101 17446 40000 17448
rect 38101 17443 38167 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 39200 17416 40000 17446
rect 19568 17375 19888 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 38009 15874 38075 15877
rect 39200 15874 40000 15904
rect 38009 15872 40000 15874
rect 38009 15816 38014 15872
rect 38070 15816 40000 15872
rect 38009 15814 40000 15816
rect 38009 15811 38075 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 39200 15784 40000 15814
rect 34928 15743 35248 15744
rect 20110 15404 20116 15468
rect 20180 15466 20186 15468
rect 36445 15466 36511 15469
rect 20180 15464 36511 15466
rect 20180 15408 36450 15464
rect 36506 15408 36511 15464
rect 20180 15406 36511 15408
rect 20180 15404 20186 15406
rect 36445 15403 36511 15406
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 10726 14860 10732 14924
rect 10796 14922 10802 14924
rect 23657 14922 23723 14925
rect 10796 14920 23723 14922
rect 10796 14864 23662 14920
rect 23718 14864 23723 14920
rect 10796 14862 23723 14864
rect 10796 14860 10802 14862
rect 23657 14859 23723 14862
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 37273 14242 37339 14245
rect 39200 14242 40000 14272
rect 37273 14240 40000 14242
rect 37273 14184 37278 14240
rect 37334 14184 40000 14240
rect 37273 14182 40000 14184
rect 37273 14179 37339 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 39200 14152 40000 14182
rect 19568 14111 19888 14112
rect 11646 13908 11652 13972
rect 11716 13970 11722 13972
rect 24301 13970 24367 13973
rect 11716 13968 24367 13970
rect 11716 13912 24306 13968
rect 24362 13912 24367 13968
rect 11716 13910 24367 13912
rect 11716 13908 11722 13910
rect 24301 13907 24367 13910
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 10910 13228 10916 13292
rect 10980 13290 10986 13292
rect 22277 13290 22343 13293
rect 23197 13290 23263 13293
rect 10980 13288 23263 13290
rect 10980 13232 22282 13288
rect 22338 13232 23202 13288
rect 23258 13232 23263 13288
rect 10980 13230 23263 13232
rect 10980 13228 10986 13230
rect 22277 13227 22343 13230
rect 23197 13227 23263 13230
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 38101 12474 38167 12477
rect 39200 12474 40000 12504
rect 38101 12472 40000 12474
rect 38101 12416 38106 12472
rect 38162 12416 40000 12472
rect 38101 12414 40000 12416
rect 38101 12411 38167 12414
rect 39200 12384 40000 12414
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 38101 10842 38167 10845
rect 39200 10842 40000 10872
rect 38101 10840 40000 10842
rect 38101 10784 38106 10840
rect 38162 10784 40000 10840
rect 38101 10782 40000 10784
rect 38101 10779 38167 10782
rect 39200 10752 40000 10782
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 0 10026 800 10056
rect 3417 10026 3483 10029
rect 0 10024 3483 10026
rect 0 9968 3422 10024
rect 3478 9968 3483 10024
rect 0 9966 3483 9968
rect 0 9936 800 9966
rect 3417 9963 3483 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 38101 9210 38167 9213
rect 39200 9210 40000 9240
rect 38101 9208 40000 9210
rect 38101 9152 38106 9208
rect 38162 9152 40000 9208
rect 38101 9150 40000 9152
rect 38101 9147 38167 9150
rect 39200 9120 40000 9150
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 1945 8394 2011 8397
rect 23473 8394 23539 8397
rect 1945 8392 23539 8394
rect 1945 8336 1950 8392
rect 2006 8336 23478 8392
rect 23534 8336 23539 8392
rect 1945 8334 23539 8336
rect 1945 8331 2011 8334
rect 23473 8331 23539 8334
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 9949 7850 10015 7853
rect 28809 7850 28875 7853
rect 9949 7848 28875 7850
rect 9949 7792 9954 7848
rect 10010 7792 28814 7848
rect 28870 7792 28875 7848
rect 9949 7790 28875 7792
rect 9949 7787 10015 7790
rect 28809 7787 28875 7790
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 38101 7578 38167 7581
rect 39200 7578 40000 7608
rect 38101 7576 40000 7578
rect 38101 7520 38106 7576
rect 38162 7520 40000 7576
rect 38101 7518 40000 7520
rect 38101 7515 38167 7518
rect 39200 7488 40000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 12065 6218 12131 6221
rect 31201 6218 31267 6221
rect 12065 6216 31267 6218
rect 12065 6160 12070 6216
rect 12126 6160 31206 6216
rect 31262 6160 31267 6216
rect 12065 6158 31267 6160
rect 12065 6155 12131 6158
rect 31201 6155 31267 6158
rect 35249 6218 35315 6221
rect 39849 6218 39915 6221
rect 35249 6216 39915 6218
rect 35249 6160 35254 6216
rect 35310 6160 39854 6216
rect 39910 6160 39915 6216
rect 35249 6158 39915 6160
rect 35249 6155 35315 6158
rect 39849 6155 39915 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 38009 5810 38075 5813
rect 39200 5810 40000 5840
rect 38009 5808 40000 5810
rect 38009 5752 38014 5808
rect 38070 5752 40000 5808
rect 38009 5750 40000 5752
rect 38009 5747 38075 5750
rect 39200 5720 40000 5750
rect 4705 5674 4771 5677
rect 4838 5674 4844 5676
rect 4705 5672 4844 5674
rect 4705 5616 4710 5672
rect 4766 5616 4844 5672
rect 4705 5614 4844 5616
rect 4705 5611 4771 5614
rect 4838 5612 4844 5614
rect 4908 5612 4914 5676
rect 34646 5476 34652 5540
rect 34716 5538 34722 5540
rect 34881 5538 34947 5541
rect 34716 5536 34947 5538
rect 34716 5480 34886 5536
rect 34942 5480 34947 5536
rect 34716 5478 34947 5480
rect 34716 5476 34722 5478
rect 34881 5475 34947 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 22645 5402 22711 5405
rect 37273 5402 37339 5405
rect 22645 5400 37339 5402
rect 22645 5344 22650 5400
rect 22706 5344 37278 5400
rect 37334 5344 37339 5400
rect 22645 5342 37339 5344
rect 22645 5339 22711 5342
rect 37273 5339 37339 5342
rect 30649 5266 30715 5269
rect 36302 5266 36308 5268
rect 30649 5264 36308 5266
rect 30649 5208 30654 5264
rect 30710 5208 36308 5264
rect 30649 5206 36308 5208
rect 30649 5203 30715 5206
rect 36302 5204 36308 5206
rect 36372 5204 36378 5268
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 33501 4858 33567 4861
rect 34462 4858 34468 4860
rect 33501 4856 34468 4858
rect 33501 4800 33506 4856
rect 33562 4800 34468 4856
rect 33501 4798 34468 4800
rect 33501 4795 33567 4798
rect 34462 4796 34468 4798
rect 34532 4796 34538 4860
rect 18505 4586 18571 4589
rect 37181 4586 37247 4589
rect 18505 4584 37247 4586
rect 18505 4528 18510 4584
rect 18566 4528 37186 4584
rect 37242 4528 37247 4584
rect 18505 4526 37247 4528
rect 18505 4523 18571 4526
rect 37181 4523 37247 4526
rect 3877 4452 3943 4453
rect 3877 4450 3924 4452
rect 3832 4448 3924 4450
rect 3832 4392 3882 4448
rect 3832 4390 3924 4392
rect 3877 4388 3924 4390
rect 3988 4388 3994 4452
rect 20805 4450 20871 4453
rect 28717 4450 28783 4453
rect 20805 4448 28783 4450
rect 20805 4392 20810 4448
rect 20866 4392 28722 4448
rect 28778 4392 28783 4448
rect 20805 4390 28783 4392
rect 3877 4387 3943 4388
rect 20805 4387 20871 4390
rect 28717 4387 28783 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 23933 4314 23999 4317
rect 32857 4314 32923 4317
rect 23933 4312 32923 4314
rect 23933 4256 23938 4312
rect 23994 4256 32862 4312
rect 32918 4256 32923 4312
rect 23933 4254 32923 4256
rect 23933 4251 23999 4254
rect 32857 4251 32923 4254
rect 9213 4178 9279 4181
rect 22093 4178 22159 4181
rect 9213 4176 22159 4178
rect 9213 4120 9218 4176
rect 9274 4120 22098 4176
rect 22154 4120 22159 4176
rect 9213 4118 22159 4120
rect 9213 4115 9279 4118
rect 22093 4115 22159 4118
rect 29729 4178 29795 4181
rect 30741 4178 30807 4181
rect 29729 4176 30807 4178
rect 29729 4120 29734 4176
rect 29790 4120 30746 4176
rect 30802 4120 30807 4176
rect 29729 4118 30807 4120
rect 29729 4115 29795 4118
rect 30741 4115 30807 4118
rect 35801 4178 35867 4181
rect 39200 4178 40000 4208
rect 35801 4176 40000 4178
rect 35801 4120 35806 4176
rect 35862 4120 40000 4176
rect 35801 4118 40000 4120
rect 35801 4115 35867 4118
rect 39200 4088 40000 4118
rect 10593 4042 10659 4045
rect 10726 4042 10732 4044
rect 10593 4040 10732 4042
rect 10593 3984 10598 4040
rect 10654 3984 10732 4040
rect 10593 3982 10732 3984
rect 10593 3979 10659 3982
rect 10726 3980 10732 3982
rect 10796 3980 10802 4044
rect 11513 4042 11579 4045
rect 11646 4042 11652 4044
rect 11513 4040 11652 4042
rect 11513 3984 11518 4040
rect 11574 3984 11652 4040
rect 11513 3982 11652 3984
rect 11513 3979 11579 3982
rect 11646 3980 11652 3982
rect 11716 3980 11722 4044
rect 12065 4042 12131 4045
rect 19057 4042 19123 4045
rect 20621 4042 20687 4045
rect 12065 4040 20687 4042
rect 12065 3984 12070 4040
rect 12126 3984 19062 4040
rect 19118 3984 20626 4040
rect 20682 3984 20687 4040
rect 12065 3982 20687 3984
rect 12065 3979 12131 3982
rect 19057 3979 19123 3982
rect 20621 3979 20687 3982
rect 8477 3906 8543 3909
rect 19885 3906 19951 3909
rect 8477 3904 19951 3906
rect 8477 3848 8482 3904
rect 8538 3848 19890 3904
rect 19946 3848 19951 3904
rect 8477 3846 19951 3848
rect 8477 3843 8543 3846
rect 19885 3843 19951 3846
rect 23013 3906 23079 3909
rect 34145 3906 34211 3909
rect 23013 3904 34211 3906
rect 23013 3848 23018 3904
rect 23074 3848 34150 3904
rect 34206 3848 34211 3904
rect 23013 3846 34211 3848
rect 23013 3843 23079 3846
rect 34145 3843 34211 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 6085 3770 6151 3773
rect 29545 3770 29611 3773
rect 6085 3768 29611 3770
rect 6085 3712 6090 3768
rect 6146 3712 29550 3768
rect 29606 3712 29611 3768
rect 6085 3710 29611 3712
rect 6085 3707 6151 3710
rect 29545 3707 29611 3710
rect 8293 3634 8359 3637
rect 12065 3634 12131 3637
rect 8293 3632 12131 3634
rect 8293 3576 8298 3632
rect 8354 3576 12070 3632
rect 12126 3576 12131 3632
rect 8293 3574 12131 3576
rect 8293 3571 8359 3574
rect 12065 3571 12131 3574
rect 16849 3634 16915 3637
rect 22318 3634 22324 3636
rect 16849 3632 22324 3634
rect 16849 3576 16854 3632
rect 16910 3576 22324 3632
rect 16849 3574 22324 3576
rect 16849 3571 16915 3574
rect 22318 3572 22324 3574
rect 22388 3572 22394 3636
rect 23381 3634 23447 3637
rect 33501 3634 33567 3637
rect 23381 3632 33567 3634
rect 23381 3576 23386 3632
rect 23442 3576 33506 3632
rect 33562 3576 33567 3632
rect 23381 3574 33567 3576
rect 23381 3571 23447 3574
rect 33501 3571 33567 3574
rect 10961 3498 11027 3501
rect 6870 3496 11027 3498
rect 6870 3440 10966 3496
rect 11022 3440 11027 3496
rect 6870 3438 11027 3440
rect 4153 3362 4219 3365
rect 6870 3362 6930 3438
rect 10961 3435 11027 3438
rect 11329 3498 11395 3501
rect 23289 3498 23355 3501
rect 11329 3496 23355 3498
rect 11329 3440 11334 3496
rect 11390 3440 23294 3496
rect 23350 3440 23355 3496
rect 11329 3438 23355 3440
rect 11329 3435 11395 3438
rect 23289 3435 23355 3438
rect 24761 3498 24827 3501
rect 36537 3498 36603 3501
rect 24761 3496 36603 3498
rect 24761 3440 24766 3496
rect 24822 3440 36542 3496
rect 36598 3440 36603 3496
rect 24761 3438 36603 3440
rect 24761 3435 24827 3438
rect 36537 3435 36603 3438
rect 4153 3360 6930 3362
rect 4153 3304 4158 3360
rect 4214 3304 6930 3360
rect 4153 3302 6930 3304
rect 8201 3362 8267 3365
rect 11053 3362 11119 3365
rect 17493 3362 17559 3365
rect 8201 3360 11119 3362
rect 8201 3304 8206 3360
rect 8262 3304 11058 3360
rect 11114 3304 11119 3360
rect 8201 3302 11119 3304
rect 4153 3299 4219 3302
rect 8201 3299 8267 3302
rect 11053 3299 11119 3302
rect 11654 3360 17559 3362
rect 11654 3304 17498 3360
rect 17554 3304 17559 3360
rect 11654 3302 17559 3304
rect 4889 3226 4955 3229
rect 11654 3226 11714 3302
rect 17493 3299 17559 3302
rect 25589 3362 25655 3365
rect 33961 3362 34027 3365
rect 25589 3360 34027 3362
rect 25589 3304 25594 3360
rect 25650 3304 33966 3360
rect 34022 3304 34027 3360
rect 25589 3302 34027 3304
rect 25589 3299 25655 3302
rect 33961 3299 34027 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 4889 3224 11714 3226
rect 4889 3168 4894 3224
rect 4950 3168 11714 3224
rect 4889 3166 11714 3168
rect 15377 3226 15443 3229
rect 15510 3226 15516 3228
rect 15377 3224 15516 3226
rect 15377 3168 15382 3224
rect 15438 3168 15516 3224
rect 15377 3166 15516 3168
rect 4889 3163 4955 3166
rect 15377 3163 15443 3166
rect 15510 3164 15516 3166
rect 15580 3164 15586 3228
rect 14549 3090 14615 3093
rect 27337 3090 27403 3093
rect 14549 3088 27403 3090
rect 14549 3032 14554 3088
rect 14610 3032 27342 3088
rect 27398 3032 27403 3088
rect 14549 3030 27403 3032
rect 14549 3027 14615 3030
rect 27337 3027 27403 3030
rect 5533 2954 5599 2957
rect 27521 2954 27587 2957
rect 5533 2952 27587 2954
rect 5533 2896 5538 2952
rect 5594 2896 27526 2952
rect 27582 2896 27587 2952
rect 5533 2894 27587 2896
rect 5533 2891 5599 2894
rect 27521 2891 27587 2894
rect 10501 2818 10567 2821
rect 12433 2818 12499 2821
rect 10501 2816 12499 2818
rect 10501 2760 10506 2816
rect 10562 2760 12438 2816
rect 12494 2760 12499 2816
rect 10501 2758 12499 2760
rect 10501 2755 10567 2758
rect 12433 2755 12499 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 10777 2682 10843 2685
rect 10910 2682 10916 2684
rect 10777 2680 10916 2682
rect 10777 2624 10782 2680
rect 10838 2624 10916 2680
rect 10777 2622 10916 2624
rect 10777 2619 10843 2622
rect 10910 2620 10916 2622
rect 10980 2620 10986 2684
rect 4838 2484 4844 2548
rect 4908 2546 4914 2548
rect 28073 2546 28139 2549
rect 4908 2544 28139 2546
rect 4908 2488 28078 2544
rect 28134 2488 28139 2544
rect 4908 2486 28139 2488
rect 4908 2484 4914 2486
rect 28073 2483 28139 2486
rect 37089 2546 37155 2549
rect 39200 2546 40000 2576
rect 37089 2544 40000 2546
rect 37089 2488 37094 2544
rect 37150 2488 40000 2544
rect 37089 2486 40000 2488
rect 37089 2483 37155 2486
rect 39200 2456 40000 2486
rect 3417 2410 3483 2413
rect 27337 2410 27403 2413
rect 3417 2408 27403 2410
rect 3417 2352 3422 2408
rect 3478 2352 27342 2408
rect 27398 2352 27403 2408
rect 3417 2350 27403 2352
rect 3417 2347 3483 2350
rect 27337 2347 27403 2350
rect 20621 2274 20687 2277
rect 33409 2274 33475 2277
rect 20621 2272 33475 2274
rect 20621 2216 20626 2272
rect 20682 2216 33414 2272
rect 33470 2216 33475 2272
rect 20621 2214 33475 2216
rect 20621 2211 20687 2214
rect 33409 2211 33475 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3918 1940 3924 2004
rect 3988 2002 3994 2004
rect 24853 2002 24919 2005
rect 3988 2000 24919 2002
rect 3988 1944 24858 2000
rect 24914 1944 24919 2000
rect 3988 1942 24919 1944
rect 3988 1940 3994 1942
rect 24853 1939 24919 1942
rect 15009 1866 15075 1869
rect 25497 1866 25563 1869
rect 15009 1864 25563 1866
rect 15009 1808 15014 1864
rect 15070 1808 25502 1864
rect 25558 1808 25563 1864
rect 15009 1806 25563 1808
rect 15009 1803 15075 1806
rect 25497 1803 25563 1806
rect 14273 1730 14339 1733
rect 25221 1730 25287 1733
rect 14273 1728 25287 1730
rect 14273 1672 14278 1728
rect 14334 1672 25226 1728
rect 25282 1672 25287 1728
rect 14273 1670 25287 1672
rect 14273 1667 14339 1670
rect 25221 1667 25287 1670
rect 8385 1594 8451 1597
rect 20437 1594 20503 1597
rect 8385 1592 20503 1594
rect 8385 1536 8390 1592
rect 8446 1536 20442 1592
rect 20498 1536 20503 1592
rect 8385 1534 20503 1536
rect 8385 1531 8451 1534
rect 20437 1531 20503 1534
rect 38101 914 38167 917
rect 39200 914 40000 944
rect 38101 912 40000 914
rect 38101 856 38106 912
rect 38162 856 40000 912
rect 38101 854 40000 856
rect 38101 851 38167 854
rect 39200 824 40000 854
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 20116 36952 20180 36956
rect 20116 36896 20166 36952
rect 20166 36896 20180 36952
rect 20116 36892 20180 36896
rect 36308 36544 36372 36548
rect 36308 36488 36322 36544
rect 36322 36488 36372 36544
rect 36308 36484 36372 36488
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 34652 34580 34716 34644
rect 22324 34368 22388 34372
rect 22324 34312 22374 34368
rect 22374 34312 22388 34368
rect 22324 34308 22388 34312
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 34468 33764 34532 33828
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 15516 21252 15580 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 20116 15404 20180 15468
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 10732 14860 10796 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 11652 13908 11716 13972
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 10916 13228 10980 13292
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4844 5612 4908 5676
rect 34652 5476 34716 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 36308 5204 36372 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 34468 4796 34532 4860
rect 3924 4448 3988 4452
rect 3924 4392 3938 4448
rect 3938 4392 3988 4448
rect 3924 4388 3988 4392
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 10732 3980 10796 4044
rect 11652 3980 11716 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 22324 3572 22388 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 15516 3164 15580 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 10916 2620 10980 2684
rect 4844 2484 4908 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 3924 1940 3988 2004
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 20115 36956 20181 36957
rect 20115 36892 20116 36956
rect 20180 36892 20181 36956
rect 20115 36891 20181 36892
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 15515 21316 15581 21317
rect 15515 21252 15516 21316
rect 15580 21252 15581 21316
rect 15515 21251 15581 21252
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 10731 14924 10797 14925
rect 10731 14860 10732 14924
rect 10796 14860 10797 14924
rect 10731 14859 10797 14860
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4843 5676 4909 5677
rect 4843 5612 4844 5676
rect 4908 5612 4909 5676
rect 4843 5611 4909 5612
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 3923 4452 3989 4453
rect 3923 4388 3924 4452
rect 3988 4388 3989 4452
rect 3923 4387 3989 4388
rect 3926 2005 3986 4387
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4846 2549 4906 5611
rect 10734 4045 10794 14859
rect 11651 13972 11717 13973
rect 11651 13908 11652 13972
rect 11716 13908 11717 13972
rect 11651 13907 11717 13908
rect 10915 13292 10981 13293
rect 10915 13228 10916 13292
rect 10980 13228 10981 13292
rect 10915 13227 10981 13228
rect 10731 4044 10797 4045
rect 10731 3980 10732 4044
rect 10796 3980 10797 4044
rect 10731 3979 10797 3980
rect 10918 2685 10978 13227
rect 11654 4045 11714 13907
rect 11651 4044 11717 4045
rect 11651 3980 11652 4044
rect 11716 3980 11717 4044
rect 11651 3979 11717 3980
rect 15518 3229 15578 21251
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 20118 15469 20178 36891
rect 34928 36480 35248 37504
rect 36307 36548 36373 36549
rect 36307 36484 36308 36548
rect 36372 36484 36373 36548
rect 36307 36483 36373 36484
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34651 34644 34717 34645
rect 34651 34580 34652 34644
rect 34716 34580 34717 34644
rect 34651 34579 34717 34580
rect 22323 34372 22389 34373
rect 22323 34308 22324 34372
rect 22388 34308 22389 34372
rect 22323 34307 22389 34308
rect 20115 15468 20181 15469
rect 20115 15404 20116 15468
rect 20180 15404 20181 15468
rect 20115 15403 20181 15404
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 22326 3637 22386 34307
rect 34467 33828 34533 33829
rect 34467 33764 34468 33828
rect 34532 33764 34533 33828
rect 34467 33763 34533 33764
rect 34470 4861 34530 33763
rect 34654 5541 34714 34579
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34651 5540 34717 5541
rect 34651 5476 34652 5540
rect 34716 5476 34717 5540
rect 34651 5475 34717 5476
rect 34928 4928 35248 5952
rect 36310 5269 36370 36483
rect 36307 5268 36373 5269
rect 36307 5204 36308 5268
rect 36372 5204 36373 5268
rect 36307 5203 36373 5204
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34467 4860 34533 4861
rect 34467 4796 34468 4860
rect 34532 4796 34533 4860
rect 34467 4795 34533 4796
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 22323 3636 22389 3637
rect 22323 3572 22324 3636
rect 22388 3572 22389 3636
rect 22323 3571 22389 3572
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 15515 3228 15581 3229
rect 15515 3164 15516 3228
rect 15580 3164 15581 3228
rect 15515 3163 15581 3164
rect 10915 2684 10981 2685
rect 10915 2620 10916 2684
rect 10980 2620 10981 2684
rect 10915 2619 10981 2620
rect 4843 2548 4909 2549
rect 4843 2484 4844 2548
rect 4908 2484 4909 2548
rect 4843 2483 4909 2484
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 3923 2004 3989 2005
rect 3923 1940 3924 2004
rect 3988 1940 3989 2004
rect 3923 1939 3989 1940
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1644511149
transform -1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B
timestamp 1644511149
transform 1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__B
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__B
timestamp 1644511149
transform -1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1644511149
transform -1 0 24564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1644511149
transform -1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1644511149
transform -1 0 23368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__B
timestamp 1644511149
transform -1 0 32568 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__B
timestamp 1644511149
transform -1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A_N
timestamp 1644511149
transform -1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B
timestamp 1644511149
transform -1 0 21712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A_N
timestamp 1644511149
transform 1 0 24472 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A_N
timestamp 1644511149
transform -1 0 29716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__B
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A_N
timestamp 1644511149
transform 1 0 24840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B
timestamp 1644511149
transform 1 0 23368 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B
timestamp 1644511149
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__B
timestamp 1644511149
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1644511149
transform -1 0 26496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B
timestamp 1644511149
transform -1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1644511149
transform -1 0 26496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__B
timestamp 1644511149
transform -1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1644511149
transform -1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 1644511149
transform -1 0 27140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__B
timestamp 1644511149
transform 1 0 27876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B
timestamp 1644511149
transform -1 0 27968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B
timestamp 1644511149
transform -1 0 31280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A_N
timestamp 1644511149
transform 1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__B
timestamp 1644511149
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1644511149
transform -1 0 34224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B
timestamp 1644511149
transform -1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B
timestamp 1644511149
transform -1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1644511149
transform -1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A_N
timestamp 1644511149
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__B
timestamp 1644511149
transform -1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1644511149
transform -1 0 36708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B
timestamp 1644511149
transform 1 0 35052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A_N
timestamp 1644511149
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1644511149
transform -1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__S
timestamp 1644511149
transform 1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1644511149
transform 1 0 3956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A0
timestamp 1644511149
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A0
timestamp 1644511149
transform -1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A0
timestamp 1644511149
transform -1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A0
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A0
timestamp 1644511149
transform -1 0 30176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A0
timestamp 1644511149
transform -1 0 32384 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A0
timestamp 1644511149
transform -1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1644511149
transform 1 0 12880 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1644511149
transform -1 0 34224 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A0
timestamp 1644511149
transform -1 0 13524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__S
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A0
timestamp 1644511149
transform -1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A0
timestamp 1644511149
transform -1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A0
timestamp 1644511149
transform -1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__S
timestamp 1644511149
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A0
timestamp 1644511149
transform -1 0 38180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A_N
timestamp 1644511149
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1644511149
transform -1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A0
timestamp 1644511149
transform -1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__S
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1644511149
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1644511149
transform -1 0 23920 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1644511149
transform -1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A0
timestamp 1644511149
transform -1 0 26680 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A0
timestamp 1644511149
transform -1 0 29072 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__B
timestamp 1644511149
transform -1 0 22448 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A0
timestamp 1644511149
transform 1 0 31464 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__B
timestamp 1644511149
transform -1 0 29716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A0
timestamp 1644511149
transform 1 0 33396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__S
timestamp 1644511149
transform -1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__S
timestamp 1644511149
transform -1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S
timestamp 1644511149
transform -1 0 23000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A_N
timestamp 1644511149
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1644511149
transform -1 0 3956 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1644511149
transform 1 0 11040 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A_N
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__B
timestamp 1644511149
transform 1 0 23552 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__B
timestamp 1644511149
transform -1 0 27876 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__B1
timestamp 1644511149
transform -1 0 31004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__B1
timestamp 1644511149
transform 1 0 31464 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1644511149
transform 1 0 26496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1644511149
transform -1 0 5888 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__B
timestamp 1644511149
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__B
timestamp 1644511149
transform -1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B
timestamp 1644511149
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1644511149
transform -1 0 4968 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__B
timestamp 1644511149
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1644511149
transform 1 0 7084 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__B
timestamp 1644511149
transform -1 0 30176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1644511149
transform -1 0 8188 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1644511149
transform -1 0 31372 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__B
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1644511149
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1644511149
transform 1 0 32936 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1644511149
transform 1 0 15640 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__B
timestamp 1644511149
transform -1 0 14812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1644511149
transform -1 0 15272 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__B
timestamp 1644511149
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1644511149
transform 1 0 14444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__B
timestamp 1644511149
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1644511149
transform -1 0 17112 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1644511149
transform -1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__B
timestamp 1644511149
transform -1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1644511149
transform -1 0 18124 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1644511149
transform 1 0 19688 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__B
timestamp 1644511149
transform -1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1644511149
transform 1 0 20700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1644511149
transform 1 0 11592 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1644511149
transform 1 0 13432 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1644511149
transform -1 0 15824 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1644511149
transform -1 0 16560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__B
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__B
timestamp 1644511149
transform -1 0 25760 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__B
timestamp 1644511149
transform -1 0 27600 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__B
timestamp 1644511149
transform -1 0 29900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1644511149
transform -1 0 24748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1644511149
transform 1 0 28244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1644511149
transform -1 0 35512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__B1
timestamp 1644511149
transform 1 0 33396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1644511149
transform 1 0 31464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__B1
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1644511149
transform 1 0 25668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__B1
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1644511149
transform 1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__B1_N
timestamp 1644511149
transform 1 0 9108 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__C1
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__B1
timestamp 1644511149
transform -1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1644511149
transform -1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1644511149
transform 1 0 6164 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1644511149
transform 1 0 5888 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1644511149
transform 1 0 5428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A
timestamp 1644511149
transform 1 0 7360 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__B1
timestamp 1644511149
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__A
timestamp 1644511149
transform 1 0 16008 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__B1
timestamp 1644511149
transform 1 0 19964 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__A
timestamp 1644511149
transform -1 0 23644 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__B1
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1644511149
transform 1 0 29624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1644511149
transform 1 0 27600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1644511149
transform -1 0 27784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1644511149
transform -1 0 23828 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1644511149
transform 1 0 16744 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1644511149
transform 1 0 15364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1644511149
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1644511149
transform 1 0 10488 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1644511149
transform 1 0 8372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1644511149
transform 1 0 3864 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1644511149
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1644511149
transform -1 0 8924 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1644511149
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1644511149
transform 1 0 4140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1644511149
transform 1 0 11224 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1644511149
transform 1 0 10488 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1644511149
transform 1 0 13524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1644511149
transform 1 0 17480 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1644511149
transform 1 0 35604 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1644511149
transform 1 0 33764 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1644511149
transform 1 0 35144 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__A
timestamp 1644511149
transform 1 0 2024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A
timestamp 1644511149
transform -1 0 29440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__A
timestamp 1644511149
transform 1 0 31188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A
timestamp 1644511149
transform -1 0 36156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__A
timestamp 1644511149
transform 1 0 36432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__A
timestamp 1644511149
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1644511149
transform -1 0 28796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1644511149
transform -1 0 38180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A
timestamp 1644511149
transform -1 0 38180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A
timestamp 1644511149
transform -1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__A
timestamp 1644511149
transform -1 0 37628 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__A
timestamp 1644511149
transform 1 0 37444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1644511149
transform -1 0 37628 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__A
timestamp 1644511149
transform 1 0 35880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1644511149
transform 1 0 10856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1644511149
transform -1 0 28336 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 33028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 33856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 34684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 35144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 36340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 34132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 33304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 36800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 28152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 28704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 28796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 29072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 29716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 30544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 32108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 34868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 25116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 32936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 34868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 36248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 37628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 36616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 35696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 35696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 27600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 28152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform -1 0 31096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 31648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 29992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 32292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 30728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 32752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 19688 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 20516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 21160 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 24380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 12420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 9476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 18308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 19044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 20516 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 21344 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 22172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1644511149
transform -1 0 23092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1644511149
transform -1 0 24656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1644511149
transform -1 0 23828 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1644511149
transform -1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1644511149
transform -1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1644511149
transform -1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1644511149
transform -1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1644511149
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1644511149
transform -1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1644511149
transform -1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1644511149
transform -1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1644511149
transform -1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1644511149
transform -1 0 1748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1644511149
transform -1 0 12328 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1644511149
transform -1 0 15180 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1644511149
transform -1 0 12880 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1644511149
transform -1 0 16100 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1644511149
transform -1 0 18584 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1644511149
transform -1 0 17664 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1644511149
transform -1 0 17020 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1644511149
transform -1 0 18216 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1644511149
transform -1 0 19412 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1644511149
transform -1 0 20148 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1644511149
transform -1 0 2300 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1644511149
transform -1 0 23828 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1644511149
transform -1 0 22632 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1644511149
transform -1 0 23920 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1644511149
transform -1 0 24472 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1644511149
transform -1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1644511149
transform -1 0 26036 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1644511149
transform -1 0 28980 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1644511149
transform -1 0 29716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1644511149
transform -1 0 31372 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1644511149
transform -1 0 29992 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1644511149
transform -1 0 2668 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1644511149
transform -1 0 34132 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1644511149
transform -1 0 33672 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1644511149
transform -1 0 35604 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1644511149
transform -1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1644511149
transform -1 0 38180 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1644511149
transform -1 0 37444 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1644511149
transform -1 0 37444 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1644511149
transform -1 0 37444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1644511149
transform -1 0 4692 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1644511149
transform -1 0 5244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1644511149
transform -1 0 6348 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1644511149
transform -1 0 6900 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1644511149
transform -1 0 10212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1644511149
transform -1 0 11684 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1644511149
transform -1 0 10028 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1644511149
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1644511149
transform -1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1644511149
transform -1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1644511149
transform -1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1644511149
transform -1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1644511149
transform -1 0 8096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1644511149
transform -1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1644511149
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1644511149
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1644511149
transform -1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1644511149
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1644511149
transform -1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1644511149
transform -1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1644511149
transform -1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1644511149
transform -1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1644511149
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1644511149
transform -1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1644511149
transform -1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1644511149
transform -1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1644511149
transform -1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1644511149
transform -1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1644511149
transform -1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1644511149
transform -1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1644511149
transform -1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1644511149
transform -1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1644511149
transform -1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1644511149
transform -1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1644511149
transform -1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1644511149
transform -1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1644511149
transform -1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1644511149
transform -1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input146_A
timestamp 1644511149
transform -1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input147_A
timestamp 1644511149
transform -1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input148_A
timestamp 1644511149
transform -1 0 37536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input149_A
timestamp 1644511149
transform -1 0 37536 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input150_A
timestamp 1644511149
transform -1 0 37536 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input151_A
timestamp 1644511149
transform -1 0 37536 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input152_A
timestamp 1644511149
transform -1 0 37444 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input153_A
timestamp 1644511149
transform -1 0 38180 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input154_A
timestamp 1644511149
transform -1 0 37536 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input155_A
timestamp 1644511149
transform -1 0 36800 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input156_A
timestamp 1644511149
transform -1 0 36800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input157_A
timestamp 1644511149
transform -1 0 36248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input158_A
timestamp 1644511149
transform -1 0 37444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input159_A
timestamp 1644511149
transform -1 0 38180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input160_A
timestamp 1644511149
transform -1 0 34868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input161_A
timestamp 1644511149
transform -1 0 37536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input162_A
timestamp 1644511149
transform -1 0 36892 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input163_A
timestamp 1644511149
transform -1 0 37536 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1644511149
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1644511149
transform -1 0 27048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output185_A
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output198_A
timestamp 1644511149
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output199_A
timestamp 1644511149
transform 1 0 16100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output204_A
timestamp 1644511149
transform -1 0 13432 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output209_A
timestamp 1644511149
transform -1 0 18768 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1644511149
transform 1 0 19872 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output223_A
timestamp 1644511149
transform 1 0 30820 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output224_A
timestamp 1644511149
transform 1 0 3036 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output225_A
timestamp 1644511149
transform 1 0 31924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1644511149
transform 1 0 32936 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1644511149
transform 1 0 34040 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output228_A
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output229_A
timestamp 1644511149
transform 1 0 35236 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1644511149
transform -1 0 36248 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1644511149
transform -1 0 34868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1644511149
transform -1 0 36892 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output233_A
timestamp 1644511149
transform -1 0 4508 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output242_A
timestamp 1644511149
transform -1 0 12972 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output243_A
timestamp 1644511149
transform 1 0 13892 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output244_A
timestamp 1644511149
transform 1 0 14536 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output245_A
timestamp 1644511149
transform 1 0 15916 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output246_A
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output247_A
timestamp 1644511149
transform -1 0 18216 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output248_A
timestamp 1644511149
transform 1 0 20424 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output249_A
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output252_A
timestamp 1644511149
transform 1 0 21896 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output253_A
timestamp 1644511149
transform 1 0 22816 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output254_A
timestamp 1644511149
transform -1 0 25024 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output255_A
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output256_A
timestamp 1644511149
transform -1 0 27140 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output261_A
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output262_A
timestamp 1644511149
transform -1 0 3772 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output263_A
timestamp 1644511149
transform -1 0 33856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output264_A
timestamp 1644511149
transform 1 0 33856 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output265_A
timestamp 1644511149
transform -1 0 34868 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output266_A
timestamp 1644511149
transform 1 0 35236 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output267_A
timestamp 1644511149
transform 1 0 35236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output268_A
timestamp 1644511149
transform 1 0 37444 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output270_A
timestamp 1644511149
transform -1 0 36340 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output271_A
timestamp 1644511149
transform -1 0 5060 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output272_A
timestamp 1644511149
transform -1 0 5612 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output273_A
timestamp 1644511149
transform -1 0 7452 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output274_A
timestamp 1644511149
transform -1 0 8004 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output275_A
timestamp 1644511149
transform -1 0 9292 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output276_A
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output277_A
timestamp 1644511149
transform -1 0 12236 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1644511149
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1644511149
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1644511149
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1644511149
transform 1 0 15640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1644511149
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1644511149
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_263
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_271
timestamp 1644511149
transform 1 0 26036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_348
timestamp 1644511149
transform 1 0 33120 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_42
timestamp 1644511149
transform 1 0 4968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_48
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1644511149
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1644511149
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 1644511149
transform 1 0 15088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1644511149
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_173
timestamp 1644511149
transform 1 0 17020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1644511149
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_207
timestamp 1644511149
transform 1 0 20148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_252
timestamp 1644511149
transform 1 0 24288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1644511149
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_313
timestamp 1644511149
transform 1 0 29900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_319
timestamp 1644511149
transform 1 0 30452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1644511149
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_351
timestamp 1644511149
transform 1 0 33396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_359
timestamp 1644511149
transform 1 0 34132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1644511149
transform 1 0 34684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1644511149
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1644511149
transform 1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_115
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_150
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1644511149
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_267
timestamp 1644511149
transform 1 0 25668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1644511149
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1644511149
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1644511149
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_324
timestamp 1644511149
transform 1 0 30912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1644511149
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_340
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_348
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_373
timestamp 1644511149
transform 1 0 35420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_385
timestamp 1644511149
transform 1 0 36524 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_61
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1644511149
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1644511149
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1644511149
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_203
timestamp 1644511149
transform 1 0 19780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_236
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_241
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_245
timestamp 1644511149
transform 1 0 23644 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_250
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_284
timestamp 1644511149
transform 1 0 27232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_291
timestamp 1644511149
transform 1 0 27876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1644511149
transform 1 0 28980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_313
timestamp 1644511149
transform 1 0 29900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_321
timestamp 1644511149
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_341
timestamp 1644511149
transform 1 0 32476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_348
timestamp 1644511149
transform 1 0 33120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_356
timestamp 1644511149
transform 1 0 33856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_375
timestamp 1644511149
transform 1 0 35604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_397
timestamp 1644511149
transform 1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 1644511149
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_37
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_45
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1644511149
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_68
timestamp 1644511149
transform 1 0 7360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1644511149
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_100
timestamp 1644511149
transform 1 0 10304 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_108
timestamp 1644511149
transform 1 0 11040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1644511149
transform 1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1644511149
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_123
timestamp 1644511149
transform 1 0 12420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1644511149
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_144
timestamp 1644511149
transform 1 0 14352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1644511149
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1644511149
transform 1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_164
timestamp 1644511149
transform 1 0 16192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 1644511149
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1644511149
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1644511149
transform 1 0 21160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_225
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_238
timestamp 1644511149
transform 1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1644511149
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_264
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1644511149
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1644511149
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_311
timestamp 1644511149
transform 1 0 29716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_317
timestamp 1644511149
transform 1 0 30268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_329
timestamp 1644511149
transform 1 0 31372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_341
timestamp 1644511149
transform 1 0 32476 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_353
timestamp 1644511149
transform 1 0 33580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_373
timestamp 1644511149
transform 1 0 35420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_379
timestamp 1644511149
transform 1 0 35972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_384
timestamp 1644511149
transform 1 0 36432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1644511149
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_5
timestamp 1644511149
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1644511149
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_59
timestamp 1644511149
transform 1 0 6532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1644511149
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_68
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_76
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1644511149
transform 1 0 8648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1644511149
transform 1 0 10304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1644511149
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1644511149
transform 1 0 12420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 1644511149
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1644511149
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_141
timestamp 1644511149
transform 1 0 14076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_147
timestamp 1644511149
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_150
timestamp 1644511149
transform 1 0 14904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1644511149
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_171
timestamp 1644511149
transform 1 0 16836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1644511149
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_192
timestamp 1644511149
transform 1 0 18768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_201
timestamp 1644511149
transform 1 0 19596 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_211
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_215
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1644511149
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_227
timestamp 1644511149
transform 1 0 21988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_239
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_247
timestamp 1644511149
transform 1 0 23828 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_253
timestamp 1644511149
transform 1 0 24380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_269
timestamp 1644511149
transform 1 0 25852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1644511149
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_285
timestamp 1644511149
transform 1 0 27324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_288
timestamp 1644511149
transform 1 0 27600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_294
timestamp 1644511149
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1644511149
transform 1 0 28520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1644511149
transform 1 0 28796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_308
timestamp 1644511149
transform 1 0 29440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1644511149
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_321
timestamp 1644511149
transform 1 0 30636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1644511149
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_340
timestamp 1644511149
transform 1 0 32384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_346
timestamp 1644511149
transform 1 0 32936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_350
timestamp 1644511149
transform 1 0 33304 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_359
timestamp 1644511149
transform 1 0 34132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_369
timestamp 1644511149
transform 1 0 35052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_377
timestamp 1644511149
transform 1 0 35788 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_383
timestamp 1644511149
transform 1 0 36340 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1644511149
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_5
timestamp 1644511149
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1644511149
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1644511149
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1644511149
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1644511149
transform 1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_62
timestamp 1644511149
transform 1 0 6808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_73
timestamp 1644511149
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1644511149
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_91 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1644511149
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1644511149
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_149
timestamp 1644511149
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1644511149
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_211
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_220
timestamp 1644511149
transform 1 0 21344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_226
timestamp 1644511149
transform 1 0 21896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1644511149
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_256
timestamp 1644511149
transform 1 0 24656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_260
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_263
timestamp 1644511149
transform 1 0 25300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1644511149
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1644511149
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_294
timestamp 1644511149
transform 1 0 28152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_317
timestamp 1644511149
transform 1 0 30268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_329
timestamp 1644511149
transform 1 0 31372 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_337
timestamp 1644511149
transform 1 0 32108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_343
timestamp 1644511149
transform 1 0 32660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_346
timestamp 1644511149
transform 1 0 32936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1644511149
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1644511149
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_368
timestamp 1644511149
transform 1 0 34960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_372
timestamp 1644511149
transform 1 0 35328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_376
timestamp 1644511149
transform 1 0 35696 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_382
timestamp 1644511149
transform 1 0 36248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_387
timestamp 1644511149
transform 1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1644511149
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_5
timestamp 1644511149
transform 1 0 1564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_17
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1644511149
transform 1 0 3220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1644511149
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1644511149
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1644511149
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1644511149
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1644511149
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_180
timestamp 1644511149
transform 1 0 17664 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_192
timestamp 1644511149
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_204
timestamp 1644511149
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1644511149
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_311
timestamp 1644511149
transform 1 0 29716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1644511149
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_326
timestamp 1644511149
transform 1 0 31096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1644511149
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_339
timestamp 1644511149
transform 1 0 32292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_347
timestamp 1644511149
transform 1 0 33028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_355
timestamp 1644511149
transform 1 0 33764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_367
timestamp 1644511149
transform 1 0 34868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_374
timestamp 1644511149
transform 1 0 35512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_381
timestamp 1644511149
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1644511149
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_401
timestamp 1644511149
transform 1 0 37996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_46
timestamp 1644511149
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1644511149
transform 1 0 6440 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1644511149
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_67
timestamp 1644511149
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_151
timestamp 1644511149
transform 1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 1644511149
transform 1 0 16192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_174
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1644511149
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1644511149
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1644511149
transform 1 0 19596 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1644511149
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_214
timestamp 1644511149
transform 1 0 20792 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_217
timestamp 1644511149
transform 1 0 21068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_229
timestamp 1644511149
transform 1 0 22172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_241
timestamp 1644511149
transform 1 0 23276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1644511149
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_261
timestamp 1644511149
transform 1 0 25116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_273
timestamp 1644511149
transform 1 0 26220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_285
timestamp 1644511149
transform 1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_291
timestamp 1644511149
transform 1 0 27876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_297
timestamp 1644511149
transform 1 0 28428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1644511149
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_314
timestamp 1644511149
transform 1 0 29992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_322
timestamp 1644511149
transform 1 0 30728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_328
timestamp 1644511149
transform 1 0 31280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_338
timestamp 1644511149
transform 1 0 32200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_344
timestamp 1644511149
transform 1 0 32752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_350
timestamp 1644511149
transform 1 0 33304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_356
timestamp 1644511149
transform 1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_367
timestamp 1644511149
transform 1 0 34868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_379
timestamp 1644511149
transform 1 0 35972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_382
timestamp 1644511149
transform 1 0 36248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_388
timestamp 1644511149
transform 1 0 36800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1644511149
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1644511149
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1644511149
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_92
timestamp 1644511149
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1644511149
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_116
timestamp 1644511149
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_128
timestamp 1644511149
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_140
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_158
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_284
timestamp 1644511149
transform 1 0 27232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_290
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1644511149
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_301
timestamp 1644511149
transform 1 0 28796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_313
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_325
timestamp 1644511149
transform 1 0 31004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1644511149
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1644511149
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_365
timestamp 1644511149
transform 1 0 34684 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_376
timestamp 1644511149
transform 1 0 35696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_382
timestamp 1644511149
transform 1 0 36248 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1644511149
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_401
timestamp 1644511149
transform 1 0 37996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1644511149
transform 1 0 11868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_129
timestamp 1644511149
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1644511149
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_211
timestamp 1644511149
transform 1 0 20516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_223
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_235
timestamp 1644511149
transform 1 0 22724 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_273
timestamp 1644511149
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_285
timestamp 1644511149
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_297
timestamp 1644511149
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1644511149
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_317
timestamp 1644511149
transform 1 0 30268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1644511149
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_342
timestamp 1644511149
transform 1 0 32568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_354
timestamp 1644511149
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1644511149
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_370
timestamp 1644511149
transform 1 0 35144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_376
timestamp 1644511149
transform 1 0 35696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_386
timestamp 1644511149
transform 1 0 36616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_394
timestamp 1644511149
transform 1 0 37352 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1644511149
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_22
timestamp 1644511149
transform 1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_35
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1644511149
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1644511149
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1644511149
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1644511149
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1644511149
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_97
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1644511149
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_119
timestamp 1644511149
transform 1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp 1644511149
transform 1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1644511149
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1644511149
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp 1644511149
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1644511149
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_254
timestamp 1644511149
transform 1 0 24472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_260
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_266
timestamp 1644511149
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1644511149
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_345
timestamp 1644511149
transform 1 0 32844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1644511149
transform 1 0 33672 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_366
timestamp 1644511149
transform 1 0 34776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_374
timestamp 1644511149
transform 1 0 35512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_377
timestamp 1644511149
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_383
timestamp 1644511149
transform 1 0 36340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_397
timestamp 1644511149
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1644511149
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_31
timestamp 1644511149
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_39
timestamp 1644511149
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1644511149
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1644511149
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_103
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1644511149
transform 1 0 11684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_127
timestamp 1644511149
transform 1 0 12788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1644511149
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1644511149
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_261
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_272
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_278
timestamp 1644511149
transform 1 0 26680 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_290
timestamp 1644511149
transform 1 0 27784 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1644511149
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_374
timestamp 1644511149
transform 1 0 35512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_381
timestamp 1644511149
transform 1 0 36156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_387
timestamp 1644511149
transform 1 0 36708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_393
timestamp 1644511149
transform 1 0 37260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_396
timestamp 1644511149
transform 1 0 37536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1644511149
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1644511149
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_146
timestamp 1644511149
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1644511149
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1644511149
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_177
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_201
timestamp 1644511149
transform 1 0 19596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1644511149
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1644511149
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_301
timestamp 1644511149
transform 1 0 28796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_306
timestamp 1644511149
transform 1 0 29256 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1644511149
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_49
timestamp 1644511149
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1644511149
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1644511149
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_157
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_175
timestamp 1644511149
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1644511149
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1644511149
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1644511149
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1644511149
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1644511149
transform 1 0 13524 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1644511149
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1644511149
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_179
timestamp 1644511149
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_191
timestamp 1644511149
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1644511149
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_289
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_292
timestamp 1644511149
transform 1 0 27968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_304
timestamp 1644511149
transform 1 0 29072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_316
timestamp 1644511149
transform 1 0 30176 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1644511149
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_381
timestamp 1644511149
transform 1 0 36156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1644511149
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_397
timestamp 1644511149
transform 1 0 37628 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1644511149
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1644511149
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1644511149
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_185
timestamp 1644511149
transform 1 0 18124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1644511149
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1644511149
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1644511149
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_283
timestamp 1644511149
transform 1 0 27140 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1644511149
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1644511149
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1644511149
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_29
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_41
timestamp 1644511149
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1644511149
transform 1 0 10028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1644511149
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_131
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_143
timestamp 1644511149
transform 1 0 14260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_155
timestamp 1644511149
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1644511149
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_202
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1644511149
transform 1 0 24748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1644511149
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_289
timestamp 1644511149
transform 1 0 27692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_299
timestamp 1644511149
transform 1 0 28612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_311
timestamp 1644511149
transform 1 0 29716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_315
timestamp 1644511149
transform 1 0 30084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_322
timestamp 1644511149
transform 1 0 30728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1644511149
transform 1 0 4508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_49
timestamp 1644511149
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_61
timestamp 1644511149
transform 1 0 6716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1644511149
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1644511149
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_100
timestamp 1644511149
transform 1 0 10304 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_112
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_124
timestamp 1644511149
transform 1 0 12512 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1644511149
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_216
timestamp 1644511149
transform 1 0 20976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_228
timestamp 1644511149
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_240
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_293
timestamp 1644511149
transform 1 0 28060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1644511149
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_331
timestamp 1644511149
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_343
timestamp 1644511149
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1644511149
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1644511149
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_85
timestamp 1644511149
transform 1 0 8924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_97
timestamp 1644511149
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1644511149
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_133
timestamp 1644511149
transform 1 0 13340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_145
timestamp 1644511149
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1644511149
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1644511149
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_204
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1644511149
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_247
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_259
timestamp 1644511149
transform 1 0 24932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1644511149
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_347
timestamp 1644511149
transform 1 0 33028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_354
timestamp 1644511149
transform 1 0 33672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_360
timestamp 1644511149
transform 1 0 34224 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_372
timestamp 1644511149
transform 1 0 35328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1644511149
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_399
timestamp 1644511149
transform 1 0 37812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1644511149
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_147
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_159
timestamp 1644511149
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_183
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_232
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_255
timestamp 1644511149
transform 1 0 24564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_267
timestamp 1644511149
transform 1 0 25668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_279
timestamp 1644511149
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_397
timestamp 1644511149
transform 1 0 37628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1644511149
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1644511149
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1644511149
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_177
timestamp 1644511149
transform 1 0 17388 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1644511149
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_255
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_263
timestamp 1644511149
transform 1 0 25300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1644511149
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_325
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_401
timestamp 1644511149
transform 1 0 37996 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1644511149
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_145
timestamp 1644511149
transform 1 0 14444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1644511149
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_229
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1644511149
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_255
timestamp 1644511149
transform 1 0 24564 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_267
timestamp 1644511149
transform 1 0 25668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_279
timestamp 1644511149
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_291
timestamp 1644511149
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1644511149
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_311
timestamp 1644511149
transform 1 0 29716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_323
timestamp 1644511149
transform 1 0 30820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_335
timestamp 1644511149
transform 1 0 31924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_347
timestamp 1644511149
transform 1 0 33028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1644511149
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_385
timestamp 1644511149
transform 1 0 36524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_72
timestamp 1644511149
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_84
timestamp 1644511149
transform 1 0 8832 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_96
timestamp 1644511149
transform 1 0 9936 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_177
timestamp 1644511149
transform 1 0 17388 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1644511149
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_239
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_242
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_248
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_260
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1644511149
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_291
timestamp 1644511149
transform 1 0 27876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_301
timestamp 1644511149
transform 1 0 28796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_311
timestamp 1644511149
transform 1 0 29716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_323
timestamp 1644511149
transform 1 0 30820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1644511149
transform 1 0 36064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_397
timestamp 1644511149
transform 1 0 37628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1644511149
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_35
timestamp 1644511149
transform 1 0 4324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_47
timestamp 1644511149
transform 1 0 5428 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_59
timestamp 1644511149
transform 1 0 6532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_71
timestamp 1644511149
transform 1 0 7636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1644511149
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1644511149
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_124
timestamp 1644511149
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1644511149
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1644511149
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1644511149
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_290
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1644511149
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_313
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_322
timestamp 1644511149
transform 1 0 30728 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_336
timestamp 1644511149
transform 1 0 32016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_342
timestamp 1644511149
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1644511149
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1644511149
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_368
timestamp 1644511149
transform 1 0 34960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_374
timestamp 1644511149
transform 1 0 35512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_382
timestamp 1644511149
transform 1 0 36248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_386
timestamp 1644511149
transform 1 0 36616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1644511149
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_398
timestamp 1644511149
transform 1 0 37720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1644511149
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_195
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_207
timestamp 1644511149
transform 1 0 20148 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_323
timestamp 1644511149
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_353
timestamp 1644511149
transform 1 0 33580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_366
timestamp 1644511149
transform 1 0 34776 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_378
timestamp 1644511149
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1644511149
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_401
timestamp 1644511149
transform 1 0 37996 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1644511149
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_67
timestamp 1644511149
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1644511149
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1644511149
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1644511149
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_183
timestamp 1644511149
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1644511149
transform 1 0 32292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1644511149
transform 1 0 33396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_397
timestamp 1644511149
transform 1 0 37628 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1644511149
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_65
timestamp 1644511149
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1644511149
transform 1 0 8004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_128
timestamp 1644511149
transform 1 0 12880 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_134
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_146
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_360
timestamp 1644511149
transform 1 0 34224 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_372
timestamp 1644511149
transform 1 0 35328 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 1644511149
transform 1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_34
timestamp 1644511149
transform 1 0 4232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_46
timestamp 1644511149
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_58
timestamp 1644511149
transform 1 0 6440 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_70
timestamp 1644511149
transform 1 0 7544 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_89
timestamp 1644511149
transform 1 0 9292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_95
timestamp 1644511149
transform 1 0 9844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_107
timestamp 1644511149
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_119
timestamp 1644511149
transform 1 0 12052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1644511149
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_255
timestamp 1644511149
transform 1 0 24564 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_267
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_279
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_291
timestamp 1644511149
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1644511149
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_397
timestamp 1644511149
transform 1 0 37628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_177
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_183
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_195
timestamp 1644511149
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_207
timestamp 1644511149
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1644511149
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_206
timestamp 1644511149
transform 1 0 20056 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_230
timestamp 1644511149
transform 1 0 22264 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_269
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_367
timestamp 1644511149
transform 1 0 34868 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_379
timestamp 1644511149
transform 1 0 35972 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_391
timestamp 1644511149
transform 1 0 37076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1644511149
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_140
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_152
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_312
timestamp 1644511149
transform 1 0 29808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_353
timestamp 1644511149
transform 1 0 33580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_363
timestamp 1644511149
transform 1 0 34500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_398
timestamp 1644511149
transform 1 0 37720 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1644511149
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_37
timestamp 1644511149
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_49
timestamp 1644511149
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1644511149
transform 1 0 6716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_69
timestamp 1644511149
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1644511149
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_100
timestamp 1644511149
transform 1 0 10304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_112
timestamp 1644511149
transform 1 0 11408 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1644511149
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_229
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_242
timestamp 1644511149
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_285
timestamp 1644511149
transform 1 0 27324 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1644511149
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_319
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_326
timestamp 1644511149
transform 1 0 31096 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_332
timestamp 1644511149
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_344
timestamp 1644511149
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1644511149
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_66
timestamp 1644511149
transform 1 0 7176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_78
timestamp 1644511149
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_90
timestamp 1644511149
transform 1 0 9384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1644511149
transform 1 0 11684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1644511149
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_299
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_323
timestamp 1644511149
transform 1 0 30820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_396
timestamp 1644511149
transform 1 0 37536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1644511149
transform 1 0 38180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_63
timestamp 1644511149
transform 1 0 6900 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_69
timestamp 1644511149
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1644511149
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1644511149
transform 1 0 12420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1644511149
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_400
timestamp 1644511149
transform 1 0 37904 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1644511149
transform 1 0 38456 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1644511149
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_26
timestamp 1644511149
transform 1 0 3496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1644511149
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1644511149
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_246
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1644511149
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp 1644511149
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1644511149
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_60
timestamp 1644511149
transform 1 0 6624 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_72
timestamp 1644511149
transform 1 0 7728 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_219
timestamp 1644511149
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_231
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1644511149
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_316
timestamp 1644511149
transform 1 0 30176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_329
timestamp 1644511149
transform 1 0 31372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_341
timestamp 1644511149
transform 1 0 32476 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1644511149
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_393
timestamp 1644511149
transform 1 0 37260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_396
timestamp 1644511149
transform 1 0 37536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_230
timestamp 1644511149
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_345
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_358
timestamp 1644511149
transform 1 0 34040 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_366
timestamp 1644511149
transform 1 0 34776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_371
timestamp 1644511149
transform 1 0 35236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1644511149
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_401
timestamp 1644511149
transform 1 0 37996 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_173
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1644511149
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1644511149
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_215
timestamp 1644511149
transform 1 0 20884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_220
timestamp 1644511149
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1644511149
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_284
timestamp 1644511149
transform 1 0 27232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_290
timestamp 1644511149
transform 1 0 27784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1644511149
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_337
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_348
timestamp 1644511149
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_397
timestamp 1644511149
transform 1 0 37628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_192
timestamp 1644511149
transform 1 0 18768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_198
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1644511149
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_316
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_324
timestamp 1644511149
transform 1 0 30912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_339
timestamp 1644511149
transform 1 0 32292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_351
timestamp 1644511149
transform 1 0 33396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_363
timestamp 1644511149
transform 1 0 34500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_375
timestamp 1644511149
transform 1 0 35604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1644511149
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_402
timestamp 1644511149
transform 1 0 38088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1644511149
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_128
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_259
timestamp 1644511149
transform 1 0 24932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1644511149
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1644511149
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_329
timestamp 1644511149
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_341
timestamp 1644511149
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1644511149
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1644511149
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1644511149
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_73
timestamp 1644511149
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_77
timestamp 1644511149
transform 1 0 8188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_94
timestamp 1644511149
transform 1 0 9752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_102
timestamp 1644511149
transform 1 0 10488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_122
timestamp 1644511149
transform 1 0 12328 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_130
timestamp 1644511149
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_61
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1644511149
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1644511149
transform 1 0 9292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_129
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_157
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_169
timestamp 1644511149
transform 1 0 16652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1644511149
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1644511149
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_334
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_340
timestamp 1644511149
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_352
timestamp 1644511149
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_11
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1644511149
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_35
timestamp 1644511149
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1644511149
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_77
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_153
timestamp 1644511149
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1644511149
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_241
timestamp 1644511149
transform 1 0 23276 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_247
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_285
timestamp 1644511149
transform 1 0 27324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_309
timestamp 1644511149
transform 1 0 29532 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1644511149
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_399
timestamp 1644511149
transform 1 0 37812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_35
timestamp 1644511149
transform 1 0 4324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_47
timestamp 1644511149
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_59
timestamp 1644511149
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_71
timestamp 1644511149
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1644511149
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_357
timestamp 1644511149
transform 1 0 33948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_377
timestamp 1644511149
transform 1 0 35788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1644511149
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_35
timestamp 1644511149
transform 1 0 4324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_48
timestamp 1644511149
transform 1 0 5520 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1644511149
transform 1 0 6072 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1644511149
transform 1 0 7176 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1644511149
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_169
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_286
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_298
timestamp 1644511149
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1644511149
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_336
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_373
timestamp 1644511149
transform 1 0 35420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_397
timestamp 1644511149
transform 1 0 37628 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1644511149
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_269
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_299
timestamp 1644511149
transform 1 0 28612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_341
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_353
timestamp 1644511149
transform 1 0 33580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_365
timestamp 1644511149
transform 1 0 34684 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_377
timestamp 1644511149
transform 1 0 35788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1644511149
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_57
timestamp 1644511149
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_181
timestamp 1644511149
transform 1 0 17756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_278
timestamp 1644511149
transform 1 0 26680 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1644511149
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_317
timestamp 1644511149
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_324
timestamp 1644511149
transform 1 0 30912 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_336
timestamp 1644511149
transform 1 0 32016 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_348
timestamp 1644511149
transform 1 0 33120 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_98
timestamp 1644511149
transform 1 0 10120 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1644511149
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_117
timestamp 1644511149
transform 1 0 11868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1644511149
transform 1 0 12420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_135
timestamp 1644511149
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_147
timestamp 1644511149
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1644511149
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_239
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_245
timestamp 1644511149
transform 1 0 23644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_257
timestamp 1644511149
transform 1 0 24748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_269
timestamp 1644511149
transform 1 0 25852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1644511149
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_93
timestamp 1644511149
transform 1 0 9660 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_99
timestamp 1644511149
transform 1 0 10212 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_107
timestamp 1644511149
transform 1 0 10948 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_112
timestamp 1644511149
transform 1 0 11408 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_124
timestamp 1644511149
transform 1 0 12512 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_266
timestamp 1644511149
transform 1 0 25576 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_278
timestamp 1644511149
transform 1 0 26680 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_290
timestamp 1644511149
transform 1 0 27784 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1644511149
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_344
timestamp 1644511149
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_393
timestamp 1644511149
transform 1 0 37260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_396
timestamp 1644511149
transform 1 0 37536 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_13
timestamp 1644511149
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_25
timestamp 1644511149
transform 1 0 3404 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_33
timestamp 1644511149
transform 1 0 4140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_41
timestamp 1644511149
transform 1 0 4876 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1644511149
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_64
timestamp 1644511149
transform 1 0 6992 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_76
timestamp 1644511149
transform 1 0 8096 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_88
timestamp 1644511149
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_100
timestamp 1644511149
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_118
timestamp 1644511149
transform 1 0 11960 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_124
timestamp 1644511149
transform 1 0 12512 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_132
timestamp 1644511149
transform 1 0 13248 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_150
timestamp 1644511149
transform 1 0 14904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_154
timestamp 1644511149
transform 1 0 15272 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_158
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_179
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_185
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1644511149
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1644511149
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_236
timestamp 1644511149
transform 1 0 22816 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_248
timestamp 1644511149
transform 1 0 23920 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_260
timestamp 1644511149
transform 1 0 25024 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1644511149
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_345
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_357
timestamp 1644511149
transform 1 0 33948 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_369
timestamp 1644511149
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_381
timestamp 1644511149
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1644511149
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_31
timestamp 1644511149
transform 1 0 3956 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_39
timestamp 1644511149
transform 1 0 4692 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_43
timestamp 1644511149
transform 1 0 5060 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_49
timestamp 1644511149
transform 1 0 5612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_61
timestamp 1644511149
transform 1 0 6716 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_73
timestamp 1644511149
transform 1 0 7820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1644511149
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1644511149
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_255
timestamp 1644511149
transform 1 0 24564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_267
timestamp 1644511149
transform 1 0 25668 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_275
timestamp 1644511149
transform 1 0 26404 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_291
timestamp 1644511149
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1644511149
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_341
timestamp 1644511149
transform 1 0 32476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_348
timestamp 1644511149
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_369
timestamp 1644511149
transform 1 0 35052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1644511149
transform 1 0 35328 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1644511149
transform 1 0 36432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_396
timestamp 1644511149
transform 1 0 37536 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_404
timestamp 1644511149
transform 1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_368
timestamp 1644511149
transform 1 0 34960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_396
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1644511149
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_268
timestamp 1644511149
transform 1 0 25760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_285
timestamp 1644511149
transform 1 0 27324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_288
timestamp 1644511149
transform 1 0 27600 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_297
timestamp 1644511149
transform 1 0 28428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1644511149
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_64
timestamp 1644511149
transform 1 0 6992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1644511149
transform 1 0 7544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1644511149
transform 1 0 8648 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1644511149
transform 1 0 9752 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1644511149
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_133
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1644511149
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1644511149
transform 1 0 25392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_346
timestamp 1644511149
transform 1 0 32936 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_370
timestamp 1644511149
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1644511149
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1644511149
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_397
timestamp 1644511149
transform 1 0 37628 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1644511149
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_201
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_207
timestamp 1644511149
transform 1 0 20148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_219
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_231
timestamp 1644511149
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_293
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1644511149
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1644511149
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_383
timestamp 1644511149
transform 1 0 36340 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_97
timestamp 1644511149
transform 1 0 10028 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp 1644511149
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1644511149
transform 1 0 12420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_135
timestamp 1644511149
transform 1 0 13524 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_147
timestamp 1644511149
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1644511149
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_187
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_194
timestamp 1644511149
transform 1 0 18952 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_206
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1644511149
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_320
timestamp 1644511149
transform 1 0 30544 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_369
timestamp 1644511149
transform 1 0 35052 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_379
timestamp 1644511149
transform 1 0 35972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_382
timestamp 1644511149
transform 1 0 36248 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1644511149
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_395
timestamp 1644511149
transform 1 0 37444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1644511149
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_106
timestamp 1644511149
transform 1 0 10856 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_112
timestamp 1644511149
transform 1 0 11408 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_124
timestamp 1644511149
transform 1 0 12512 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_163
timestamp 1644511149
transform 1 0 16100 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_171
timestamp 1644511149
transform 1 0 16836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_175
timestamp 1644511149
transform 1 0 17204 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_183
timestamp 1644511149
transform 1 0 17940 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1644511149
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1644511149
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_241
timestamp 1644511149
transform 1 0 23276 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 1644511149
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_327
timestamp 1644511149
transform 1 0 31188 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_355
timestamp 1644511149
transform 1 0 33764 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_358
timestamp 1644511149
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_367
timestamp 1644511149
transform 1 0 34868 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_373
timestamp 1644511149
transform 1 0 35420 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_379
timestamp 1644511149
transform 1 0 35972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_386
timestamp 1644511149
transform 1 0 36616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_394
timestamp 1644511149
transform 1 0 37352 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_402
timestamp 1644511149
transform 1 0 38088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1644511149
transform 1 0 38456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_17
timestamp 1644511149
transform 1 0 2668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_23
timestamp 1644511149
transform 1 0 3220 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_29
timestamp 1644511149
transform 1 0 3772 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_35
timestamp 1644511149
transform 1 0 4324 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1644511149
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_59
timestamp 1644511149
transform 1 0 6532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_71
timestamp 1644511149
transform 1 0 7636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_83
timestamp 1644511149
transform 1 0 8740 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_89
timestamp 1644511149
transform 1 0 9292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_95
timestamp 1644511149
transform 1 0 9844 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_103
timestamp 1644511149
transform 1 0 10580 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_106
timestamp 1644511149
transform 1 0 10856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_115
timestamp 1644511149
transform 1 0 11684 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_121
timestamp 1644511149
transform 1 0 12236 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_129
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_141
timestamp 1644511149
transform 1 0 14076 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_145
timestamp 1644511149
transform 1 0 14444 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_148
timestamp 1644511149
transform 1 0 14720 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_154
timestamp 1644511149
transform 1 0 15272 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_160
timestamp 1644511149
transform 1 0 15824 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_173
timestamp 1644511149
transform 1 0 17020 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_177
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1644511149
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 1644511149
transform 1 0 19504 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_206
timestamp 1644511149
transform 1 0 20056 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_212
timestamp 1644511149
transform 1 0 20608 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_229
timestamp 1644511149
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_232
timestamp 1644511149
transform 1 0 22448 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_242
timestamp 1644511149
transform 1 0 23368 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_252
timestamp 1644511149
transform 1 0 24288 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_345
timestamp 1644511149
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_348
timestamp 1644511149
transform 1 0 33120 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_356
timestamp 1644511149
transform 1 0 33856 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_364
timestamp 1644511149
transform 1 0 34592 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1644511149
transform 1 0 34868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_380
timestamp 1644511149
transform 1 0 36064 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_395
timestamp 1644511149
transform 1 0 37444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1644511149
transform 1 0 38180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_13
timestamp 1644511149
transform 1 0 2300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1644511149
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_31
timestamp 1644511149
transform 1 0 3956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_37
timestamp 1644511149
transform 1 0 4508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_43
timestamp 1644511149
transform 1 0 5060 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_49
timestamp 1644511149
transform 1 0 5612 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_57
timestamp 1644511149
transform 1 0 6348 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_63
timestamp 1644511149
transform 1 0 6900 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_69
timestamp 1644511149
transform 1 0 7452 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_75
timestamp 1644511149
transform 1 0 8004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_87
timestamp 1644511149
transform 1 0 9108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_104
timestamp 1644511149
transform 1 0 10672 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_110
timestamp 1644511149
transform 1 0 11224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_116
timestamp 1644511149
transform 1 0 11776 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_122
timestamp 1644511149
transform 1 0 12328 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1644511149
transform 1 0 12880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_134
timestamp 1644511149
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_147
timestamp 1644511149
transform 1 0 14628 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_151
timestamp 1644511149
transform 1 0 14996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_155
timestamp 1644511149
transform 1 0 15364 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_162
timestamp 1644511149
transform 1 0 16008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_168
timestamp 1644511149
transform 1 0 16560 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1644511149
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_180
timestamp 1644511149
transform 1 0 17664 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_186
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_199
timestamp 1644511149
transform 1 0 19412 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_207
timestamp 1644511149
transform 1 0 20148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_213
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_219
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_235
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1644511149
transform 1 0 27600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_300
timestamp 1644511149
transform 1 0 28704 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_322
timestamp 1644511149
transform 1 0 30728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_331
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_337
timestamp 1644511149
transform 1 0 32108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_348
timestamp 1644511149
transform 1 0 33120 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_354
timestamp 1644511149
transform 1 0 33672 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_367
timestamp 1644511149
transform 1 0 34868 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_375
timestamp 1644511149
transform 1 0 35604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_395
timestamp 1644511149
transform 1 0 37444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_13
timestamp 1644511149
transform 1 0 2300 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_20
timestamp 1644511149
transform 1 0 2944 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_33
timestamp 1644511149
transform 1 0 4140 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_45
timestamp 1644511149
transform 1 0 5244 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_49
timestamp 1644511149
transform 1 0 5612 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1644511149
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_61
timestamp 1644511149
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_67
timestamp 1644511149
transform 1 0 7268 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_77
timestamp 1644511149
transform 1 0 8188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_84
timestamp 1644511149
transform 1 0 8832 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_92
timestamp 1644511149
transform 1 0 9568 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_97
timestamp 1644511149
transform 1 0 10028 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1644511149
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_116
timestamp 1644511149
transform 1 0 11776 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_120
timestamp 1644511149
transform 1 0 12144 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_124
timestamp 1644511149
transform 1 0 12512 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_130
timestamp 1644511149
transform 1 0 13064 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_136
timestamp 1644511149
transform 1 0 13616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_145
timestamp 1644511149
transform 1 0 14444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_152
timestamp 1644511149
transform 1 0 15088 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_156
timestamp 1644511149
transform 1 0 15456 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_172
timestamp 1644511149
transform 1 0 16928 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_179
timestamp 1644511149
transform 1 0 17572 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_185
timestamp 1644511149
transform 1 0 18124 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_196
timestamp 1644511149
transform 1 0 19136 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_203
timestamp 1644511149
transform 1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_209
timestamp 1644511149
transform 1 0 20332 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1644511149
transform 1 0 22632 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_242
timestamp 1644511149
transform 1 0 23368 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1644511149
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_254
timestamp 1644511149
transform 1 0 24472 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_266
timestamp 1644511149
transform 1 0 25576 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_272
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_283
timestamp 1644511149
transform 1 0 27140 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_297
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_303
timestamp 1644511149
transform 1 0 28980 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_314
timestamp 1644511149
transform 1 0 29992 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_322
timestamp 1644511149
transform 1 0 30728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_326
timestamp 1644511149
transform 1 0 31096 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_341
timestamp 1644511149
transform 1 0 32476 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_346
timestamp 1644511149
transform 1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_354
timestamp 1644511149
transform 1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1644511149
transform 1 0 34408 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_366
timestamp 1644511149
transform 1 0 34776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_371
timestamp 1644511149
transform 1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_379
timestamp 1644511149
transform 1 0 35972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_383
timestamp 1644511149
transform 1 0 36340 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1644511149
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_395
timestamp 1644511149
transform 1 0 37444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_35
timestamp 1644511149
transform 1 0 4324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_39
timestamp 1644511149
transform 1 0 4692 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_42
timestamp 1644511149
transform 1 0 4968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_49
timestamp 1644511149
transform 1 0 5612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_58
timestamp 1644511149
transform 1 0 6440 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_70
timestamp 1644511149
transform 1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_89
timestamp 1644511149
transform 1 0 9292 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_95
timestamp 1644511149
transform 1 0 9844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_100
timestamp 1644511149
transform 1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_108
timestamp 1644511149
transform 1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_116
timestamp 1644511149
transform 1 0 11776 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_122
timestamp 1644511149
transform 1 0 12328 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_127
timestamp 1644511149
transform 1 0 12788 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_145
timestamp 1644511149
transform 1 0 14444 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1644511149
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_159
timestamp 1644511149
transform 1 0 15732 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_164
timestamp 1644511149
transform 1 0 16192 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_173
timestamp 1644511149
transform 1 0 17020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_179
timestamp 1644511149
transform 1 0 17572 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_184
timestamp 1644511149
transform 1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1644511149
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_201
timestamp 1644511149
transform 1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_208
timestamp 1644511149
transform 1 0 20240 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_215
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1644511149
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1644511149
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_264
timestamp 1644511149
transform 1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_268
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_271
timestamp 1644511149
transform 1 0 26036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_278
timestamp 1644511149
transform 1 0 26680 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_285
timestamp 1644511149
transform 1 0 27324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_291
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1644511149
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_311
timestamp 1644511149
transform 1 0 29716 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_315
timestamp 1644511149
transform 1 0 30084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_320
timestamp 1644511149
transform 1 0 30544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_328
timestamp 1644511149
transform 1 0 31280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_336
timestamp 1644511149
transform 1 0 32016 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_344
timestamp 1644511149
transform 1 0 32752 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_354
timestamp 1644511149
transform 1 0 33672 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_369
timestamp 1644511149
transform 1 0 35052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_375
timestamp 1644511149
transform 1 0 35604 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_11
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_35
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_61
timestamp 1644511149
transform 1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_77
timestamp 1644511149
transform 1 0 8188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_85
timestamp 1644511149
transform 1 0 8924 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_103
timestamp 1644511149
transform 1 0 10580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_115
timestamp 1644511149
transform 1 0 11684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_123
timestamp 1644511149
transform 1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1644511149
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_139
timestamp 1644511149
transform 1 0 13892 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_147
timestamp 1644511149
transform 1 0 14628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_153
timestamp 1644511149
transform 1 0 15180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_157
timestamp 1644511149
transform 1 0 15548 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1644511149
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_177
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1644511149
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_211
timestamp 1644511149
transform 1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1644511149
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_253
timestamp 1644511149
transform 1 0 24380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_269
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_285
timestamp 1644511149
transform 1 0 27324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1644511149
transform 1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_324
timestamp 1644511149
transform 1 0 30912 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_341
timestamp 1644511149
transform 1 0 32476 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_347
timestamp 1644511149
transform 1 0 33028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_352
timestamp 1644511149
transform 1 0 33488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_364
timestamp 1644511149
transform 1 0 34592 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_370
timestamp 1644511149
transform 1 0 35144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_375
timestamp 1644511149
transform 1 0 35604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_387
timestamp 1644511149
transform 1 0 36708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1644511149
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1644511149
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_13
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1644511149
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_52
timestamp 1644511149
transform 1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_67
timestamp 1644511149
transform 1 0 7268 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_75
timestamp 1644511149
transform 1 0 8004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_95
timestamp 1644511149
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_103
timestamp 1644511149
transform 1 0 10580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1644511149
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_123
timestamp 1644511149
transform 1 0 12420 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_149
timestamp 1644511149
transform 1 0 14812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_157
timestamp 1644511149
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_163
timestamp 1644511149
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1644511149
transform 1 0 17940 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_190
timestamp 1644511149
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_201
timestamp 1644511149
transform 1 0 19596 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_211
timestamp 1644511149
transform 1 0 20516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 1644511149
transform 1 0 21252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1644511149
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_241
timestamp 1644511149
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1644511149
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_257
timestamp 1644511149
transform 1 0 24748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_263
timestamp 1644511149
transform 1 0 25300 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_268
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1644511149
transform 1 0 26496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_285
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1644511149
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1644511149
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_313
timestamp 1644511149
transform 1 0 29900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1644511149
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 1644511149
transform 1 0 34132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_369
timestamp 1644511149
transform 1 0 35052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1644511149
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1644511149
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_397
timestamp 1644511149
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _193_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _194_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _195_
timestamp 1644511149
transform 1 0 9200 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1644511149
transform -1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _197_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1644511149
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _199_
timestamp 1644511149
transform 1 0 12052 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1644511149
transform -1 0 12420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _201_
timestamp 1644511149
transform 1 0 14444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1644511149
transform -1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _203_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27876 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _204_
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _205_
timestamp 1644511149
transform -1 0 23828 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _206_
timestamp 1644511149
transform 1 0 25944 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _207_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _208_
timestamp 1644511149
transform 1 0 22356 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _209_
timestamp 1644511149
transform -1 0 23184 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _210_
timestamp 1644511149
transform -1 0 32016 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1644511149
transform -1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _212_
timestamp 1644511149
transform 1 0 20332 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1644511149
transform 1 0 19320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _214_
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1644511149
transform -1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _216_
timestamp 1644511149
transform 1 0 25668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _218_
timestamp 1644511149
transform -1 0 29900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _220_
timestamp 1644511149
transform -1 0 24472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1644511149
transform -1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _222_
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _223_
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _224_
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1644511149
transform -1 0 25944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _226_
timestamp 1644511149
transform 1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1644511149
transform -1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _228_
timestamp 1644511149
transform 1 0 6532 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1644511149
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _230_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _231_
timestamp 1644511149
transform -1 0 27692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1644511149
transform -1 0 28704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _233_
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1644511149
transform -1 0 29256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _235_
timestamp 1644511149
transform 1 0 27968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1644511149
transform -1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _237_
timestamp 1644511149
transform -1 0 32200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1644511149
transform -1 0 33120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _239_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1644511149
transform -1 0 33672 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _241_
timestamp 1644511149
transform 1 0 14260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1644511149
transform -1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _243_
timestamp 1644511149
transform 1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1644511149
transform -1 0 35696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _245_
timestamp 1644511149
transform 1 0 16652 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1644511149
transform -1 0 36156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _247_
timestamp 1644511149
transform 1 0 35604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _248_
timestamp 1644511149
transform 1 0 36984 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_4  _249_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1644511149
transform 1 0 2668 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _251_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 3312 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _253_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _254_
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1644511149
transform -1 0 3496 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1644511149
transform 1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _258_
timestamp 1644511149
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1644511149
transform 1 0 6164 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp 1644511149
transform 1 0 5888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _261_
timestamp 1644511149
transform 1 0 32200 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _263_
timestamp 1644511149
transform -1 0 30544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _265_
timestamp 1644511149
transform -1 0 31280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _266_
timestamp 1644511149
transform -1 0 31648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _267_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _268_
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _269_
timestamp 1644511149
transform -1 0 32752 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_4  _270_
timestamp 1644511149
transform -1 0 32844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1644511149
transform 1 0 12236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _272_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _273_
timestamp 1644511149
transform -1 0 33672 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _274_
timestamp 1644511149
transform -1 0 13248 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _275_
timestamp 1644511149
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _277_
timestamp 1644511149
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1644511149
transform -1 0 16560 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _279_
timestamp 1644511149
transform -1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _281_
timestamp 1644511149
transform -1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _283_
timestamp 1644511149
transform -1 0 36892 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _284_
timestamp 1644511149
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1644511149
transform -1 0 20240 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1644511149
transform -1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _288_
timestamp 1644511149
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _289_
timestamp 1644511149
transform 1 0 22172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _290_
timestamp 1644511149
transform -1 0 10764 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _291_
timestamp 1644511149
transform 1 0 23552 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _292_
timestamp 1644511149
transform -1 0 11684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _293_
timestamp 1644511149
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp 1644511149
transform -1 0 13156 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _295_
timestamp 1644511149
transform 1 0 24748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _296_
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1644511149
transform 1 0 27048 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1644511149
transform -1 0 27324 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1644511149
transform 1 0 28612 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _301_
timestamp 1644511149
transform 1 0 22816 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1644511149
transform -1 0 28244 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1644511149
transform 1 0 31280 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _305_
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _306_
timestamp 1644511149
transform 1 0 30452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1644511149
transform 1 0 33948 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _308_
timestamp 1644511149
transform -1 0 34224 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1644511149
transform -1 0 19780 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _310_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1644511149
transform -1 0 20976 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _312_
timestamp 1644511149
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1644511149
transform -1 0 22632 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1644511149
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1644511149
transform -1 0 23828 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _316_
timestamp 1644511149
transform -1 0 35788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_4  _317_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 2668 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _319_
timestamp 1644511149
transform -1 0 30728 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _320_
timestamp 1644511149
transform -1 0 26036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_4  _321_
timestamp 1644511149
transform -1 0 32568 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _323_
timestamp 1644511149
transform -1 0 18216 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform -1 0 19780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _325_
timestamp 1644511149
transform 1 0 23736 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1644511149
transform -1 0 27784 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _327_
timestamp 1644511149
transform -1 0 28796 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _328_
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _329_
timestamp 1644511149
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _330_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27324 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _331_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22264 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _332_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20240 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _333_
timestamp 1644511149
transform -1 0 12880 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _334_
timestamp 1644511149
transform -1 0 13156 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _335_
timestamp 1644511149
transform -1 0 7728 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _336_
timestamp 1644511149
transform -1 0 7176 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _337_
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _338_
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _339_
timestamp 1644511149
transform 1 0 19780 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1644511149
transform -1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _341_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32476 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _342_
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _343_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32016 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _344_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _345_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _346_
timestamp 1644511149
transform -1 0 32752 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _347_
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1644511149
transform -1 0 34960 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _349_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26128 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1644511149
transform 1 0 5612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _351_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3128 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _352_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _353_
timestamp 1644511149
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _354_
timestamp 1644511149
transform 1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _355_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1644511149
transform 1 0 5336 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _357_
timestamp 1644511149
transform -1 0 7912 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1644511149
transform -1 0 6716 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _359_
timestamp 1644511149
transform -1 0 29992 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _360_
timestamp 1644511149
transform 1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _361_
timestamp 1644511149
transform -1 0 30820 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _363_
timestamp 1644511149
transform -1 0 31648 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1644511149
transform 1 0 10396 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _365_
timestamp 1644511149
transform -1 0 33672 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _366_
timestamp 1644511149
transform -1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _367_
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _369_
timestamp 1644511149
transform -1 0 15640 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1644511149
transform 1 0 14168 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _371_
timestamp 1644511149
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _373_
timestamp 1644511149
transform -1 0 18032 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp 1644511149
transform 1 0 17296 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _375_
timestamp 1644511149
transform -1 0 37720 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _376_
timestamp 1644511149
transform 1 0 37260 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _377_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1644511149
transform -1 0 20884 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _379_
timestamp 1644511149
transform 1 0 10120 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1644511149
transform -1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _381_
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _382_
timestamp 1644511149
transform -1 0 13616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _383_
timestamp 1644511149
transform -1 0 13064 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1644511149
transform -1 0 15364 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _385_
timestamp 1644511149
transform -1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1644511149
transform -1 0 16008 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1644511149
transform -1 0 26496 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _389_
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _390_
timestamp 1644511149
transform -1 0 26680 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _391_
timestamp 1644511149
transform 1 0 27968 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1644511149
transform -1 0 29440 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _393_
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _394_
timestamp 1644511149
transform 1 0 31372 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _395_
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _396_
timestamp 1644511149
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _397_
timestamp 1644511149
transform 1 0 20516 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _398_
timestamp 1644511149
transform 1 0 33028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _399_
timestamp 1644511149
transform 1 0 25208 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _400_
timestamp 1644511149
transform 1 0 33948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _401_
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _402_
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _403_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34960 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _404_
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _405_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33948 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _406_
timestamp 1644511149
transform -1 0 30452 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _407_
timestamp 1644511149
transform 1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _408_
timestamp 1644511149
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _409_
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _410_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23552 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _411_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _412_
timestamp 1644511149
transform -1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _413_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _414_
timestamp 1644511149
transform -1 0 27324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _415_
timestamp 1644511149
transform -1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _416_
timestamp 1644511149
transform 1 0 25024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _417_
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _418_
timestamp 1644511149
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _419_
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _420_
timestamp 1644511149
transform -1 0 21252 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _421_
timestamp 1644511149
transform 1 0 20976 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _422_
timestamp 1644511149
transform -1 0 18124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _423_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _424_
timestamp 1644511149
transform -1 0 20056 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _425_
timestamp 1644511149
transform -1 0 17940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _426_
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _427_
timestamp 1644511149
transform -1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _428_
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _429_
timestamp 1644511149
transform -1 0 13432 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _430_
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _431_
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _432_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _433_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1644511149
transform -1 0 9752 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1644511149
transform 1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1644511149
transform -1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _437_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13064 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _438_
timestamp 1644511149
transform 1 0 8096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _439_
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _440_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _441_
timestamp 1644511149
transform -1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1644511149
transform -1 0 4232 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _443_
timestamp 1644511149
transform -1 0 3312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _444_
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _445_
timestamp 1644511149
transform -1 0 7268 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _446_
timestamp 1644511149
transform -1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _447_
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _448_
timestamp 1644511149
transform 1 0 7360 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _449_
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _450_
timestamp 1644511149
transform 1 0 6808 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _451_
timestamp 1644511149
transform 1 0 6348 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _452_
timestamp 1644511149
transform 1 0 6716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _453_
timestamp 1644511149
transform 1 0 4416 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _454_
timestamp 1644511149
transform 1 0 5244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _455_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _456_
timestamp 1644511149
transform -1 0 5428 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _457_
timestamp 1644511149
transform 1 0 4784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _458_
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _459_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _460_
timestamp 1644511149
transform -1 0 6992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _461_
timestamp 1644511149
transform 1 0 5244 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _462_
timestamp 1644511149
transform -1 0 11868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _463_
timestamp 1644511149
transform 1 0 10120 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _464_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _465_
timestamp 1644511149
transform -1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _466_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _467_
timestamp 1644511149
transform -1 0 17572 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _468_
timestamp 1644511149
transform -1 0 15640 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _469_
timestamp 1644511149
transform 1 0 14352 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _470_
timestamp 1644511149
transform -1 0 19596 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _471_
timestamp 1644511149
transform 1 0 18400 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _472_
timestamp 1644511149
transform -1 0 19412 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _473_
timestamp 1644511149
transform -1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _474_
timestamp 1644511149
transform -1 0 18492 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _475_
timestamp 1644511149
transform -1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _476_
timestamp 1644511149
transform -1 0 22816 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _477_
timestamp 1644511149
transform -1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _478_
timestamp 1644511149
transform -1 0 27416 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _479_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _480_
timestamp 1644511149
transform -1 0 31648 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _481_
timestamp 1644511149
transform -1 0 23828 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1644511149
transform 1 0 25760 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1644511149
transform 1 0 25760 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1644511149
transform 1 0 17296 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1644511149
transform 1 0 6900 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1644511149
transform -1 0 15548 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1644511149
transform 1 0 2024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1644511149
transform 1 0 2668 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1644511149
transform 1 0 6900 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1644511149
transform 1 0 4600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1644511149
transform 1 0 2300 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1644511149
transform 1 0 1840 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1644511149
transform 1 0 4416 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1644511149
transform 1 0 9384 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1644511149
transform 1 0 8648 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1644511149
transform 1 0 14076 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1644511149
transform -1 0 23736 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1644511149
transform 1 0 27140 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1644511149
transform 1 0 36156 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1644511149
transform 1 0 35972 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1644511149
transform -1 0 35788 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1644511149
transform -1 0 36800 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _510__280 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _511__281
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _512__282
timestamp 1644511149
transform 1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _513__283
timestamp 1644511149
transform 1 0 37904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514__284
timestamp 1644511149
transform 1 0 37904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515__285
timestamp 1644511149
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _516_
timestamp 1644511149
transform 1 0 2576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1644511149
transform -1 0 30084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _518_
timestamp 1644511149
transform -1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1644511149
transform -1 0 36800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _520_
timestamp 1644511149
transform -1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1644511149
transform -1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _522_
timestamp 1644511149
transform -1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _523_
timestamp 1644511149
transform -1 0 30268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _524_
timestamp 1644511149
transform -1 0 36524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _525_
timestamp 1644511149
transform -1 0 37996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _526_
timestamp 1644511149
transform -1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _527_
timestamp 1644511149
transform -1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _528_
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _529_
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _530_
timestamp 1644511149
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _531_
timestamp 1644511149
transform 1 0 36984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _532_
timestamp 1644511149
transform 1 0 37628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _533_
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _534_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _535_
timestamp 1644511149
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _536_
timestamp 1644511149
transform 1 0 36432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform -1 0 10488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform -1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform -1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform -1 0 28612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform -1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 33028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 33856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform -1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1644511149
transform -1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform -1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 37444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform -1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform -1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform -1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1644511149
transform -1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 30544 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1644511149
transform 1 0 32200 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 33304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform -1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform -1 0 35420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform -1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 35880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform -1 0 38180 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform -1 0 35512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 27600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform -1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform -1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1644511149
transform -1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform -1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1644511149
transform 1 0 29992 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform -1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1644511149
transform 1 0 32476 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform -1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform -1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform -1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform -1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1644511149
transform 1 0 9476 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform -1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform -1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform -1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 24472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1644511149
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1644511149
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 11868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 12788 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1644511149
transform 1 0 12788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1644511149
transform -1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1644511149
transform 1 0 17020 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input85
timestamp 1644511149
transform 1 0 18032 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1644511149
transform 1 0 20148 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input88
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1644511149
transform -1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1644511149
transform -1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input93
timestamp 1644511149
transform 1 0 25392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1644511149
transform -1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1644511149
transform 1 0 31372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1644511149
transform -1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1644511149
transform 1 0 2668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1644511149
transform -1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1644511149
transform -1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1644511149
transform -1 0 35052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1644511149
transform -1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1644511149
transform -1 0 36524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1644511149
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1644511149
transform -1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1644511149
transform -1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1644511149
transform -1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input111
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 1644511149
transform 1 0 7636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input113
timestamp 1644511149
transform 1 0 9292 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1644511149
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input115
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1644511149
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input123
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input124
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1644511149
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input129
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1644511149
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1644511149
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1644511149
transform -1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1644511149
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1644511149
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input136
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input137
timestamp 1644511149
transform 1 0 8648 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1644511149
transform -1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1644511149
transform -1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1644511149
transform -1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1644511149
transform -1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1644511149
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1644511149
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1644511149
transform -1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input147
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1644511149
transform 1 0 37904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1644511149
transform 1 0 37904 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1644511149
transform 1 0 37904 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1644511149
transform -1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input153
timestamp 1644511149
transform -1 0 38180 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1644511149
transform 1 0 36340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1644511149
transform -1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input157
timestamp 1644511149
transform -1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input158
timestamp 1644511149
transform -1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1644511149
transform -1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1644511149
transform 1 0 35880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1644511149
transform 1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input162
timestamp 1644511149
transform 1 0 37260 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1644511149
transform 1 0 37904 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 32752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 35236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 36064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 36432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 37076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform -1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform -1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform 1 0 31004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform 1 0 32016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform -1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform -1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform -1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform -1 0 21068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform -1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform -1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform -1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform -1 0 24104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1644511149
transform -1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1644511149
transform -1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1644511149
transform -1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1644511149
transform -1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1644511149
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1644511149
transform 1 0 10672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1644511149
transform -1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1644511149
transform -1 0 13892 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1644511149
transform 1 0 14260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1644511149
transform -1 0 16008 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1644511149
transform -1 0 16192 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1644511149
transform -1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1644511149
transform -1 0 18860 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1644511149
transform -1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1644511149
transform -1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1644511149
transform 1 0 24748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1644511149
transform 1 0 27876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1644511149
transform 1 0 3220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1644511149
transform 1 0 33120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1644511149
transform 1 0 34224 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1644511149
transform 1 0 35236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1644511149
transform 1 0 36340 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1644511149
transform 1 0 36432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1644511149
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1644511149
transform 1 0 37812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1644511149
transform -1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1644511149
transform -1 0 5060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1644511149
transform 1 0 7084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1644511149
transform -1 0 8188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1644511149
transform -1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1644511149
transform -1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1644511149
transform -1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1644511149
transform -1 0 11776 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1644511149
transform -1 0 12788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1644511149
transform 1 0 14996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1644511149
transform -1 0 15916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1644511149
transform -1 0 17020 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1644511149
transform -1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1644511149
transform -1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1644511149
transform -1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1644511149
transform -1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1644511149
transform -1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1644511149
transform 1 0 23000 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1644511149
transform -1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1644511149
transform 1 0 27692 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1644511149
transform -1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1644511149
transform -1 0 30728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1644511149
transform 1 0 31648 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1644511149
transform -1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1644511149
transform -1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1644511149
transform 1 0 34040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1644511149
transform 1 0 35604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1644511149
transform -1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1644511149
transform 1 0 37720 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1644511149
transform 1 0 37812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1644511149
transform 1 0 36984 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1644511149
transform -1 0 4324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1644511149
transform 1 0 5428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1644511149
transform -1 0 6440 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1644511149
transform -1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1644511149
transform -1 0 9292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1644511149
transform -1 0 10028 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1644511149
transform -1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1644511149
transform -1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1644511149
transform -1 0 35604 0 1 34816
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 9936 800 10056 6 clk
port 0 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 gpio0_input[0]
port 1 nsew signal tristate
rlabel metal2 s 32678 0 32734 800 6 gpio0_input[10]
port 2 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 gpio0_input[11]
port 3 nsew signal tristate
rlabel metal2 s 34334 0 34390 800 6 gpio0_input[12]
port 4 nsew signal tristate
rlabel metal2 s 35162 0 35218 800 6 gpio0_input[13]
port 5 nsew signal tristate
rlabel metal2 s 35990 0 36046 800 6 gpio0_input[14]
port 6 nsew signal tristate
rlabel metal2 s 36818 0 36874 800 6 gpio0_input[15]
port 7 nsew signal tristate
rlabel metal2 s 37646 0 37702 800 6 gpio0_input[16]
port 8 nsew signal tristate
rlabel metal2 s 38474 0 38530 800 6 gpio0_input[17]
port 9 nsew signal tristate
rlabel metal2 s 39302 0 39358 800 6 gpio0_input[18]
port 10 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 gpio0_input[1]
port 11 nsew signal tristate
rlabel metal2 s 26146 0 26202 800 6 gpio0_input[2]
port 12 nsew signal tristate
rlabel metal2 s 26882 0 26938 800 6 gpio0_input[3]
port 13 nsew signal tristate
rlabel metal2 s 27710 0 27766 800 6 gpio0_input[4]
port 14 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 gpio0_input[5]
port 15 nsew signal tristate
rlabel metal2 s 29366 0 29422 800 6 gpio0_input[6]
port 16 nsew signal tristate
rlabel metal2 s 30194 0 30250 800 6 gpio0_input[7]
port 17 nsew signal tristate
rlabel metal2 s 31022 0 31078 800 6 gpio0_input[8]
port 18 nsew signal tristate
rlabel metal2 s 31850 0 31906 800 6 gpio0_input[9]
port 19 nsew signal tristate
rlabel metal2 s 24766 0 24822 800 6 gpio0_oe[0]
port 20 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 gpio0_oe[10]
port 21 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 gpio0_oe[11]
port 22 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 gpio0_oe[12]
port 23 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 gpio0_oe[13]
port 24 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 gpio0_oe[14]
port 25 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 gpio0_oe[15]
port 26 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 gpio0_oe[16]
port 27 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 gpio0_oe[17]
port 28 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 gpio0_oe[18]
port 29 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 gpio0_oe[1]
port 30 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 gpio0_oe[2]
port 31 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 gpio0_oe[3]
port 32 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 gpio0_oe[4]
port 33 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 gpio0_oe[5]
port 34 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 gpio0_oe[6]
port 35 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 gpio0_oe[7]
port 36 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 gpio0_oe[8]
port 37 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 gpio0_oe[9]
port 38 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 gpio0_output[0]
port 39 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 gpio0_output[10]
port 40 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 gpio0_output[11]
port 41 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 gpio0_output[12]
port 42 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 gpio0_output[13]
port 43 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 gpio0_output[14]
port 44 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 gpio0_output[15]
port 45 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 gpio0_output[16]
port 46 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 gpio0_output[17]
port 47 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 gpio0_output[18]
port 48 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 gpio0_output[1]
port 49 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 gpio0_output[2]
port 50 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 gpio0_output[3]
port 51 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 gpio0_output[4]
port 52 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 gpio0_output[5]
port 53 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 gpio0_output[6]
port 54 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gpio0_output[7]
port 55 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 gpio0_output[8]
port 56 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 gpio0_output[9]
port 57 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 gpio1_input[0]
port 58 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 gpio1_input[10]
port 59 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 gpio1_input[11]
port 60 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 gpio1_input[12]
port 61 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 gpio1_input[13]
port 62 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 gpio1_input[14]
port 63 nsew signal tristate
rlabel metal2 s 21178 0 21234 800 6 gpio1_input[15]
port 64 nsew signal tristate
rlabel metal2 s 22006 0 22062 800 6 gpio1_input[16]
port 65 nsew signal tristate
rlabel metal2 s 22834 0 22890 800 6 gpio1_input[17]
port 66 nsew signal tristate
rlabel metal2 s 23662 0 23718 800 6 gpio1_input[18]
port 67 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 gpio1_input[1]
port 68 nsew signal tristate
rlabel metal2 s 10506 0 10562 800 6 gpio1_input[2]
port 69 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 gpio1_input[3]
port 70 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 gpio1_input[4]
port 71 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 gpio1_input[5]
port 72 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 gpio1_input[6]
port 73 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 gpio1_input[7]
port 74 nsew signal tristate
rlabel metal2 s 15382 0 15438 800 6 gpio1_input[8]
port 75 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 gpio1_input[9]
port 76 nsew signal tristate
rlabel metal2 s 9126 0 9182 800 6 gpio1_oe[0]
port 77 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 gpio1_oe[10]
port 78 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 gpio1_oe[11]
port 79 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 gpio1_oe[12]
port 80 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 gpio1_oe[13]
port 81 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 gpio1_oe[14]
port 82 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 gpio1_oe[15]
port 83 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 gpio1_oe[16]
port 84 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 gpio1_oe[17]
port 85 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 gpio1_oe[18]
port 86 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 gpio1_oe[1]
port 87 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 gpio1_oe[2]
port 88 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 gpio1_oe[3]
port 89 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 gpio1_oe[4]
port 90 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 gpio1_oe[5]
port 91 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 gpio1_oe[6]
port 92 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 gpio1_oe[7]
port 93 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 gpio1_oe[8]
port 94 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 gpio1_oe[9]
port 95 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 gpio1_output[0]
port 96 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 gpio1_output[10]
port 97 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 gpio1_output[11]
port 98 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 gpio1_output[12]
port 99 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 gpio1_output[13]
port 100 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 gpio1_output[14]
port 101 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 gpio1_output[15]
port 102 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 gpio1_output[16]
port 103 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 gpio1_output[17]
port 104 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 gpio1_output[18]
port 105 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 gpio1_output[1]
port 106 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 gpio1_output[2]
port 107 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 gpio1_output[3]
port 108 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 gpio1_output[4]
port 109 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 gpio1_output[5]
port 110 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 gpio1_output[6]
port 111 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 gpio1_output[7]
port 112 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 gpio1_output[8]
port 113 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 gpio1_output[9]
port 114 nsew signal input
rlabel metal2 s 110 39200 166 40000 6 io_in[0]
port 115 nsew signal input
rlabel metal2 s 10598 39200 10654 40000 6 io_in[10]
port 116 nsew signal input
rlabel metal2 s 11610 39200 11666 40000 6 io_in[11]
port 117 nsew signal input
rlabel metal2 s 12714 39200 12770 40000 6 io_in[12]
port 118 nsew signal input
rlabel metal2 s 13726 39200 13782 40000 6 io_in[13]
port 119 nsew signal input
rlabel metal2 s 14830 39200 14886 40000 6 io_in[14]
port 120 nsew signal input
rlabel metal2 s 15842 39200 15898 40000 6 io_in[15]
port 121 nsew signal input
rlabel metal2 s 16946 39200 17002 40000 6 io_in[16]
port 122 nsew signal input
rlabel metal2 s 17958 39200 18014 40000 6 io_in[17]
port 123 nsew signal input
rlabel metal2 s 19062 39200 19118 40000 6 io_in[18]
port 124 nsew signal input
rlabel metal2 s 20074 39200 20130 40000 6 io_in[19]
port 125 nsew signal input
rlabel metal2 s 1122 39200 1178 40000 6 io_in[1]
port 126 nsew signal input
rlabel metal2 s 21086 39200 21142 40000 6 io_in[20]
port 127 nsew signal input
rlabel metal2 s 22190 39200 22246 40000 6 io_in[21]
port 128 nsew signal input
rlabel metal2 s 23202 39200 23258 40000 6 io_in[22]
port 129 nsew signal input
rlabel metal2 s 24306 39200 24362 40000 6 io_in[23]
port 130 nsew signal input
rlabel metal2 s 25318 39200 25374 40000 6 io_in[24]
port 131 nsew signal input
rlabel metal2 s 26422 39200 26478 40000 6 io_in[25]
port 132 nsew signal input
rlabel metal2 s 27434 39200 27490 40000 6 io_in[26]
port 133 nsew signal input
rlabel metal2 s 28538 39200 28594 40000 6 io_in[27]
port 134 nsew signal input
rlabel metal2 s 29550 39200 29606 40000 6 io_in[28]
port 135 nsew signal input
rlabel metal2 s 30562 39200 30618 40000 6 io_in[29]
port 136 nsew signal input
rlabel metal2 s 2134 39200 2190 40000 6 io_in[2]
port 137 nsew signal input
rlabel metal2 s 31666 39200 31722 40000 6 io_in[30]
port 138 nsew signal input
rlabel metal2 s 32678 39200 32734 40000 6 io_in[31]
port 139 nsew signal input
rlabel metal2 s 33782 39200 33838 40000 6 io_in[32]
port 140 nsew signal input
rlabel metal2 s 34794 39200 34850 40000 6 io_in[33]
port 141 nsew signal input
rlabel metal2 s 35898 39200 35954 40000 6 io_in[34]
port 142 nsew signal input
rlabel metal2 s 36910 39200 36966 40000 6 io_in[35]
port 143 nsew signal input
rlabel metal2 s 38014 39200 38070 40000 6 io_in[36]
port 144 nsew signal input
rlabel metal2 s 39026 39200 39082 40000 6 io_in[37]
port 145 nsew signal input
rlabel metal2 s 3238 39200 3294 40000 6 io_in[3]
port 146 nsew signal input
rlabel metal2 s 4250 39200 4306 40000 6 io_in[4]
port 147 nsew signal input
rlabel metal2 s 5354 39200 5410 40000 6 io_in[5]
port 148 nsew signal input
rlabel metal2 s 6366 39200 6422 40000 6 io_in[6]
port 149 nsew signal input
rlabel metal2 s 7470 39200 7526 40000 6 io_in[7]
port 150 nsew signal input
rlabel metal2 s 8482 39200 8538 40000 6 io_in[8]
port 151 nsew signal input
rlabel metal2 s 9586 39200 9642 40000 6 io_in[9]
port 152 nsew signal input
rlabel metal2 s 386 39200 442 40000 6 io_oeb[0]
port 153 nsew signal tristate
rlabel metal2 s 10966 39200 11022 40000 6 io_oeb[10]
port 154 nsew signal tristate
rlabel metal2 s 11978 39200 12034 40000 6 io_oeb[11]
port 155 nsew signal tristate
rlabel metal2 s 13082 39200 13138 40000 6 io_oeb[12]
port 156 nsew signal tristate
rlabel metal2 s 14094 39200 14150 40000 6 io_oeb[13]
port 157 nsew signal tristate
rlabel metal2 s 15198 39200 15254 40000 6 io_oeb[14]
port 158 nsew signal tristate
rlabel metal2 s 16210 39200 16266 40000 6 io_oeb[15]
port 159 nsew signal tristate
rlabel metal2 s 17222 39200 17278 40000 6 io_oeb[16]
port 160 nsew signal tristate
rlabel metal2 s 18326 39200 18382 40000 6 io_oeb[17]
port 161 nsew signal tristate
rlabel metal2 s 19338 39200 19394 40000 6 io_oeb[18]
port 162 nsew signal tristate
rlabel metal2 s 20442 39200 20498 40000 6 io_oeb[19]
port 163 nsew signal tristate
rlabel metal2 s 1490 39200 1546 40000 6 io_oeb[1]
port 164 nsew signal tristate
rlabel metal2 s 21454 39200 21510 40000 6 io_oeb[20]
port 165 nsew signal tristate
rlabel metal2 s 22558 39200 22614 40000 6 io_oeb[21]
port 166 nsew signal tristate
rlabel metal2 s 23570 39200 23626 40000 6 io_oeb[22]
port 167 nsew signal tristate
rlabel metal2 s 24674 39200 24730 40000 6 io_oeb[23]
port 168 nsew signal tristate
rlabel metal2 s 25686 39200 25742 40000 6 io_oeb[24]
port 169 nsew signal tristate
rlabel metal2 s 26790 39200 26846 40000 6 io_oeb[25]
port 170 nsew signal tristate
rlabel metal2 s 27802 39200 27858 40000 6 io_oeb[26]
port 171 nsew signal tristate
rlabel metal2 s 28814 39200 28870 40000 6 io_oeb[27]
port 172 nsew signal tristate
rlabel metal2 s 29918 39200 29974 40000 6 io_oeb[28]
port 173 nsew signal tristate
rlabel metal2 s 30930 39200 30986 40000 6 io_oeb[29]
port 174 nsew signal tristate
rlabel metal2 s 2502 39200 2558 40000 6 io_oeb[2]
port 175 nsew signal tristate
rlabel metal2 s 32034 39200 32090 40000 6 io_oeb[30]
port 176 nsew signal tristate
rlabel metal2 s 33046 39200 33102 40000 6 io_oeb[31]
port 177 nsew signal tristate
rlabel metal2 s 34150 39200 34206 40000 6 io_oeb[32]
port 178 nsew signal tristate
rlabel metal2 s 35162 39200 35218 40000 6 io_oeb[33]
port 179 nsew signal tristate
rlabel metal2 s 36266 39200 36322 40000 6 io_oeb[34]
port 180 nsew signal tristate
rlabel metal2 s 37278 39200 37334 40000 6 io_oeb[35]
port 181 nsew signal tristate
rlabel metal2 s 38290 39200 38346 40000 6 io_oeb[36]
port 182 nsew signal tristate
rlabel metal2 s 39394 39200 39450 40000 6 io_oeb[37]
port 183 nsew signal tristate
rlabel metal2 s 3606 39200 3662 40000 6 io_oeb[3]
port 184 nsew signal tristate
rlabel metal2 s 4618 39200 4674 40000 6 io_oeb[4]
port 185 nsew signal tristate
rlabel metal2 s 5722 39200 5778 40000 6 io_oeb[5]
port 186 nsew signal tristate
rlabel metal2 s 6734 39200 6790 40000 6 io_oeb[6]
port 187 nsew signal tristate
rlabel metal2 s 7746 39200 7802 40000 6 io_oeb[7]
port 188 nsew signal tristate
rlabel metal2 s 8850 39200 8906 40000 6 io_oeb[8]
port 189 nsew signal tristate
rlabel metal2 s 9862 39200 9918 40000 6 io_oeb[9]
port 190 nsew signal tristate
rlabel metal2 s 754 39200 810 40000 6 io_out[0]
port 191 nsew signal tristate
rlabel metal2 s 11334 39200 11390 40000 6 io_out[10]
port 192 nsew signal tristate
rlabel metal2 s 12346 39200 12402 40000 6 io_out[11]
port 193 nsew signal tristate
rlabel metal2 s 13450 39200 13506 40000 6 io_out[12]
port 194 nsew signal tristate
rlabel metal2 s 14462 39200 14518 40000 6 io_out[13]
port 195 nsew signal tristate
rlabel metal2 s 15474 39200 15530 40000 6 io_out[14]
port 196 nsew signal tristate
rlabel metal2 s 16578 39200 16634 40000 6 io_out[15]
port 197 nsew signal tristate
rlabel metal2 s 17590 39200 17646 40000 6 io_out[16]
port 198 nsew signal tristate
rlabel metal2 s 18694 39200 18750 40000 6 io_out[17]
port 199 nsew signal tristate
rlabel metal2 s 19706 39200 19762 40000 6 io_out[18]
port 200 nsew signal tristate
rlabel metal2 s 20810 39200 20866 40000 6 io_out[19]
port 201 nsew signal tristate
rlabel metal2 s 1858 39200 1914 40000 6 io_out[1]
port 202 nsew signal tristate
rlabel metal2 s 21822 39200 21878 40000 6 io_out[20]
port 203 nsew signal tristate
rlabel metal2 s 22926 39200 22982 40000 6 io_out[21]
port 204 nsew signal tristate
rlabel metal2 s 23938 39200 23994 40000 6 io_out[22]
port 205 nsew signal tristate
rlabel metal2 s 24950 39200 25006 40000 6 io_out[23]
port 206 nsew signal tristate
rlabel metal2 s 26054 39200 26110 40000 6 io_out[24]
port 207 nsew signal tristate
rlabel metal2 s 27066 39200 27122 40000 6 io_out[25]
port 208 nsew signal tristate
rlabel metal2 s 28170 39200 28226 40000 6 io_out[26]
port 209 nsew signal tristate
rlabel metal2 s 29182 39200 29238 40000 6 io_out[27]
port 210 nsew signal tristate
rlabel metal2 s 30286 39200 30342 40000 6 io_out[28]
port 211 nsew signal tristate
rlabel metal2 s 31298 39200 31354 40000 6 io_out[29]
port 212 nsew signal tristate
rlabel metal2 s 2870 39200 2926 40000 6 io_out[2]
port 213 nsew signal tristate
rlabel metal2 s 32402 39200 32458 40000 6 io_out[30]
port 214 nsew signal tristate
rlabel metal2 s 33414 39200 33470 40000 6 io_out[31]
port 215 nsew signal tristate
rlabel metal2 s 34426 39200 34482 40000 6 io_out[32]
port 216 nsew signal tristate
rlabel metal2 s 35530 39200 35586 40000 6 io_out[33]
port 217 nsew signal tristate
rlabel metal2 s 36542 39200 36598 40000 6 io_out[34]
port 218 nsew signal tristate
rlabel metal2 s 37646 39200 37702 40000 6 io_out[35]
port 219 nsew signal tristate
rlabel metal2 s 38658 39200 38714 40000 6 io_out[36]
port 220 nsew signal tristate
rlabel metal2 s 39762 39200 39818 40000 6 io_out[37]
port 221 nsew signal tristate
rlabel metal2 s 3882 39200 3938 40000 6 io_out[3]
port 222 nsew signal tristate
rlabel metal2 s 4986 39200 5042 40000 6 io_out[4]
port 223 nsew signal tristate
rlabel metal2 s 5998 39200 6054 40000 6 io_out[5]
port 224 nsew signal tristate
rlabel metal2 s 7102 39200 7158 40000 6 io_out[6]
port 225 nsew signal tristate
rlabel metal2 s 8114 39200 8170 40000 6 io_out[7]
port 226 nsew signal tristate
rlabel metal2 s 9218 39200 9274 40000 6 io_out[8]
port 227 nsew signal tristate
rlabel metal2 s 10230 39200 10286 40000 6 io_out[9]
port 228 nsew signal tristate
rlabel metal3 s 39200 37408 40000 37528 6 la_blink[0]
port 229 nsew signal tristate
rlabel metal3 s 39200 39040 40000 39160 6 la_blink[1]
port 230 nsew signal tristate
rlabel metal2 s 110 0 166 800 6 pwm_en[0]
port 231 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 pwm_en[10]
port 232 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 pwm_en[11]
port 233 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 pwm_en[12]
port 234 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 pwm_en[13]
port 235 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 pwm_en[14]
port 236 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 pwm_en[15]
port 237 nsew signal input
rlabel metal2 s 570 0 626 800 6 pwm_en[1]
port 238 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 pwm_en[2]
port 239 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 pwm_en[3]
port 240 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 pwm_en[4]
port 241 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 pwm_en[5]
port 242 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 pwm_en[6]
port 243 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 pwm_en[7]
port 244 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 pwm_en[8]
port 245 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 pwm_en[9]
port 246 nsew signal input
rlabel metal2 s 294 0 350 800 6 pwm_out[0]
port 247 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 pwm_out[10]
port 248 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 pwm_out[11]
port 249 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 pwm_out[12]
port 250 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 pwm_out[13]
port 251 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 pwm_out[14]
port 252 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 pwm_out[15]
port 253 nsew signal input
rlabel metal2 s 846 0 902 800 6 pwm_out[1]
port 254 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 pwm_out[2]
port 255 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 pwm_out[3]
port 256 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 pwm_out[4]
port 257 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 pwm_out[5]
port 258 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 pwm_out[6]
port 259 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 pwm_out[7]
port 260 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 pwm_out[8]
port 261 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 pwm_out[9]
port 262 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 rst
port 263 nsew signal input
rlabel metal3 s 39200 20816 40000 20936 6 spi_clk[0]
port 264 nsew signal input
rlabel metal3 s 39200 29112 40000 29232 6 spi_clk[1]
port 265 nsew signal input
rlabel metal3 s 39200 22448 40000 22568 6 spi_cs[0]
port 266 nsew signal input
rlabel metal3 s 39200 30744 40000 30864 6 spi_cs[1]
port 267 nsew signal input
rlabel metal3 s 39200 24080 40000 24200 6 spi_en[0]
port 268 nsew signal input
rlabel metal3 s 39200 32376 40000 32496 6 spi_en[1]
port 269 nsew signal input
rlabel metal3 s 39200 25712 40000 25832 6 spi_miso[0]
port 270 nsew signal tristate
rlabel metal3 s 39200 34144 40000 34264 6 spi_miso[1]
port 271 nsew signal tristate
rlabel metal3 s 39200 27480 40000 27600 6 spi_mosi[0]
port 272 nsew signal input
rlabel metal3 s 39200 35776 40000 35896 6 spi_mosi[1]
port 273 nsew signal input
rlabel metal3 s 39200 824 40000 944 6 uart_en[0]
port 274 nsew signal input
rlabel metal3 s 39200 5720 40000 5840 6 uart_en[1]
port 275 nsew signal input
rlabel metal3 s 39200 10752 40000 10872 6 uart_en[2]
port 276 nsew signal input
rlabel metal3 s 39200 15784 40000 15904 6 uart_en[3]
port 277 nsew signal input
rlabel metal3 s 39200 2456 40000 2576 6 uart_rx[0]
port 278 nsew signal tristate
rlabel metal3 s 39200 7488 40000 7608 6 uart_rx[1]
port 279 nsew signal tristate
rlabel metal3 s 39200 12384 40000 12504 6 uart_rx[2]
port 280 nsew signal tristate
rlabel metal3 s 39200 17416 40000 17536 6 uart_rx[3]
port 281 nsew signal tristate
rlabel metal3 s 39200 4088 40000 4208 6 uart_tx[0]
port 282 nsew signal input
rlabel metal3 s 39200 9120 40000 9240 6 uart_tx[1]
port 283 nsew signal input
rlabel metal3 s 39200 14152 40000 14272 6 uart_tx[2]
port 284 nsew signal input
rlabel metal3 s 39200 19048 40000 19168 6 uart_tx[3]
port 285 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 286 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 286 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 287 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
