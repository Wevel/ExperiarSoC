magic
tech sky130A
magscale 1 2
timestamp 1652645824
<< obsli1 >>
rect 1104 2159 118864 97393
<< obsm1 >>
rect 474 1300 119494 98116
<< metal2 >>
rect 478 99200 534 100000
rect 1398 99200 1454 100000
rect 2318 99200 2374 100000
rect 3330 99200 3386 100000
rect 4250 99200 4306 100000
rect 5262 99200 5318 100000
rect 6182 99200 6238 100000
rect 7194 99200 7250 100000
rect 8114 99200 8170 100000
rect 9034 99200 9090 100000
rect 10046 99200 10102 100000
rect 10966 99200 11022 100000
rect 11978 99200 12034 100000
rect 12898 99200 12954 100000
rect 13910 99200 13966 100000
rect 14830 99200 14886 100000
rect 15750 99200 15806 100000
rect 16762 99200 16818 100000
rect 17682 99200 17738 100000
rect 18694 99200 18750 100000
rect 19614 99200 19670 100000
rect 20626 99200 20682 100000
rect 21546 99200 21602 100000
rect 22466 99200 22522 100000
rect 23478 99200 23534 100000
rect 24398 99200 24454 100000
rect 25410 99200 25466 100000
rect 26330 99200 26386 100000
rect 27342 99200 27398 100000
rect 28262 99200 28318 100000
rect 29182 99200 29238 100000
rect 30194 99200 30250 100000
rect 31114 99200 31170 100000
rect 32126 99200 32182 100000
rect 33046 99200 33102 100000
rect 34058 99200 34114 100000
rect 34978 99200 35034 100000
rect 35898 99200 35954 100000
rect 36910 99200 36966 100000
rect 37830 99200 37886 100000
rect 38842 99200 38898 100000
rect 39762 99200 39818 100000
rect 40774 99200 40830 100000
rect 41694 99200 41750 100000
rect 42706 99200 42762 100000
rect 43626 99200 43682 100000
rect 44546 99200 44602 100000
rect 45558 99200 45614 100000
rect 46478 99200 46534 100000
rect 47490 99200 47546 100000
rect 48410 99200 48466 100000
rect 49422 99200 49478 100000
rect 50342 99200 50398 100000
rect 51262 99200 51318 100000
rect 52274 99200 52330 100000
rect 53194 99200 53250 100000
rect 54206 99200 54262 100000
rect 55126 99200 55182 100000
rect 56138 99200 56194 100000
rect 57058 99200 57114 100000
rect 57978 99200 58034 100000
rect 58990 99200 59046 100000
rect 59910 99200 59966 100000
rect 60922 99200 60978 100000
rect 61842 99200 61898 100000
rect 62854 99200 62910 100000
rect 63774 99200 63830 100000
rect 64694 99200 64750 100000
rect 65706 99200 65762 100000
rect 66626 99200 66682 100000
rect 67638 99200 67694 100000
rect 68558 99200 68614 100000
rect 69570 99200 69626 100000
rect 70490 99200 70546 100000
rect 71410 99200 71466 100000
rect 72422 99200 72478 100000
rect 73342 99200 73398 100000
rect 74354 99200 74410 100000
rect 75274 99200 75330 100000
rect 76286 99200 76342 100000
rect 77206 99200 77262 100000
rect 78126 99200 78182 100000
rect 79138 99200 79194 100000
rect 80058 99200 80114 100000
rect 81070 99200 81126 100000
rect 81990 99200 82046 100000
rect 83002 99200 83058 100000
rect 83922 99200 83978 100000
rect 84934 99200 84990 100000
rect 85854 99200 85910 100000
rect 86774 99200 86830 100000
rect 87786 99200 87842 100000
rect 88706 99200 88762 100000
rect 89718 99200 89774 100000
rect 90638 99200 90694 100000
rect 91650 99200 91706 100000
rect 92570 99200 92626 100000
rect 93490 99200 93546 100000
rect 94502 99200 94558 100000
rect 95422 99200 95478 100000
rect 96434 99200 96490 100000
rect 97354 99200 97410 100000
rect 98366 99200 98422 100000
rect 99286 99200 99342 100000
rect 100206 99200 100262 100000
rect 101218 99200 101274 100000
rect 102138 99200 102194 100000
rect 103150 99200 103206 100000
rect 104070 99200 104126 100000
rect 105082 99200 105138 100000
rect 106002 99200 106058 100000
rect 106922 99200 106978 100000
rect 107934 99200 107990 100000
rect 108854 99200 108910 100000
rect 109866 99200 109922 100000
rect 110786 99200 110842 100000
rect 111798 99200 111854 100000
rect 112718 99200 112774 100000
rect 113638 99200 113694 100000
rect 114650 99200 114706 100000
rect 115570 99200 115626 100000
rect 116582 99200 116638 100000
rect 117502 99200 117558 100000
rect 118514 99200 118570 100000
rect 119434 99200 119490 100000
rect 1490 0 1546 800
rect 4434 0 4490 800
rect 7470 0 7526 800
rect 10414 0 10470 800
rect 13450 0 13506 800
rect 16486 0 16542 800
rect 19430 0 19486 800
rect 22466 0 22522 800
rect 25410 0 25466 800
rect 28446 0 28502 800
rect 31482 0 31538 800
rect 34426 0 34482 800
rect 37462 0 37518 800
rect 40406 0 40462 800
rect 43442 0 43498 800
rect 46478 0 46534 800
rect 49422 0 49478 800
rect 52458 0 52514 800
rect 55402 0 55458 800
rect 58438 0 58494 800
rect 61474 0 61530 800
rect 64418 0 64474 800
rect 67454 0 67510 800
rect 70398 0 70454 800
rect 73434 0 73490 800
rect 76470 0 76526 800
rect 79414 0 79470 800
rect 82450 0 82506 800
rect 85394 0 85450 800
rect 88430 0 88486 800
rect 91466 0 91522 800
rect 94410 0 94466 800
rect 97446 0 97502 800
rect 100390 0 100446 800
rect 103426 0 103482 800
rect 106462 0 106518 800
rect 109406 0 109462 800
rect 112442 0 112498 800
rect 115386 0 115442 800
rect 118422 0 118478 800
<< obsm2 >>
rect 590 99144 1342 99657
rect 1510 99144 2262 99657
rect 2430 99144 3274 99657
rect 3442 99144 4194 99657
rect 4362 99144 5206 99657
rect 5374 99144 6126 99657
rect 6294 99144 7138 99657
rect 7306 99144 8058 99657
rect 8226 99144 8978 99657
rect 9146 99144 9990 99657
rect 10158 99144 10910 99657
rect 11078 99144 11922 99657
rect 12090 99144 12842 99657
rect 13010 99144 13854 99657
rect 14022 99144 14774 99657
rect 14942 99144 15694 99657
rect 15862 99144 16706 99657
rect 16874 99144 17626 99657
rect 17794 99144 18638 99657
rect 18806 99144 19558 99657
rect 19726 99144 20570 99657
rect 20738 99144 21490 99657
rect 21658 99144 22410 99657
rect 22578 99144 23422 99657
rect 23590 99144 24342 99657
rect 24510 99144 25354 99657
rect 25522 99144 26274 99657
rect 26442 99144 27286 99657
rect 27454 99144 28206 99657
rect 28374 99144 29126 99657
rect 29294 99144 30138 99657
rect 30306 99144 31058 99657
rect 31226 99144 32070 99657
rect 32238 99144 32990 99657
rect 33158 99144 34002 99657
rect 34170 99144 34922 99657
rect 35090 99144 35842 99657
rect 36010 99144 36854 99657
rect 37022 99144 37774 99657
rect 37942 99144 38786 99657
rect 38954 99144 39706 99657
rect 39874 99144 40718 99657
rect 40886 99144 41638 99657
rect 41806 99144 42650 99657
rect 42818 99144 43570 99657
rect 43738 99144 44490 99657
rect 44658 99144 45502 99657
rect 45670 99144 46422 99657
rect 46590 99144 47434 99657
rect 47602 99144 48354 99657
rect 48522 99144 49366 99657
rect 49534 99144 50286 99657
rect 50454 99144 51206 99657
rect 51374 99144 52218 99657
rect 52386 99144 53138 99657
rect 53306 99144 54150 99657
rect 54318 99144 55070 99657
rect 55238 99144 56082 99657
rect 56250 99144 57002 99657
rect 57170 99144 57922 99657
rect 58090 99144 58934 99657
rect 59102 99144 59854 99657
rect 60022 99144 60866 99657
rect 61034 99144 61786 99657
rect 61954 99144 62798 99657
rect 62966 99144 63718 99657
rect 63886 99144 64638 99657
rect 64806 99144 65650 99657
rect 65818 99144 66570 99657
rect 66738 99144 67582 99657
rect 67750 99144 68502 99657
rect 68670 99144 69514 99657
rect 69682 99144 70434 99657
rect 70602 99144 71354 99657
rect 71522 99144 72366 99657
rect 72534 99144 73286 99657
rect 73454 99144 74298 99657
rect 74466 99144 75218 99657
rect 75386 99144 76230 99657
rect 76398 99144 77150 99657
rect 77318 99144 78070 99657
rect 78238 99144 79082 99657
rect 79250 99144 80002 99657
rect 80170 99144 81014 99657
rect 81182 99144 81934 99657
rect 82102 99144 82946 99657
rect 83114 99144 83866 99657
rect 84034 99144 84878 99657
rect 85046 99144 85798 99657
rect 85966 99144 86718 99657
rect 86886 99144 87730 99657
rect 87898 99144 88650 99657
rect 88818 99144 89662 99657
rect 89830 99144 90582 99657
rect 90750 99144 91594 99657
rect 91762 99144 92514 99657
rect 92682 99144 93434 99657
rect 93602 99144 94446 99657
rect 94614 99144 95366 99657
rect 95534 99144 96378 99657
rect 96546 99144 97298 99657
rect 97466 99144 98310 99657
rect 98478 99144 99230 99657
rect 99398 99144 100150 99657
rect 100318 99144 101162 99657
rect 101330 99144 102082 99657
rect 102250 99144 103094 99657
rect 103262 99144 104014 99657
rect 104182 99144 105026 99657
rect 105194 99144 105946 99657
rect 106114 99144 106866 99657
rect 107034 99144 107878 99657
rect 108046 99144 108798 99657
rect 108966 99144 109810 99657
rect 109978 99144 110730 99657
rect 110898 99144 111742 99657
rect 111910 99144 112662 99657
rect 112830 99144 113582 99657
rect 113750 99144 114594 99657
rect 114762 99144 115514 99657
rect 115682 99144 116526 99657
rect 116694 99144 117446 99657
rect 117614 99144 118458 99657
rect 118626 99144 119378 99657
rect 480 856 119488 99144
rect 480 167 1434 856
rect 1602 167 4378 856
rect 4546 167 7414 856
rect 7582 167 10358 856
rect 10526 167 13394 856
rect 13562 167 16430 856
rect 16598 167 19374 856
rect 19542 167 22410 856
rect 22578 167 25354 856
rect 25522 167 28390 856
rect 28558 167 31426 856
rect 31594 167 34370 856
rect 34538 167 37406 856
rect 37574 167 40350 856
rect 40518 167 43386 856
rect 43554 167 46422 856
rect 46590 167 49366 856
rect 49534 167 52402 856
rect 52570 167 55346 856
rect 55514 167 58382 856
rect 58550 167 61418 856
rect 61586 167 64362 856
rect 64530 167 67398 856
rect 67566 167 70342 856
rect 70510 167 73378 856
rect 73546 167 76414 856
rect 76582 167 79358 856
rect 79526 167 82394 856
rect 82562 167 85338 856
rect 85506 167 88374 856
rect 88542 167 91410 856
rect 91578 167 94354 856
rect 94522 167 97390 856
rect 97558 167 100334 856
rect 100502 167 103370 856
rect 103538 167 106406 856
rect 106574 167 109350 856
rect 109518 167 112386 856
rect 112554 167 115330 856
rect 115498 167 118366 856
rect 118534 167 119488 856
<< metal3 >>
rect 119200 99560 120000 99680
rect 0 98880 800 99000
rect 119200 99016 120000 99136
rect 119200 98608 120000 98728
rect 119200 98064 120000 98184
rect 119200 97520 120000 97640
rect 0 97112 800 97232
rect 119200 97112 120000 97232
rect 119200 96568 120000 96688
rect 119200 96160 120000 96280
rect 119200 95616 120000 95736
rect 0 95208 800 95328
rect 119200 95072 120000 95192
rect 119200 94664 120000 94784
rect 119200 94120 120000 94240
rect 0 93440 800 93560
rect 119200 93576 120000 93696
rect 119200 93168 120000 93288
rect 119200 92624 120000 92744
rect 119200 92216 120000 92336
rect 0 91672 800 91792
rect 119200 91672 120000 91792
rect 119200 91128 120000 91248
rect 119200 90720 120000 90840
rect 119200 90176 120000 90296
rect 0 89768 800 89888
rect 119200 89632 120000 89752
rect 119200 89224 120000 89344
rect 119200 88680 120000 88800
rect 119200 88272 120000 88392
rect 0 88000 800 88120
rect 119200 87728 120000 87848
rect 119200 87184 120000 87304
rect 119200 86776 120000 86896
rect 0 86232 800 86352
rect 119200 86232 120000 86352
rect 119200 85824 120000 85944
rect 119200 85280 120000 85400
rect 119200 84736 120000 84856
rect 0 84328 800 84448
rect 119200 84328 120000 84448
rect 119200 83784 120000 83904
rect 119200 83240 120000 83360
rect 119200 82832 120000 82952
rect 0 82560 800 82680
rect 119200 82288 120000 82408
rect 119200 81880 120000 82000
rect 119200 81336 120000 81456
rect 0 80792 800 80912
rect 119200 80792 120000 80912
rect 119200 80384 120000 80504
rect 119200 79840 120000 79960
rect 119200 79296 120000 79416
rect 0 78888 800 79008
rect 119200 78888 120000 79008
rect 119200 78344 120000 78464
rect 119200 77936 120000 78056
rect 119200 77392 120000 77512
rect 0 77120 800 77240
rect 119200 76848 120000 76968
rect 119200 76440 120000 76560
rect 119200 75896 120000 76016
rect 0 75216 800 75336
rect 119200 75352 120000 75472
rect 119200 74944 120000 75064
rect 119200 74400 120000 74520
rect 119200 73992 120000 74112
rect 0 73448 800 73568
rect 119200 73448 120000 73568
rect 119200 72904 120000 73024
rect 119200 72496 120000 72616
rect 119200 71952 120000 72072
rect 0 71680 800 71800
rect 119200 71544 120000 71664
rect 119200 71000 120000 71120
rect 119200 70456 120000 70576
rect 119200 70048 120000 70168
rect 0 69776 800 69896
rect 119200 69504 120000 69624
rect 119200 68960 120000 69080
rect 119200 68552 120000 68672
rect 0 68008 800 68128
rect 119200 68008 120000 68128
rect 119200 67600 120000 67720
rect 119200 67056 120000 67176
rect 119200 66512 120000 66632
rect 0 66240 800 66360
rect 119200 66104 120000 66224
rect 119200 65560 120000 65680
rect 119200 65016 120000 65136
rect 119200 64608 120000 64728
rect 0 64336 800 64456
rect 119200 64064 120000 64184
rect 119200 63656 120000 63776
rect 119200 63112 120000 63232
rect 0 62568 800 62688
rect 119200 62568 120000 62688
rect 119200 62160 120000 62280
rect 119200 61616 120000 61736
rect 119200 61072 120000 61192
rect 0 60800 800 60920
rect 119200 60664 120000 60784
rect 119200 60120 120000 60240
rect 119200 59712 120000 59832
rect 119200 59168 120000 59288
rect 0 58896 800 59016
rect 119200 58624 120000 58744
rect 119200 58216 120000 58336
rect 119200 57672 120000 57792
rect 0 57128 800 57248
rect 119200 57264 120000 57384
rect 119200 56720 120000 56840
rect 119200 56176 120000 56296
rect 119200 55768 120000 55888
rect 0 55224 800 55344
rect 119200 55224 120000 55344
rect 119200 54680 120000 54800
rect 119200 54272 120000 54392
rect 119200 53728 120000 53848
rect 0 53456 800 53576
rect 119200 53320 120000 53440
rect 119200 52776 120000 52896
rect 119200 52232 120000 52352
rect 0 51688 800 51808
rect 119200 51824 120000 51944
rect 119200 51280 120000 51400
rect 119200 50736 120000 50856
rect 119200 50328 120000 50448
rect 0 49784 800 49904
rect 119200 49784 120000 49904
rect 119200 49376 120000 49496
rect 119200 48832 120000 48952
rect 119200 48288 120000 48408
rect 0 48016 800 48136
rect 119200 47880 120000 48000
rect 119200 47336 120000 47456
rect 119200 46792 120000 46912
rect 0 46248 800 46368
rect 119200 46384 120000 46504
rect 119200 45840 120000 45960
rect 119200 45432 120000 45552
rect 119200 44888 120000 45008
rect 0 44344 800 44464
rect 119200 44344 120000 44464
rect 119200 43936 120000 44056
rect 119200 43392 120000 43512
rect 119200 42984 120000 43104
rect 0 42576 800 42696
rect 119200 42440 120000 42560
rect 119200 41896 120000 42016
rect 119200 41488 120000 41608
rect 0 40808 800 40928
rect 119200 40944 120000 41064
rect 119200 40400 120000 40520
rect 119200 39992 120000 40112
rect 119200 39448 120000 39568
rect 0 38904 800 39024
rect 119200 39040 120000 39160
rect 119200 38496 120000 38616
rect 119200 37952 120000 38072
rect 119200 37544 120000 37664
rect 0 37136 800 37256
rect 119200 37000 120000 37120
rect 119200 36456 120000 36576
rect 119200 36048 120000 36168
rect 119200 35504 120000 35624
rect 0 35232 800 35352
rect 119200 35096 120000 35216
rect 119200 34552 120000 34672
rect 119200 34008 120000 34128
rect 0 33464 800 33584
rect 119200 33600 120000 33720
rect 119200 33056 120000 33176
rect 119200 32512 120000 32632
rect 119200 32104 120000 32224
rect 0 31696 800 31816
rect 119200 31560 120000 31680
rect 119200 31152 120000 31272
rect 119200 30608 120000 30728
rect 119200 30064 120000 30184
rect 0 29792 800 29912
rect 119200 29656 120000 29776
rect 119200 29112 120000 29232
rect 119200 28704 120000 28824
rect 0 28024 800 28144
rect 119200 28160 120000 28280
rect 119200 27616 120000 27736
rect 119200 27208 120000 27328
rect 119200 26664 120000 26784
rect 0 26256 800 26376
rect 119200 26120 120000 26240
rect 119200 25712 120000 25832
rect 119200 25168 120000 25288
rect 119200 24760 120000 24880
rect 0 24352 800 24472
rect 119200 24216 120000 24336
rect 119200 23672 120000 23792
rect 119200 23264 120000 23384
rect 0 22584 800 22704
rect 119200 22720 120000 22840
rect 119200 22176 120000 22296
rect 119200 21768 120000 21888
rect 119200 21224 120000 21344
rect 0 20816 800 20936
rect 119200 20816 120000 20936
rect 119200 20272 120000 20392
rect 119200 19728 120000 19848
rect 119200 19320 120000 19440
rect 0 18912 800 19032
rect 119200 18776 120000 18896
rect 119200 18232 120000 18352
rect 119200 17824 120000 17944
rect 0 17144 800 17264
rect 119200 17280 120000 17400
rect 119200 16872 120000 16992
rect 119200 16328 120000 16448
rect 119200 15784 120000 15904
rect 0 15240 800 15360
rect 119200 15376 120000 15496
rect 119200 14832 120000 14952
rect 119200 14424 120000 14544
rect 119200 13880 120000 14000
rect 0 13472 800 13592
rect 119200 13336 120000 13456
rect 119200 12928 120000 13048
rect 119200 12384 120000 12504
rect 0 11704 800 11824
rect 119200 11840 120000 11960
rect 119200 11432 120000 11552
rect 119200 10888 120000 11008
rect 119200 10480 120000 10600
rect 0 9800 800 9920
rect 119200 9936 120000 10056
rect 119200 9392 120000 9512
rect 119200 8984 120000 9104
rect 119200 8440 120000 8560
rect 0 8032 800 8152
rect 119200 7896 120000 8016
rect 119200 7488 120000 7608
rect 119200 6944 120000 7064
rect 119200 6536 120000 6656
rect 0 6264 800 6384
rect 119200 5992 120000 6112
rect 119200 5448 120000 5568
rect 119200 5040 120000 5160
rect 0 4360 800 4480
rect 119200 4496 120000 4616
rect 119200 3952 120000 4072
rect 119200 3544 120000 3664
rect 119200 3000 120000 3120
rect 0 2592 800 2712
rect 119200 2592 120000 2712
rect 119200 2048 120000 2168
rect 119200 1504 120000 1624
rect 119200 1096 120000 1216
rect 0 824 800 944
rect 119200 552 120000 672
rect 119200 144 120000 264
<< obsm3 >>
rect 800 99480 119120 99653
rect 800 99216 119219 99480
rect 800 99080 119120 99216
rect 880 98936 119120 99080
rect 880 98808 119219 98936
rect 880 98800 119120 98808
rect 800 98528 119120 98800
rect 800 98264 119219 98528
rect 800 97984 119120 98264
rect 800 97720 119219 97984
rect 800 97440 119120 97720
rect 800 97312 119219 97440
rect 880 97032 119120 97312
rect 800 96768 119219 97032
rect 800 96488 119120 96768
rect 800 96360 119219 96488
rect 800 96080 119120 96360
rect 800 95816 119219 96080
rect 800 95536 119120 95816
rect 800 95408 119219 95536
rect 880 95272 119219 95408
rect 880 95128 119120 95272
rect 800 94992 119120 95128
rect 800 94864 119219 94992
rect 800 94584 119120 94864
rect 800 94320 119219 94584
rect 800 94040 119120 94320
rect 800 93776 119219 94040
rect 800 93640 119120 93776
rect 880 93496 119120 93640
rect 880 93368 119219 93496
rect 880 93360 119120 93368
rect 800 93088 119120 93360
rect 800 92824 119219 93088
rect 800 92544 119120 92824
rect 800 92416 119219 92544
rect 800 92136 119120 92416
rect 800 91872 119219 92136
rect 880 91592 119120 91872
rect 800 91328 119219 91592
rect 800 91048 119120 91328
rect 800 90920 119219 91048
rect 800 90640 119120 90920
rect 800 90376 119219 90640
rect 800 90096 119120 90376
rect 800 89968 119219 90096
rect 880 89832 119219 89968
rect 880 89688 119120 89832
rect 800 89552 119120 89688
rect 800 89424 119219 89552
rect 800 89144 119120 89424
rect 800 88880 119219 89144
rect 800 88600 119120 88880
rect 800 88472 119219 88600
rect 800 88200 119120 88472
rect 880 88192 119120 88200
rect 880 87928 119219 88192
rect 880 87920 119120 87928
rect 800 87648 119120 87920
rect 800 87384 119219 87648
rect 800 87104 119120 87384
rect 800 86976 119219 87104
rect 800 86696 119120 86976
rect 800 86432 119219 86696
rect 880 86152 119120 86432
rect 800 86024 119219 86152
rect 800 85744 119120 86024
rect 800 85480 119219 85744
rect 800 85200 119120 85480
rect 800 84936 119219 85200
rect 800 84656 119120 84936
rect 800 84528 119219 84656
rect 880 84248 119120 84528
rect 800 83984 119219 84248
rect 800 83704 119120 83984
rect 800 83440 119219 83704
rect 800 83160 119120 83440
rect 800 83032 119219 83160
rect 800 82760 119120 83032
rect 880 82752 119120 82760
rect 880 82488 119219 82752
rect 880 82480 119120 82488
rect 800 82208 119120 82480
rect 800 82080 119219 82208
rect 800 81800 119120 82080
rect 800 81536 119219 81800
rect 800 81256 119120 81536
rect 800 80992 119219 81256
rect 880 80712 119120 80992
rect 800 80584 119219 80712
rect 800 80304 119120 80584
rect 800 80040 119219 80304
rect 800 79760 119120 80040
rect 800 79496 119219 79760
rect 800 79216 119120 79496
rect 800 79088 119219 79216
rect 880 78808 119120 79088
rect 800 78544 119219 78808
rect 800 78264 119120 78544
rect 800 78136 119219 78264
rect 800 77856 119120 78136
rect 800 77592 119219 77856
rect 800 77320 119120 77592
rect 880 77312 119120 77320
rect 880 77048 119219 77312
rect 880 77040 119120 77048
rect 800 76768 119120 77040
rect 800 76640 119219 76768
rect 800 76360 119120 76640
rect 800 76096 119219 76360
rect 800 75816 119120 76096
rect 800 75552 119219 75816
rect 800 75416 119120 75552
rect 880 75272 119120 75416
rect 880 75144 119219 75272
rect 880 75136 119120 75144
rect 800 74864 119120 75136
rect 800 74600 119219 74864
rect 800 74320 119120 74600
rect 800 74192 119219 74320
rect 800 73912 119120 74192
rect 800 73648 119219 73912
rect 880 73368 119120 73648
rect 800 73104 119219 73368
rect 800 72824 119120 73104
rect 800 72696 119219 72824
rect 800 72416 119120 72696
rect 800 72152 119219 72416
rect 800 71880 119120 72152
rect 880 71872 119120 71880
rect 880 71744 119219 71872
rect 880 71600 119120 71744
rect 800 71464 119120 71600
rect 800 71200 119219 71464
rect 800 70920 119120 71200
rect 800 70656 119219 70920
rect 800 70376 119120 70656
rect 800 70248 119219 70376
rect 800 69976 119120 70248
rect 880 69968 119120 69976
rect 880 69704 119219 69968
rect 880 69696 119120 69704
rect 800 69424 119120 69696
rect 800 69160 119219 69424
rect 800 68880 119120 69160
rect 800 68752 119219 68880
rect 800 68472 119120 68752
rect 800 68208 119219 68472
rect 880 67928 119120 68208
rect 800 67800 119219 67928
rect 800 67520 119120 67800
rect 800 67256 119219 67520
rect 800 66976 119120 67256
rect 800 66712 119219 66976
rect 800 66440 119120 66712
rect 880 66432 119120 66440
rect 880 66304 119219 66432
rect 880 66160 119120 66304
rect 800 66024 119120 66160
rect 800 65760 119219 66024
rect 800 65480 119120 65760
rect 800 65216 119219 65480
rect 800 64936 119120 65216
rect 800 64808 119219 64936
rect 800 64536 119120 64808
rect 880 64528 119120 64536
rect 880 64264 119219 64528
rect 880 64256 119120 64264
rect 800 63984 119120 64256
rect 800 63856 119219 63984
rect 800 63576 119120 63856
rect 800 63312 119219 63576
rect 800 63032 119120 63312
rect 800 62768 119219 63032
rect 880 62488 119120 62768
rect 800 62360 119219 62488
rect 800 62080 119120 62360
rect 800 61816 119219 62080
rect 800 61536 119120 61816
rect 800 61272 119219 61536
rect 800 61000 119120 61272
rect 880 60992 119120 61000
rect 880 60864 119219 60992
rect 880 60720 119120 60864
rect 800 60584 119120 60720
rect 800 60320 119219 60584
rect 800 60040 119120 60320
rect 800 59912 119219 60040
rect 800 59632 119120 59912
rect 800 59368 119219 59632
rect 800 59096 119120 59368
rect 880 59088 119120 59096
rect 880 58824 119219 59088
rect 880 58816 119120 58824
rect 800 58544 119120 58816
rect 800 58416 119219 58544
rect 800 58136 119120 58416
rect 800 57872 119219 58136
rect 800 57592 119120 57872
rect 800 57464 119219 57592
rect 800 57328 119120 57464
rect 880 57184 119120 57328
rect 880 57048 119219 57184
rect 800 56920 119219 57048
rect 800 56640 119120 56920
rect 800 56376 119219 56640
rect 800 56096 119120 56376
rect 800 55968 119219 56096
rect 800 55688 119120 55968
rect 800 55424 119219 55688
rect 880 55144 119120 55424
rect 800 54880 119219 55144
rect 800 54600 119120 54880
rect 800 54472 119219 54600
rect 800 54192 119120 54472
rect 800 53928 119219 54192
rect 800 53656 119120 53928
rect 880 53648 119120 53656
rect 880 53520 119219 53648
rect 880 53376 119120 53520
rect 800 53240 119120 53376
rect 800 52976 119219 53240
rect 800 52696 119120 52976
rect 800 52432 119219 52696
rect 800 52152 119120 52432
rect 800 52024 119219 52152
rect 800 51888 119120 52024
rect 880 51744 119120 51888
rect 880 51608 119219 51744
rect 800 51480 119219 51608
rect 800 51200 119120 51480
rect 800 50936 119219 51200
rect 800 50656 119120 50936
rect 800 50528 119219 50656
rect 800 50248 119120 50528
rect 800 49984 119219 50248
rect 880 49704 119120 49984
rect 800 49576 119219 49704
rect 800 49296 119120 49576
rect 800 49032 119219 49296
rect 800 48752 119120 49032
rect 800 48488 119219 48752
rect 800 48216 119120 48488
rect 880 48208 119120 48216
rect 880 48080 119219 48208
rect 880 47936 119120 48080
rect 800 47800 119120 47936
rect 800 47536 119219 47800
rect 800 47256 119120 47536
rect 800 46992 119219 47256
rect 800 46712 119120 46992
rect 800 46584 119219 46712
rect 800 46448 119120 46584
rect 880 46304 119120 46448
rect 880 46168 119219 46304
rect 800 46040 119219 46168
rect 800 45760 119120 46040
rect 800 45632 119219 45760
rect 800 45352 119120 45632
rect 800 45088 119219 45352
rect 800 44808 119120 45088
rect 800 44544 119219 44808
rect 880 44264 119120 44544
rect 800 44136 119219 44264
rect 800 43856 119120 44136
rect 800 43592 119219 43856
rect 800 43312 119120 43592
rect 800 43184 119219 43312
rect 800 42904 119120 43184
rect 800 42776 119219 42904
rect 880 42640 119219 42776
rect 880 42496 119120 42640
rect 800 42360 119120 42496
rect 800 42096 119219 42360
rect 800 41816 119120 42096
rect 800 41688 119219 41816
rect 800 41408 119120 41688
rect 800 41144 119219 41408
rect 800 41008 119120 41144
rect 880 40864 119120 41008
rect 880 40728 119219 40864
rect 800 40600 119219 40728
rect 800 40320 119120 40600
rect 800 40192 119219 40320
rect 800 39912 119120 40192
rect 800 39648 119219 39912
rect 800 39368 119120 39648
rect 800 39240 119219 39368
rect 800 39104 119120 39240
rect 880 38960 119120 39104
rect 880 38824 119219 38960
rect 800 38696 119219 38824
rect 800 38416 119120 38696
rect 800 38152 119219 38416
rect 800 37872 119120 38152
rect 800 37744 119219 37872
rect 800 37464 119120 37744
rect 800 37336 119219 37464
rect 880 37200 119219 37336
rect 880 37056 119120 37200
rect 800 36920 119120 37056
rect 800 36656 119219 36920
rect 800 36376 119120 36656
rect 800 36248 119219 36376
rect 800 35968 119120 36248
rect 800 35704 119219 35968
rect 800 35432 119120 35704
rect 880 35424 119120 35432
rect 880 35296 119219 35424
rect 880 35152 119120 35296
rect 800 35016 119120 35152
rect 800 34752 119219 35016
rect 800 34472 119120 34752
rect 800 34208 119219 34472
rect 800 33928 119120 34208
rect 800 33800 119219 33928
rect 800 33664 119120 33800
rect 880 33520 119120 33664
rect 880 33384 119219 33520
rect 800 33256 119219 33384
rect 800 32976 119120 33256
rect 800 32712 119219 32976
rect 800 32432 119120 32712
rect 800 32304 119219 32432
rect 800 32024 119120 32304
rect 800 31896 119219 32024
rect 880 31760 119219 31896
rect 880 31616 119120 31760
rect 800 31480 119120 31616
rect 800 31352 119219 31480
rect 800 31072 119120 31352
rect 800 30808 119219 31072
rect 800 30528 119120 30808
rect 800 30264 119219 30528
rect 800 29992 119120 30264
rect 880 29984 119120 29992
rect 880 29856 119219 29984
rect 880 29712 119120 29856
rect 800 29576 119120 29712
rect 800 29312 119219 29576
rect 800 29032 119120 29312
rect 800 28904 119219 29032
rect 800 28624 119120 28904
rect 800 28360 119219 28624
rect 800 28224 119120 28360
rect 880 28080 119120 28224
rect 880 27944 119219 28080
rect 800 27816 119219 27944
rect 800 27536 119120 27816
rect 800 27408 119219 27536
rect 800 27128 119120 27408
rect 800 26864 119219 27128
rect 800 26584 119120 26864
rect 800 26456 119219 26584
rect 880 26320 119219 26456
rect 880 26176 119120 26320
rect 800 26040 119120 26176
rect 800 25912 119219 26040
rect 800 25632 119120 25912
rect 800 25368 119219 25632
rect 800 25088 119120 25368
rect 800 24960 119219 25088
rect 800 24680 119120 24960
rect 800 24552 119219 24680
rect 880 24416 119219 24552
rect 880 24272 119120 24416
rect 800 24136 119120 24272
rect 800 23872 119219 24136
rect 800 23592 119120 23872
rect 800 23464 119219 23592
rect 800 23184 119120 23464
rect 800 22920 119219 23184
rect 800 22784 119120 22920
rect 880 22640 119120 22784
rect 880 22504 119219 22640
rect 800 22376 119219 22504
rect 800 22096 119120 22376
rect 800 21968 119219 22096
rect 800 21688 119120 21968
rect 800 21424 119219 21688
rect 800 21144 119120 21424
rect 800 21016 119219 21144
rect 880 20736 119120 21016
rect 800 20472 119219 20736
rect 800 20192 119120 20472
rect 800 19928 119219 20192
rect 800 19648 119120 19928
rect 800 19520 119219 19648
rect 800 19240 119120 19520
rect 800 19112 119219 19240
rect 880 18976 119219 19112
rect 880 18832 119120 18976
rect 800 18696 119120 18832
rect 800 18432 119219 18696
rect 800 18152 119120 18432
rect 800 18024 119219 18152
rect 800 17744 119120 18024
rect 800 17480 119219 17744
rect 800 17344 119120 17480
rect 880 17200 119120 17344
rect 880 17072 119219 17200
rect 880 17064 119120 17072
rect 800 16792 119120 17064
rect 800 16528 119219 16792
rect 800 16248 119120 16528
rect 800 15984 119219 16248
rect 800 15704 119120 15984
rect 800 15576 119219 15704
rect 800 15440 119120 15576
rect 880 15296 119120 15440
rect 880 15160 119219 15296
rect 800 15032 119219 15160
rect 800 14752 119120 15032
rect 800 14624 119219 14752
rect 800 14344 119120 14624
rect 800 14080 119219 14344
rect 800 13800 119120 14080
rect 800 13672 119219 13800
rect 880 13536 119219 13672
rect 880 13392 119120 13536
rect 800 13256 119120 13392
rect 800 13128 119219 13256
rect 800 12848 119120 13128
rect 800 12584 119219 12848
rect 800 12304 119120 12584
rect 800 12040 119219 12304
rect 800 11904 119120 12040
rect 880 11760 119120 11904
rect 880 11632 119219 11760
rect 880 11624 119120 11632
rect 800 11352 119120 11624
rect 800 11088 119219 11352
rect 800 10808 119120 11088
rect 800 10680 119219 10808
rect 800 10400 119120 10680
rect 800 10136 119219 10400
rect 800 10000 119120 10136
rect 880 9856 119120 10000
rect 880 9720 119219 9856
rect 800 9592 119219 9720
rect 800 9312 119120 9592
rect 800 9184 119219 9312
rect 800 8904 119120 9184
rect 800 8640 119219 8904
rect 800 8360 119120 8640
rect 800 8232 119219 8360
rect 880 8096 119219 8232
rect 880 7952 119120 8096
rect 800 7816 119120 7952
rect 800 7688 119219 7816
rect 800 7408 119120 7688
rect 800 7144 119219 7408
rect 800 6864 119120 7144
rect 800 6736 119219 6864
rect 800 6464 119120 6736
rect 880 6456 119120 6464
rect 880 6192 119219 6456
rect 880 6184 119120 6192
rect 800 5912 119120 6184
rect 800 5648 119219 5912
rect 800 5368 119120 5648
rect 800 5240 119219 5368
rect 800 4960 119120 5240
rect 800 4696 119219 4960
rect 800 4560 119120 4696
rect 880 4416 119120 4560
rect 880 4280 119219 4416
rect 800 4152 119219 4280
rect 800 3872 119120 4152
rect 800 3744 119219 3872
rect 800 3464 119120 3744
rect 800 3200 119219 3464
rect 800 2920 119120 3200
rect 800 2792 119219 2920
rect 880 2512 119120 2792
rect 800 2248 119219 2512
rect 800 1968 119120 2248
rect 800 1704 119219 1968
rect 800 1424 119120 1704
rect 800 1296 119219 1424
rect 800 1024 119120 1296
rect 880 1016 119120 1024
rect 880 752 119219 1016
rect 880 744 119120 752
rect 800 472 119120 744
rect 800 344 119219 472
rect 800 171 119120 344
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
rect 111728 2128 112048 97424
<< obsm4 >>
rect 20115 4523 34848 96661
rect 35328 4523 50208 96661
rect 50688 4523 65568 96661
rect 66048 4523 80928 96661
rect 81408 4523 96288 96661
rect 96768 4523 111648 96661
rect 112128 4523 116597 96661
<< labels >>
rlabel metal2 s 7194 99200 7250 100000 6 addr0[0]
port 1 nsew signal output
rlabel metal2 s 8114 99200 8170 100000 6 addr0[1]
port 2 nsew signal output
rlabel metal2 s 9034 99200 9090 100000 6 addr0[2]
port 3 nsew signal output
rlabel metal2 s 10046 99200 10102 100000 6 addr0[3]
port 4 nsew signal output
rlabel metal2 s 10966 99200 11022 100000 6 addr0[4]
port 5 nsew signal output
rlabel metal2 s 11978 99200 12034 100000 6 addr0[5]
port 6 nsew signal output
rlabel metal2 s 12898 99200 12954 100000 6 addr0[6]
port 7 nsew signal output
rlabel metal2 s 13910 99200 13966 100000 6 addr0[7]
port 8 nsew signal output
rlabel metal2 s 14830 99200 14886 100000 6 addr0[8]
port 9 nsew signal output
rlabel metal2 s 79138 99200 79194 100000 6 addr1[0]
port 10 nsew signal output
rlabel metal2 s 80058 99200 80114 100000 6 addr1[1]
port 11 nsew signal output
rlabel metal2 s 81070 99200 81126 100000 6 addr1[2]
port 12 nsew signal output
rlabel metal2 s 81990 99200 82046 100000 6 addr1[3]
port 13 nsew signal output
rlabel metal2 s 83002 99200 83058 100000 6 addr1[4]
port 14 nsew signal output
rlabel metal2 s 83922 99200 83978 100000 6 addr1[5]
port 15 nsew signal output
rlabel metal2 s 84934 99200 84990 100000 6 addr1[6]
port 16 nsew signal output
rlabel metal2 s 85854 99200 85910 100000 6 addr1[7]
port 17 nsew signal output
rlabel metal2 s 86774 99200 86830 100000 6 addr1[8]
port 18 nsew signal output
rlabel metal2 s 478 99200 534 100000 6 clk0
port 19 nsew signal output
rlabel metal2 s 77206 99200 77262 100000 6 clk1
port 20 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 119200 1096 120000 1216 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 119200 3952 120000 4072 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 119200 20816 120000 20936 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 119200 22176 120000 22296 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 119200 23672 120000 23792 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 119200 25168 120000 25288 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 119200 26664 120000 26784 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 119200 28160 120000 28280 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 119200 29656 120000 29776 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 119200 31152 120000 31272 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 119200 32512 120000 32632 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 119200 34008 120000 34128 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 119200 5992 120000 6112 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 119200 35504 120000 35624 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 119200 37000 120000 37120 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 119200 38496 120000 38616 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 119200 39992 120000 40112 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 119200 41488 120000 41608 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 119200 42984 120000 43104 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 119200 44344 120000 44464 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 119200 45840 120000 45960 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 119200 7896 120000 8016 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 119200 9936 120000 10056 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 119200 11840 120000 11960 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 119200 13336 120000 13456 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 119200 14832 120000 14952 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 119200 16328 120000 16448 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 119200 17824 120000 17944 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 119200 19320 120000 19440 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 119200 1504 120000 1624 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 119200 4496 120000 4616 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 119200 21224 120000 21344 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 119200 22720 120000 22840 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 119200 24216 120000 24336 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 119200 25712 120000 25832 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 119200 27208 120000 27328 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 119200 28704 120000 28824 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 119200 30064 120000 30184 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 119200 31560 120000 31680 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 119200 33056 120000 33176 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 119200 34552 120000 34672 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 119200 6536 120000 6656 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 119200 36048 120000 36168 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 119200 37544 120000 37664 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 119200 39040 120000 39160 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 119200 40400 120000 40520 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 119200 41896 120000 42016 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 119200 43392 120000 43512 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 119200 44888 120000 45008 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 119200 46384 120000 46504 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 119200 47336 120000 47456 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 119200 48288 120000 48408 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 119200 8440 120000 8560 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 119200 49376 120000 49496 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 119200 50328 120000 50448 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 119200 10480 120000 10600 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 119200 12384 120000 12504 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 119200 13880 120000 14000 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 119200 15376 120000 15496 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 119200 16872 120000 16992 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 119200 18232 120000 18352 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 119200 19728 120000 19848 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 119200 5040 120000 5160 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 119200 21768 120000 21888 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 119200 23264 120000 23384 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 119200 24760 120000 24880 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 119200 26120 120000 26240 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 119200 27616 120000 27736 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 119200 29112 120000 29232 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 119200 30608 120000 30728 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 119200 32104 120000 32224 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 119200 33600 120000 33720 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 119200 35096 120000 35216 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 119200 6944 120000 7064 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 119200 36456 120000 36576 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 119200 37952 120000 38072 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 119200 39448 120000 39568 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 119200 40944 120000 41064 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 119200 42440 120000 42560 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 119200 43936 120000 44056 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 119200 45432 120000 45552 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 119200 46792 120000 46912 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 119200 47880 120000 48000 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 119200 48832 120000 48952 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 119200 8984 120000 9104 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 119200 49784 120000 49904 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 119200 50736 120000 50856 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 119200 10888 120000 11008 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 119200 12928 120000 13048 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 119200 14424 120000 14544 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 119200 15784 120000 15904 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 119200 17280 120000 17400 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 119200 18776 120000 18896 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 119200 20272 120000 20392 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 119200 2048 120000 2168 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 119200 5448 120000 5568 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 119200 7488 120000 7608 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 119200 9392 120000 9512 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 119200 11432 120000 11552 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 119200 2592 120000 2712 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 119200 3000 120000 3120 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 119200 3544 120000 3664 6 core_wb_we_o
port 130 nsew signal output
rlabel metal2 s 1398 99200 1454 100000 6 csb0
port 131 nsew signal output
rlabel metal2 s 78126 99200 78182 100000 6 csb1
port 132 nsew signal output
rlabel metal2 s 15750 99200 15806 100000 6 din0[0]
port 133 nsew signal output
rlabel metal2 s 25410 99200 25466 100000 6 din0[10]
port 134 nsew signal output
rlabel metal2 s 26330 99200 26386 100000 6 din0[11]
port 135 nsew signal output
rlabel metal2 s 27342 99200 27398 100000 6 din0[12]
port 136 nsew signal output
rlabel metal2 s 28262 99200 28318 100000 6 din0[13]
port 137 nsew signal output
rlabel metal2 s 29182 99200 29238 100000 6 din0[14]
port 138 nsew signal output
rlabel metal2 s 30194 99200 30250 100000 6 din0[15]
port 139 nsew signal output
rlabel metal2 s 31114 99200 31170 100000 6 din0[16]
port 140 nsew signal output
rlabel metal2 s 32126 99200 32182 100000 6 din0[17]
port 141 nsew signal output
rlabel metal2 s 33046 99200 33102 100000 6 din0[18]
port 142 nsew signal output
rlabel metal2 s 34058 99200 34114 100000 6 din0[19]
port 143 nsew signal output
rlabel metal2 s 16762 99200 16818 100000 6 din0[1]
port 144 nsew signal output
rlabel metal2 s 34978 99200 35034 100000 6 din0[20]
port 145 nsew signal output
rlabel metal2 s 35898 99200 35954 100000 6 din0[21]
port 146 nsew signal output
rlabel metal2 s 36910 99200 36966 100000 6 din0[22]
port 147 nsew signal output
rlabel metal2 s 37830 99200 37886 100000 6 din0[23]
port 148 nsew signal output
rlabel metal2 s 38842 99200 38898 100000 6 din0[24]
port 149 nsew signal output
rlabel metal2 s 39762 99200 39818 100000 6 din0[25]
port 150 nsew signal output
rlabel metal2 s 40774 99200 40830 100000 6 din0[26]
port 151 nsew signal output
rlabel metal2 s 41694 99200 41750 100000 6 din0[27]
port 152 nsew signal output
rlabel metal2 s 42706 99200 42762 100000 6 din0[28]
port 153 nsew signal output
rlabel metal2 s 43626 99200 43682 100000 6 din0[29]
port 154 nsew signal output
rlabel metal2 s 17682 99200 17738 100000 6 din0[2]
port 155 nsew signal output
rlabel metal2 s 44546 99200 44602 100000 6 din0[30]
port 156 nsew signal output
rlabel metal2 s 45558 99200 45614 100000 6 din0[31]
port 157 nsew signal output
rlabel metal2 s 18694 99200 18750 100000 6 din0[3]
port 158 nsew signal output
rlabel metal2 s 19614 99200 19670 100000 6 din0[4]
port 159 nsew signal output
rlabel metal2 s 20626 99200 20682 100000 6 din0[5]
port 160 nsew signal output
rlabel metal2 s 21546 99200 21602 100000 6 din0[6]
port 161 nsew signal output
rlabel metal2 s 22466 99200 22522 100000 6 din0[7]
port 162 nsew signal output
rlabel metal2 s 23478 99200 23534 100000 6 din0[8]
port 163 nsew signal output
rlabel metal2 s 24398 99200 24454 100000 6 din0[9]
port 164 nsew signal output
rlabel metal2 s 46478 99200 46534 100000 6 dout0[0]
port 165 nsew signal input
rlabel metal2 s 56138 99200 56194 100000 6 dout0[10]
port 166 nsew signal input
rlabel metal2 s 57058 99200 57114 100000 6 dout0[11]
port 167 nsew signal input
rlabel metal2 s 57978 99200 58034 100000 6 dout0[12]
port 168 nsew signal input
rlabel metal2 s 58990 99200 59046 100000 6 dout0[13]
port 169 nsew signal input
rlabel metal2 s 59910 99200 59966 100000 6 dout0[14]
port 170 nsew signal input
rlabel metal2 s 60922 99200 60978 100000 6 dout0[15]
port 171 nsew signal input
rlabel metal2 s 61842 99200 61898 100000 6 dout0[16]
port 172 nsew signal input
rlabel metal2 s 62854 99200 62910 100000 6 dout0[17]
port 173 nsew signal input
rlabel metal2 s 63774 99200 63830 100000 6 dout0[18]
port 174 nsew signal input
rlabel metal2 s 64694 99200 64750 100000 6 dout0[19]
port 175 nsew signal input
rlabel metal2 s 47490 99200 47546 100000 6 dout0[1]
port 176 nsew signal input
rlabel metal2 s 65706 99200 65762 100000 6 dout0[20]
port 177 nsew signal input
rlabel metal2 s 66626 99200 66682 100000 6 dout0[21]
port 178 nsew signal input
rlabel metal2 s 67638 99200 67694 100000 6 dout0[22]
port 179 nsew signal input
rlabel metal2 s 68558 99200 68614 100000 6 dout0[23]
port 180 nsew signal input
rlabel metal2 s 69570 99200 69626 100000 6 dout0[24]
port 181 nsew signal input
rlabel metal2 s 70490 99200 70546 100000 6 dout0[25]
port 182 nsew signal input
rlabel metal2 s 71410 99200 71466 100000 6 dout0[26]
port 183 nsew signal input
rlabel metal2 s 72422 99200 72478 100000 6 dout0[27]
port 184 nsew signal input
rlabel metal2 s 73342 99200 73398 100000 6 dout0[28]
port 185 nsew signal input
rlabel metal2 s 74354 99200 74410 100000 6 dout0[29]
port 186 nsew signal input
rlabel metal2 s 48410 99200 48466 100000 6 dout0[2]
port 187 nsew signal input
rlabel metal2 s 75274 99200 75330 100000 6 dout0[30]
port 188 nsew signal input
rlabel metal2 s 76286 99200 76342 100000 6 dout0[31]
port 189 nsew signal input
rlabel metal2 s 49422 99200 49478 100000 6 dout0[3]
port 190 nsew signal input
rlabel metal2 s 50342 99200 50398 100000 6 dout0[4]
port 191 nsew signal input
rlabel metal2 s 51262 99200 51318 100000 6 dout0[5]
port 192 nsew signal input
rlabel metal2 s 52274 99200 52330 100000 6 dout0[6]
port 193 nsew signal input
rlabel metal2 s 53194 99200 53250 100000 6 dout0[7]
port 194 nsew signal input
rlabel metal2 s 54206 99200 54262 100000 6 dout0[8]
port 195 nsew signal input
rlabel metal2 s 55126 99200 55182 100000 6 dout0[9]
port 196 nsew signal input
rlabel metal2 s 87786 99200 87842 100000 6 dout1[0]
port 197 nsew signal input
rlabel metal2 s 97354 99200 97410 100000 6 dout1[10]
port 198 nsew signal input
rlabel metal2 s 98366 99200 98422 100000 6 dout1[11]
port 199 nsew signal input
rlabel metal2 s 99286 99200 99342 100000 6 dout1[12]
port 200 nsew signal input
rlabel metal2 s 100206 99200 100262 100000 6 dout1[13]
port 201 nsew signal input
rlabel metal2 s 101218 99200 101274 100000 6 dout1[14]
port 202 nsew signal input
rlabel metal2 s 102138 99200 102194 100000 6 dout1[15]
port 203 nsew signal input
rlabel metal2 s 103150 99200 103206 100000 6 dout1[16]
port 204 nsew signal input
rlabel metal2 s 104070 99200 104126 100000 6 dout1[17]
port 205 nsew signal input
rlabel metal2 s 105082 99200 105138 100000 6 dout1[18]
port 206 nsew signal input
rlabel metal2 s 106002 99200 106058 100000 6 dout1[19]
port 207 nsew signal input
rlabel metal2 s 88706 99200 88762 100000 6 dout1[1]
port 208 nsew signal input
rlabel metal2 s 106922 99200 106978 100000 6 dout1[20]
port 209 nsew signal input
rlabel metal2 s 107934 99200 107990 100000 6 dout1[21]
port 210 nsew signal input
rlabel metal2 s 108854 99200 108910 100000 6 dout1[22]
port 211 nsew signal input
rlabel metal2 s 109866 99200 109922 100000 6 dout1[23]
port 212 nsew signal input
rlabel metal2 s 110786 99200 110842 100000 6 dout1[24]
port 213 nsew signal input
rlabel metal2 s 111798 99200 111854 100000 6 dout1[25]
port 214 nsew signal input
rlabel metal2 s 112718 99200 112774 100000 6 dout1[26]
port 215 nsew signal input
rlabel metal2 s 113638 99200 113694 100000 6 dout1[27]
port 216 nsew signal input
rlabel metal2 s 114650 99200 114706 100000 6 dout1[28]
port 217 nsew signal input
rlabel metal2 s 115570 99200 115626 100000 6 dout1[29]
port 218 nsew signal input
rlabel metal2 s 89718 99200 89774 100000 6 dout1[2]
port 219 nsew signal input
rlabel metal2 s 116582 99200 116638 100000 6 dout1[30]
port 220 nsew signal input
rlabel metal2 s 117502 99200 117558 100000 6 dout1[31]
port 221 nsew signal input
rlabel metal2 s 90638 99200 90694 100000 6 dout1[3]
port 222 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 dout1[4]
port 223 nsew signal input
rlabel metal2 s 92570 99200 92626 100000 6 dout1[5]
port 224 nsew signal input
rlabel metal2 s 93490 99200 93546 100000 6 dout1[6]
port 225 nsew signal input
rlabel metal2 s 94502 99200 94558 100000 6 dout1[7]
port 226 nsew signal input
rlabel metal2 s 95422 99200 95478 100000 6 dout1[8]
port 227 nsew signal input
rlabel metal2 s 96434 99200 96490 100000 6 dout1[9]
port 228 nsew signal input
rlabel metal2 s 118514 99200 118570 100000 6 jtag_tck
port 229 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 jtag_tdi
port 230 nsew signal input
rlabel metal2 s 119434 99200 119490 100000 6 jtag_tdo
port 231 nsew signal output
rlabel metal3 s 119200 99560 120000 99680 6 jtag_tms
port 232 nsew signal input
rlabel metal3 s 119200 51280 120000 51400 6 localMemory_wb_ack_o
port 233 nsew signal output
rlabel metal3 s 119200 54272 120000 54392 6 localMemory_wb_adr_i[0]
port 234 nsew signal input
rlabel metal3 s 119200 71000 120000 71120 6 localMemory_wb_adr_i[10]
port 235 nsew signal input
rlabel metal3 s 119200 72496 120000 72616 6 localMemory_wb_adr_i[11]
port 236 nsew signal input
rlabel metal3 s 119200 73992 120000 74112 6 localMemory_wb_adr_i[12]
port 237 nsew signal input
rlabel metal3 s 119200 75352 120000 75472 6 localMemory_wb_adr_i[13]
port 238 nsew signal input
rlabel metal3 s 119200 76848 120000 76968 6 localMemory_wb_adr_i[14]
port 239 nsew signal input
rlabel metal3 s 119200 78344 120000 78464 6 localMemory_wb_adr_i[15]
port 240 nsew signal input
rlabel metal3 s 119200 79840 120000 79960 6 localMemory_wb_adr_i[16]
port 241 nsew signal input
rlabel metal3 s 119200 81336 120000 81456 6 localMemory_wb_adr_i[17]
port 242 nsew signal input
rlabel metal3 s 119200 82832 120000 82952 6 localMemory_wb_adr_i[18]
port 243 nsew signal input
rlabel metal3 s 119200 84328 120000 84448 6 localMemory_wb_adr_i[19]
port 244 nsew signal input
rlabel metal3 s 119200 56176 120000 56296 6 localMemory_wb_adr_i[1]
port 245 nsew signal input
rlabel metal3 s 119200 85824 120000 85944 6 localMemory_wb_adr_i[20]
port 246 nsew signal input
rlabel metal3 s 119200 87184 120000 87304 6 localMemory_wb_adr_i[21]
port 247 nsew signal input
rlabel metal3 s 119200 88680 120000 88800 6 localMemory_wb_adr_i[22]
port 248 nsew signal input
rlabel metal3 s 119200 90176 120000 90296 6 localMemory_wb_adr_i[23]
port 249 nsew signal input
rlabel metal3 s 119200 58216 120000 58336 6 localMemory_wb_adr_i[2]
port 250 nsew signal input
rlabel metal3 s 119200 60120 120000 60240 6 localMemory_wb_adr_i[3]
port 251 nsew signal input
rlabel metal3 s 119200 62160 120000 62280 6 localMemory_wb_adr_i[4]
port 252 nsew signal input
rlabel metal3 s 119200 63656 120000 63776 6 localMemory_wb_adr_i[5]
port 253 nsew signal input
rlabel metal3 s 119200 65016 120000 65136 6 localMemory_wb_adr_i[6]
port 254 nsew signal input
rlabel metal3 s 119200 66512 120000 66632 6 localMemory_wb_adr_i[7]
port 255 nsew signal input
rlabel metal3 s 119200 68008 120000 68128 6 localMemory_wb_adr_i[8]
port 256 nsew signal input
rlabel metal3 s 119200 69504 120000 69624 6 localMemory_wb_adr_i[9]
port 257 nsew signal input
rlabel metal3 s 119200 51824 120000 51944 6 localMemory_wb_cyc_i
port 258 nsew signal input
rlabel metal3 s 119200 54680 120000 54800 6 localMemory_wb_data_i[0]
port 259 nsew signal input
rlabel metal3 s 119200 71544 120000 71664 6 localMemory_wb_data_i[10]
port 260 nsew signal input
rlabel metal3 s 119200 72904 120000 73024 6 localMemory_wb_data_i[11]
port 261 nsew signal input
rlabel metal3 s 119200 74400 120000 74520 6 localMemory_wb_data_i[12]
port 262 nsew signal input
rlabel metal3 s 119200 75896 120000 76016 6 localMemory_wb_data_i[13]
port 263 nsew signal input
rlabel metal3 s 119200 77392 120000 77512 6 localMemory_wb_data_i[14]
port 264 nsew signal input
rlabel metal3 s 119200 78888 120000 79008 6 localMemory_wb_data_i[15]
port 265 nsew signal input
rlabel metal3 s 119200 80384 120000 80504 6 localMemory_wb_data_i[16]
port 266 nsew signal input
rlabel metal3 s 119200 81880 120000 82000 6 localMemory_wb_data_i[17]
port 267 nsew signal input
rlabel metal3 s 119200 83240 120000 83360 6 localMemory_wb_data_i[18]
port 268 nsew signal input
rlabel metal3 s 119200 84736 120000 84856 6 localMemory_wb_data_i[19]
port 269 nsew signal input
rlabel metal3 s 119200 56720 120000 56840 6 localMemory_wb_data_i[1]
port 270 nsew signal input
rlabel metal3 s 119200 86232 120000 86352 6 localMemory_wb_data_i[20]
port 271 nsew signal input
rlabel metal3 s 119200 87728 120000 87848 6 localMemory_wb_data_i[21]
port 272 nsew signal input
rlabel metal3 s 119200 89224 120000 89344 6 localMemory_wb_data_i[22]
port 273 nsew signal input
rlabel metal3 s 119200 90720 120000 90840 6 localMemory_wb_data_i[23]
port 274 nsew signal input
rlabel metal3 s 119200 91672 120000 91792 6 localMemory_wb_data_i[24]
port 275 nsew signal input
rlabel metal3 s 119200 92624 120000 92744 6 localMemory_wb_data_i[25]
port 276 nsew signal input
rlabel metal3 s 119200 93576 120000 93696 6 localMemory_wb_data_i[26]
port 277 nsew signal input
rlabel metal3 s 119200 94664 120000 94784 6 localMemory_wb_data_i[27]
port 278 nsew signal input
rlabel metal3 s 119200 95616 120000 95736 6 localMemory_wb_data_i[28]
port 279 nsew signal input
rlabel metal3 s 119200 96568 120000 96688 6 localMemory_wb_data_i[29]
port 280 nsew signal input
rlabel metal3 s 119200 58624 120000 58744 6 localMemory_wb_data_i[2]
port 281 nsew signal input
rlabel metal3 s 119200 97520 120000 97640 6 localMemory_wb_data_i[30]
port 282 nsew signal input
rlabel metal3 s 119200 98608 120000 98728 6 localMemory_wb_data_i[31]
port 283 nsew signal input
rlabel metal3 s 119200 60664 120000 60784 6 localMemory_wb_data_i[3]
port 284 nsew signal input
rlabel metal3 s 119200 62568 120000 62688 6 localMemory_wb_data_i[4]
port 285 nsew signal input
rlabel metal3 s 119200 64064 120000 64184 6 localMemory_wb_data_i[5]
port 286 nsew signal input
rlabel metal3 s 119200 65560 120000 65680 6 localMemory_wb_data_i[6]
port 287 nsew signal input
rlabel metal3 s 119200 67056 120000 67176 6 localMemory_wb_data_i[7]
port 288 nsew signal input
rlabel metal3 s 119200 68552 120000 68672 6 localMemory_wb_data_i[8]
port 289 nsew signal input
rlabel metal3 s 119200 70048 120000 70168 6 localMemory_wb_data_i[9]
port 290 nsew signal input
rlabel metal3 s 119200 55224 120000 55344 6 localMemory_wb_data_o[0]
port 291 nsew signal output
rlabel metal3 s 119200 71952 120000 72072 6 localMemory_wb_data_o[10]
port 292 nsew signal output
rlabel metal3 s 119200 73448 120000 73568 6 localMemory_wb_data_o[11]
port 293 nsew signal output
rlabel metal3 s 119200 74944 120000 75064 6 localMemory_wb_data_o[12]
port 294 nsew signal output
rlabel metal3 s 119200 76440 120000 76560 6 localMemory_wb_data_o[13]
port 295 nsew signal output
rlabel metal3 s 119200 77936 120000 78056 6 localMemory_wb_data_o[14]
port 296 nsew signal output
rlabel metal3 s 119200 79296 120000 79416 6 localMemory_wb_data_o[15]
port 297 nsew signal output
rlabel metal3 s 119200 80792 120000 80912 6 localMemory_wb_data_o[16]
port 298 nsew signal output
rlabel metal3 s 119200 82288 120000 82408 6 localMemory_wb_data_o[17]
port 299 nsew signal output
rlabel metal3 s 119200 83784 120000 83904 6 localMemory_wb_data_o[18]
port 300 nsew signal output
rlabel metal3 s 119200 85280 120000 85400 6 localMemory_wb_data_o[19]
port 301 nsew signal output
rlabel metal3 s 119200 57264 120000 57384 6 localMemory_wb_data_o[1]
port 302 nsew signal output
rlabel metal3 s 119200 86776 120000 86896 6 localMemory_wb_data_o[20]
port 303 nsew signal output
rlabel metal3 s 119200 88272 120000 88392 6 localMemory_wb_data_o[21]
port 304 nsew signal output
rlabel metal3 s 119200 89632 120000 89752 6 localMemory_wb_data_o[22]
port 305 nsew signal output
rlabel metal3 s 119200 91128 120000 91248 6 localMemory_wb_data_o[23]
port 306 nsew signal output
rlabel metal3 s 119200 92216 120000 92336 6 localMemory_wb_data_o[24]
port 307 nsew signal output
rlabel metal3 s 119200 93168 120000 93288 6 localMemory_wb_data_o[25]
port 308 nsew signal output
rlabel metal3 s 119200 94120 120000 94240 6 localMemory_wb_data_o[26]
port 309 nsew signal output
rlabel metal3 s 119200 95072 120000 95192 6 localMemory_wb_data_o[27]
port 310 nsew signal output
rlabel metal3 s 119200 96160 120000 96280 6 localMemory_wb_data_o[28]
port 311 nsew signal output
rlabel metal3 s 119200 97112 120000 97232 6 localMemory_wb_data_o[29]
port 312 nsew signal output
rlabel metal3 s 119200 59168 120000 59288 6 localMemory_wb_data_o[2]
port 313 nsew signal output
rlabel metal3 s 119200 98064 120000 98184 6 localMemory_wb_data_o[30]
port 314 nsew signal output
rlabel metal3 s 119200 99016 120000 99136 6 localMemory_wb_data_o[31]
port 315 nsew signal output
rlabel metal3 s 119200 61072 120000 61192 6 localMemory_wb_data_o[3]
port 316 nsew signal output
rlabel metal3 s 119200 63112 120000 63232 6 localMemory_wb_data_o[4]
port 317 nsew signal output
rlabel metal3 s 119200 64608 120000 64728 6 localMemory_wb_data_o[5]
port 318 nsew signal output
rlabel metal3 s 119200 66104 120000 66224 6 localMemory_wb_data_o[6]
port 319 nsew signal output
rlabel metal3 s 119200 67600 120000 67720 6 localMemory_wb_data_o[7]
port 320 nsew signal output
rlabel metal3 s 119200 68960 120000 69080 6 localMemory_wb_data_o[8]
port 321 nsew signal output
rlabel metal3 s 119200 70456 120000 70576 6 localMemory_wb_data_o[9]
port 322 nsew signal output
rlabel metal3 s 119200 52232 120000 52352 6 localMemory_wb_error_o
port 323 nsew signal output
rlabel metal3 s 119200 55768 120000 55888 6 localMemory_wb_sel_i[0]
port 324 nsew signal input
rlabel metal3 s 119200 57672 120000 57792 6 localMemory_wb_sel_i[1]
port 325 nsew signal input
rlabel metal3 s 119200 59712 120000 59832 6 localMemory_wb_sel_i[2]
port 326 nsew signal input
rlabel metal3 s 119200 61616 120000 61736 6 localMemory_wb_sel_i[3]
port 327 nsew signal input
rlabel metal3 s 119200 52776 120000 52896 6 localMemory_wb_stall_o
port 328 nsew signal output
rlabel metal3 s 119200 53320 120000 53440 6 localMemory_wb_stb_i
port 329 nsew signal input
rlabel metal3 s 119200 53728 120000 53848 6 localMemory_wb_we_i
port 330 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 manufacturerID[0]
port 331 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 manufacturerID[10]
port 332 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 manufacturerID[1]
port 333 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 manufacturerID[2]
port 334 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 manufacturerID[3]
port 335 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 manufacturerID[4]
port 336 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 manufacturerID[5]
port 337 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 manufacturerID[6]
port 338 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 manufacturerID[7]
port 339 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 manufacturerID[8]
port 340 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 manufacturerID[9]
port 341 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 partID[0]
port 342 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 partID[10]
port 343 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 partID[11]
port 344 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 partID[12]
port 345 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 partID[13]
port 346 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 partID[14]
port 347 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 partID[15]
port 348 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 partID[1]
port 349 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 partID[2]
port 350 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 partID[3]
port 351 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 partID[4]
port 352 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 partID[5]
port 353 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 partID[6]
port 354 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 partID[7]
port 355 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 partID[8]
port 356 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 partID[9]
port 357 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 probe_errorCode[0]
port 358 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 probe_errorCode[1]
port 359 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 probe_errorCode[2]
port 360 nsew signal output
rlabel metal3 s 0 35232 800 35352 6 probe_errorCode[3]
port 361 nsew signal output
rlabel metal3 s 0 824 800 944 6 probe_isBranch
port 362 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 probe_isCompressed
port 363 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 probe_isLoad
port 364 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 probe_isStore
port 365 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 probe_jtagInstruction[0]
port 366 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 probe_jtagInstruction[1]
port 367 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 probe_jtagInstruction[2]
port 368 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 probe_jtagInstruction[3]
port 369 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 probe_jtagInstruction[4]
port 370 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 probe_opcode[0]
port 371 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 probe_opcode[1]
port 372 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 probe_opcode[2]
port 373 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 probe_opcode[3]
port 374 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 probe_opcode[4]
port 375 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 probe_opcode[5]
port 376 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 probe_opcode[6]
port 377 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 probe_programCounter[0]
port 378 nsew signal output
rlabel metal3 s 0 60800 800 60920 6 probe_programCounter[10]
port 379 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 probe_programCounter[11]
port 380 nsew signal output
rlabel metal3 s 0 64336 800 64456 6 probe_programCounter[12]
port 381 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 probe_programCounter[13]
port 382 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 probe_programCounter[14]
port 383 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 probe_programCounter[15]
port 384 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 probe_programCounter[16]
port 385 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 probe_programCounter[17]
port 386 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 probe_programCounter[18]
port 387 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 probe_programCounter[19]
port 388 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 probe_programCounter[1]
port 389 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 probe_programCounter[20]
port 390 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 probe_programCounter[21]
port 391 nsew signal output
rlabel metal3 s 0 82560 800 82680 6 probe_programCounter[22]
port 392 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 probe_programCounter[23]
port 393 nsew signal output
rlabel metal3 s 0 86232 800 86352 6 probe_programCounter[24]
port 394 nsew signal output
rlabel metal3 s 0 88000 800 88120 6 probe_programCounter[25]
port 395 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 probe_programCounter[26]
port 396 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 probe_programCounter[27]
port 397 nsew signal output
rlabel metal3 s 0 93440 800 93560 6 probe_programCounter[28]
port 398 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 probe_programCounter[29]
port 399 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 probe_programCounter[2]
port 400 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 probe_programCounter[30]
port 401 nsew signal output
rlabel metal3 s 0 98880 800 99000 6 probe_programCounter[31]
port 402 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 probe_programCounter[3]
port 403 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 probe_programCounter[4]
port 404 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 probe_programCounter[5]
port 405 nsew signal output
rlabel metal3 s 0 53456 800 53576 6 probe_programCounter[6]
port 406 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 probe_programCounter[7]
port 407 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 probe_programCounter[8]
port 408 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 probe_programCounter[9]
port 409 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 probe_state[0]
port 410 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 probe_state[1]
port 411 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 probe_takeBranch
port 412 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 413 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 413 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 413 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 413 nsew power input
rlabel metal2 s 106462 0 106518 800 6 versionID[0]
port 414 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 versionID[1]
port 415 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 versionID[2]
port 416 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 versionID[3]
port 417 nsew signal input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 418 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 418 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 418 nsew ground input
rlabel metal4 s 111728 2128 112048 97424 6 vssd1
port 418 nsew ground input
rlabel metal3 s 119200 144 120000 264 6 wb_clk_i
port 419 nsew signal input
rlabel metal3 s 119200 552 120000 672 6 wb_rst_i
port 420 nsew signal input
rlabel metal2 s 2318 99200 2374 100000 6 web0
port 421 nsew signal output
rlabel metal2 s 3330 99200 3386 100000 6 wmask0[0]
port 422 nsew signal output
rlabel metal2 s 4250 99200 4306 100000 6 wmask0[1]
port 423 nsew signal output
rlabel metal2 s 5262 99200 5318 100000 6 wmask0[2]
port 424 nsew signal output
rlabel metal2 s 6182 99200 6238 100000 6 wmask0[3]
port 425 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 28218602
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/finishing/ExperiarCore.magic.gds
string GDS_START 1389434
<< end >>

