VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 800.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 796.000 5.430 800.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 796.000 15.550 800.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 796.000 25.670 800.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 796.000 35.790 800.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 796.000 46.370 800.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 796.000 56.490 800.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 796.000 66.610 800.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 796.000 77.190 800.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.880 400.000 9.480 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 32.680 400.000 33.280 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 167.320 400.000 167.920 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.880 400.000 179.480 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.120 400.000 191.720 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.680 400.000 203.280 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.920 400.000 215.520 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 226.480 400.000 227.080 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.720 400.000 239.320 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.280 400.000 250.880 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 262.520 400.000 263.120 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.080 400.000 274.680 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 48.320 400.000 48.920 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 286.320 400.000 286.920 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.880 400.000 298.480 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 310.120 400.000 310.720 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.680 400.000 322.280 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 345.480 400.000 346.080 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.040 400.000 357.640 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 369.280 400.000 369.880 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.280 400.000 80.880 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.160 400.000 108.760 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.720 400.000 120.320 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.960 400.000 132.560 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 143.520 400.000 144.120 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 155.760 400.000 156.360 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 12.960 400.000 13.560 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.760 400.000 37.360 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 171.400 400.000 172.000 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 182.960 400.000 183.560 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 195.200 400.000 195.800 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.760 400.000 207.360 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.000 400.000 219.600 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 230.560 400.000 231.160 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 242.800 400.000 243.400 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 254.360 400.000 254.960 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 266.600 400.000 267.200 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.160 400.000 278.760 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 52.400 400.000 53.000 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.720 400.000 290.320 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.960 400.000 302.560 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 313.520 400.000 314.120 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.760 400.000 326.360 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 337.320 400.000 337.920 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 349.560 400.000 350.160 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.120 400.000 361.720 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 373.360 400.000 373.960 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.840 400.000 381.440 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.160 400.000 397.760 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 404.640 400.000 405.240 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 84.360 400.000 84.960 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 100.000 400.000 100.600 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.800 400.000 124.400 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 135.360 400.000 135.960 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 147.600 400.000 148.200 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.160 400.000 159.760 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 40.840 400.000 41.440 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 175.480 400.000 176.080 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 400.000 187.640 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 199.280 400.000 199.880 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 223.080 400.000 223.680 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 234.640 400.000 235.240 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.200 400.000 246.800 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 270.000 400.000 270.600 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.240 400.000 282.840 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 56.480 400.000 57.080 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.800 400.000 294.400 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 317.600 400.000 318.200 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.840 400.000 330.440 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 341.400 400.000 342.000 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 353.640 400.000 354.240 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.200 400.000 365.800 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 377.440 400.000 378.040 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 384.920 400.000 385.520 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.080 400.000 393.680 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.120 400.000 72.720 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 401.240 400.000 401.840 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 408.720 400.000 409.320 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.080 400.000 104.680 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.880 400.000 128.480 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 139.440 400.000 140.040 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.680 400.000 152.280 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.240 400.000 163.840 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.040 400.000 17.640 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.920 400.000 45.520 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 60.560 400.000 61.160 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.200 400.000 76.800 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.840 400.000 92.440 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 21.120 400.000 21.720 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 24.520 400.000 25.120 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 28.600 400.000 29.200 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.000 4.000 644.600 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.720 4.000 715.320 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.800 4.000 719.400 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.200 4.000 739.800 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END dout1[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 412.800 400.000 413.400 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 436.600 400.000 437.200 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 571.240 400.000 571.840 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 582.800 400.000 583.400 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 595.040 400.000 595.640 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 606.600 400.000 607.200 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 618.840 400.000 619.440 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 630.400 400.000 631.000 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 642.640 400.000 643.240 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 654.200 400.000 654.800 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 666.440 400.000 667.040 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 678.000 400.000 678.600 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 452.240 400.000 452.840 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 689.560 400.000 690.160 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 701.800 400.000 702.400 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 713.360 400.000 713.960 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 725.600 400.000 726.200 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 467.880 400.000 468.480 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 484.200 400.000 484.800 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 499.840 400.000 500.440 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 512.080 400.000 512.680 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 523.640 400.000 524.240 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 535.200 400.000 535.800 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 547.440 400.000 548.040 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 559.000 400.000 559.600 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 416.880 400.000 417.480 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 440.680 400.000 441.280 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 575.320 400.000 575.920 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 586.880 400.000 587.480 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 599.120 400.000 599.720 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 610.680 400.000 611.280 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 622.920 400.000 623.520 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 634.480 400.000 635.080 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 646.040 400.000 646.640 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 658.280 400.000 658.880 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 669.840 400.000 670.440 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 682.080 400.000 682.680 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 456.320 400.000 456.920 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 693.640 400.000 694.240 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 705.880 400.000 706.480 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 717.440 400.000 718.040 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 729.680 400.000 730.280 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 737.160 400.000 737.760 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 745.320 400.000 745.920 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 753.480 400.000 754.080 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 760.960 400.000 761.560 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 769.120 400.000 769.720 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 777.280 400.000 777.880 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 471.960 400.000 472.560 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 784.760 400.000 785.360 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 792.920 400.000 793.520 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 488.280 400.000 488.880 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 503.920 400.000 504.520 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 515.480 400.000 516.080 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 527.720 400.000 528.320 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 539.280 400.000 539.880 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 551.520 400.000 552.120 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 563.080 400.000 563.680 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 444.760 400.000 445.360 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 578.720 400.000 579.320 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 590.960 400.000 591.560 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 602.520 400.000 603.120 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 614.760 400.000 615.360 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 626.320 400.000 626.920 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 638.560 400.000 639.160 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 650.120 400.000 650.720 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 662.360 400.000 662.960 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 673.920 400.000 674.520 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 686.160 400.000 686.760 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 460.400 400.000 461.000 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 697.720 400.000 698.320 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 709.960 400.000 710.560 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 721.520 400.000 722.120 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 733.760 400.000 734.360 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 741.240 400.000 741.840 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 749.400 400.000 750.000 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 756.880 400.000 757.480 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 765.040 400.000 765.640 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 773.200 400.000 773.800 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 780.680 400.000 781.280 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 476.040 400.000 476.640 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 788.840 400.000 789.440 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 797.000 400.000 797.600 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 491.680 400.000 492.280 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 508.000 400.000 508.600 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 519.560 400.000 520.160 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 531.800 400.000 532.400 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 543.360 400.000 543.960 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 555.600 400.000 556.200 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 567.160 400.000 567.760 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 420.960 400.000 421.560 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 448.160 400.000 448.760 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 464.480 400.000 465.080 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 480.120 400.000 480.720 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 495.760 400.000 496.360 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 424.360 400.000 424.960 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 428.440 400.000 429.040 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 432.520 400.000 433.120 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 796.000 87.310 800.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 796.000 189.890 800.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 796.000 97.430 800.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 796.000 108.010 800.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 796.000 118.130 800.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 796.000 128.250 800.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 796.000 138.830 800.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 796.000 148.950 800.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 796.000 159.070 800.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 796.000 169.190 800.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 796.000 179.770 800.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 796.000 200.010 800.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 796.000 302.590 800.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 796.000 313.170 800.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 796.000 323.290 800.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 796.000 333.410 800.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 796.000 343.990 800.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 796.000 354.110 800.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 796.000 210.590 800.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 796.000 220.710 800.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 796.000 230.830 800.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 796.000 241.410 800.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 796.000 251.530 800.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 796.000 261.650 800.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 796.000 272.230 800.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 796.000 282.350 800.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 796.000 292.470 800.000 ;
    END
  END partID[9]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END probe_errorCode[1]
  PIN probe_errorCode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END probe_errorCode[2]
  PIN probe_errorCode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END probe_errorCode[3]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 796.000 364.230 800.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 796.000 374.810 800.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 796.000 384.930 800.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 796.000 395.050 800.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1.400 400.000 2.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.800 400.000 5.400 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 788.885 ;
      LAYER met1 ;
        RECT 3.290 6.500 396.450 792.160 ;
      LAYER met2 ;
        RECT 3.320 795.720 4.870 797.485 ;
        RECT 5.710 795.720 14.990 797.485 ;
        RECT 15.830 795.720 25.110 797.485 ;
        RECT 25.950 795.720 35.230 797.485 ;
        RECT 36.070 795.720 45.810 797.485 ;
        RECT 46.650 795.720 55.930 797.485 ;
        RECT 56.770 795.720 66.050 797.485 ;
        RECT 66.890 795.720 76.630 797.485 ;
        RECT 77.470 795.720 86.750 797.485 ;
        RECT 87.590 795.720 96.870 797.485 ;
        RECT 97.710 795.720 107.450 797.485 ;
        RECT 108.290 795.720 117.570 797.485 ;
        RECT 118.410 795.720 127.690 797.485 ;
        RECT 128.530 795.720 138.270 797.485 ;
        RECT 139.110 795.720 148.390 797.485 ;
        RECT 149.230 795.720 158.510 797.485 ;
        RECT 159.350 795.720 168.630 797.485 ;
        RECT 169.470 795.720 179.210 797.485 ;
        RECT 180.050 795.720 189.330 797.485 ;
        RECT 190.170 795.720 199.450 797.485 ;
        RECT 200.290 795.720 210.030 797.485 ;
        RECT 210.870 795.720 220.150 797.485 ;
        RECT 220.990 795.720 230.270 797.485 ;
        RECT 231.110 795.720 240.850 797.485 ;
        RECT 241.690 795.720 250.970 797.485 ;
        RECT 251.810 795.720 261.090 797.485 ;
        RECT 261.930 795.720 271.670 797.485 ;
        RECT 272.510 795.720 281.790 797.485 ;
        RECT 282.630 795.720 291.910 797.485 ;
        RECT 292.750 795.720 302.030 797.485 ;
        RECT 302.870 795.720 312.610 797.485 ;
        RECT 313.450 795.720 322.730 797.485 ;
        RECT 323.570 795.720 332.850 797.485 ;
        RECT 333.690 795.720 343.430 797.485 ;
        RECT 344.270 795.720 353.550 797.485 ;
        RECT 354.390 795.720 363.670 797.485 ;
        RECT 364.510 795.720 374.250 797.485 ;
        RECT 375.090 795.720 384.370 797.485 ;
        RECT 385.210 795.720 394.490 797.485 ;
        RECT 395.330 795.720 396.420 797.485 ;
        RECT 3.320 4.280 396.420 795.720 ;
        RECT 3.870 1.515 9.930 4.280 ;
        RECT 10.770 1.515 17.290 4.280 ;
        RECT 18.130 1.515 24.650 4.280 ;
        RECT 25.490 1.515 32.010 4.280 ;
        RECT 32.850 1.515 39.370 4.280 ;
        RECT 40.210 1.515 46.270 4.280 ;
        RECT 47.110 1.515 53.630 4.280 ;
        RECT 54.470 1.515 60.990 4.280 ;
        RECT 61.830 1.515 68.350 4.280 ;
        RECT 69.190 1.515 75.710 4.280 ;
        RECT 76.550 1.515 83.070 4.280 ;
        RECT 83.910 1.515 89.970 4.280 ;
        RECT 90.810 1.515 97.330 4.280 ;
        RECT 98.170 1.515 104.690 4.280 ;
        RECT 105.530 1.515 112.050 4.280 ;
        RECT 112.890 1.515 119.410 4.280 ;
        RECT 120.250 1.515 126.310 4.280 ;
        RECT 127.150 1.515 133.670 4.280 ;
        RECT 134.510 1.515 141.030 4.280 ;
        RECT 141.870 1.515 148.390 4.280 ;
        RECT 149.230 1.515 155.750 4.280 ;
        RECT 156.590 1.515 163.110 4.280 ;
        RECT 163.950 1.515 170.010 4.280 ;
        RECT 170.850 1.515 177.370 4.280 ;
        RECT 178.210 1.515 184.730 4.280 ;
        RECT 185.570 1.515 192.090 4.280 ;
        RECT 192.930 1.515 199.450 4.280 ;
        RECT 200.290 1.515 206.350 4.280 ;
        RECT 207.190 1.515 213.710 4.280 ;
        RECT 214.550 1.515 221.070 4.280 ;
        RECT 221.910 1.515 228.430 4.280 ;
        RECT 229.270 1.515 235.790 4.280 ;
        RECT 236.630 1.515 243.150 4.280 ;
        RECT 243.990 1.515 250.050 4.280 ;
        RECT 250.890 1.515 257.410 4.280 ;
        RECT 258.250 1.515 264.770 4.280 ;
        RECT 265.610 1.515 272.130 4.280 ;
        RECT 272.970 1.515 279.490 4.280 ;
        RECT 280.330 1.515 286.390 4.280 ;
        RECT 287.230 1.515 293.750 4.280 ;
        RECT 294.590 1.515 301.110 4.280 ;
        RECT 301.950 1.515 308.470 4.280 ;
        RECT 309.310 1.515 315.830 4.280 ;
        RECT 316.670 1.515 323.190 4.280 ;
        RECT 324.030 1.515 330.090 4.280 ;
        RECT 330.930 1.515 337.450 4.280 ;
        RECT 338.290 1.515 344.810 4.280 ;
        RECT 345.650 1.515 352.170 4.280 ;
        RECT 353.010 1.515 359.530 4.280 ;
        RECT 360.370 1.515 366.430 4.280 ;
        RECT 367.270 1.515 373.790 4.280 ;
        RECT 374.630 1.515 381.150 4.280 ;
        RECT 381.990 1.515 388.510 4.280 ;
        RECT 389.350 1.515 395.870 4.280 ;
      LAYER met3 ;
        RECT 4.400 796.600 395.600 797.465 ;
        RECT 4.000 793.920 396.000 796.600 ;
        RECT 4.400 792.520 395.600 793.920 ;
        RECT 4.000 789.840 396.000 792.520 ;
        RECT 4.400 788.440 395.600 789.840 ;
        RECT 4.000 785.760 396.000 788.440 ;
        RECT 4.400 784.360 395.600 785.760 ;
        RECT 4.000 781.680 396.000 784.360 ;
        RECT 4.400 780.280 395.600 781.680 ;
        RECT 4.000 778.280 396.000 780.280 ;
        RECT 4.000 777.600 395.600 778.280 ;
        RECT 4.400 776.880 395.600 777.600 ;
        RECT 4.400 776.200 396.000 776.880 ;
        RECT 4.000 774.200 396.000 776.200 ;
        RECT 4.000 773.520 395.600 774.200 ;
        RECT 4.400 772.800 395.600 773.520 ;
        RECT 4.400 772.120 396.000 772.800 ;
        RECT 4.000 770.120 396.000 772.120 ;
        RECT 4.000 769.440 395.600 770.120 ;
        RECT 4.400 768.720 395.600 769.440 ;
        RECT 4.400 768.040 396.000 768.720 ;
        RECT 4.000 766.040 396.000 768.040 ;
        RECT 4.000 765.360 395.600 766.040 ;
        RECT 4.400 764.640 395.600 765.360 ;
        RECT 4.400 763.960 396.000 764.640 ;
        RECT 4.000 761.960 396.000 763.960 ;
        RECT 4.000 761.280 395.600 761.960 ;
        RECT 4.400 760.560 395.600 761.280 ;
        RECT 4.400 759.880 396.000 760.560 ;
        RECT 4.000 757.880 396.000 759.880 ;
        RECT 4.000 756.520 395.600 757.880 ;
        RECT 4.400 756.480 395.600 756.520 ;
        RECT 4.400 755.120 396.000 756.480 ;
        RECT 4.000 754.480 396.000 755.120 ;
        RECT 4.000 753.080 395.600 754.480 ;
        RECT 4.000 752.440 396.000 753.080 ;
        RECT 4.400 751.040 396.000 752.440 ;
        RECT 4.000 750.400 396.000 751.040 ;
        RECT 4.000 749.000 395.600 750.400 ;
        RECT 4.000 748.360 396.000 749.000 ;
        RECT 4.400 746.960 396.000 748.360 ;
        RECT 4.000 746.320 396.000 746.960 ;
        RECT 4.000 744.920 395.600 746.320 ;
        RECT 4.000 744.280 396.000 744.920 ;
        RECT 4.400 742.880 396.000 744.280 ;
        RECT 4.000 742.240 396.000 742.880 ;
        RECT 4.000 740.840 395.600 742.240 ;
        RECT 4.000 740.200 396.000 740.840 ;
        RECT 4.400 738.800 396.000 740.200 ;
        RECT 4.000 738.160 396.000 738.800 ;
        RECT 4.000 736.760 395.600 738.160 ;
        RECT 4.000 736.120 396.000 736.760 ;
        RECT 4.400 734.760 396.000 736.120 ;
        RECT 4.400 734.720 395.600 734.760 ;
        RECT 4.000 733.360 395.600 734.720 ;
        RECT 4.000 732.040 396.000 733.360 ;
        RECT 4.400 730.680 396.000 732.040 ;
        RECT 4.400 730.640 395.600 730.680 ;
        RECT 4.000 729.280 395.600 730.640 ;
        RECT 4.000 727.960 396.000 729.280 ;
        RECT 4.400 726.600 396.000 727.960 ;
        RECT 4.400 726.560 395.600 726.600 ;
        RECT 4.000 725.200 395.600 726.560 ;
        RECT 4.000 723.880 396.000 725.200 ;
        RECT 4.400 722.520 396.000 723.880 ;
        RECT 4.400 722.480 395.600 722.520 ;
        RECT 4.000 721.120 395.600 722.480 ;
        RECT 4.000 719.800 396.000 721.120 ;
        RECT 4.400 718.440 396.000 719.800 ;
        RECT 4.400 718.400 395.600 718.440 ;
        RECT 4.000 717.040 395.600 718.400 ;
        RECT 4.000 715.720 396.000 717.040 ;
        RECT 4.400 714.360 396.000 715.720 ;
        RECT 4.400 714.320 395.600 714.360 ;
        RECT 4.000 712.960 395.600 714.320 ;
        RECT 4.000 710.960 396.000 712.960 ;
        RECT 4.400 709.560 395.600 710.960 ;
        RECT 4.000 706.880 396.000 709.560 ;
        RECT 4.400 705.480 395.600 706.880 ;
        RECT 4.000 702.800 396.000 705.480 ;
        RECT 4.400 701.400 395.600 702.800 ;
        RECT 4.000 698.720 396.000 701.400 ;
        RECT 4.400 697.320 395.600 698.720 ;
        RECT 4.000 694.640 396.000 697.320 ;
        RECT 4.400 693.240 395.600 694.640 ;
        RECT 4.000 690.560 396.000 693.240 ;
        RECT 4.400 689.160 395.600 690.560 ;
        RECT 4.000 687.160 396.000 689.160 ;
        RECT 4.000 686.480 395.600 687.160 ;
        RECT 4.400 685.760 395.600 686.480 ;
        RECT 4.400 685.080 396.000 685.760 ;
        RECT 4.000 683.080 396.000 685.080 ;
        RECT 4.000 682.400 395.600 683.080 ;
        RECT 4.400 681.680 395.600 682.400 ;
        RECT 4.400 681.000 396.000 681.680 ;
        RECT 4.000 679.000 396.000 681.000 ;
        RECT 4.000 678.320 395.600 679.000 ;
        RECT 4.400 677.600 395.600 678.320 ;
        RECT 4.400 676.920 396.000 677.600 ;
        RECT 4.000 674.920 396.000 676.920 ;
        RECT 4.000 674.240 395.600 674.920 ;
        RECT 4.400 673.520 395.600 674.240 ;
        RECT 4.400 672.840 396.000 673.520 ;
        RECT 4.000 670.840 396.000 672.840 ;
        RECT 4.000 670.160 395.600 670.840 ;
        RECT 4.400 669.440 395.600 670.160 ;
        RECT 4.400 668.760 396.000 669.440 ;
        RECT 4.000 667.440 396.000 668.760 ;
        RECT 4.000 666.040 395.600 667.440 ;
        RECT 4.000 665.400 396.000 666.040 ;
        RECT 4.400 664.000 396.000 665.400 ;
        RECT 4.000 663.360 396.000 664.000 ;
        RECT 4.000 661.960 395.600 663.360 ;
        RECT 4.000 661.320 396.000 661.960 ;
        RECT 4.400 659.920 396.000 661.320 ;
        RECT 4.000 659.280 396.000 659.920 ;
        RECT 4.000 657.880 395.600 659.280 ;
        RECT 4.000 657.240 396.000 657.880 ;
        RECT 4.400 655.840 396.000 657.240 ;
        RECT 4.000 655.200 396.000 655.840 ;
        RECT 4.000 653.800 395.600 655.200 ;
        RECT 4.000 653.160 396.000 653.800 ;
        RECT 4.400 651.760 396.000 653.160 ;
        RECT 4.000 651.120 396.000 651.760 ;
        RECT 4.000 649.720 395.600 651.120 ;
        RECT 4.000 649.080 396.000 649.720 ;
        RECT 4.400 647.680 396.000 649.080 ;
        RECT 4.000 647.040 396.000 647.680 ;
        RECT 4.000 645.640 395.600 647.040 ;
        RECT 4.000 645.000 396.000 645.640 ;
        RECT 4.400 643.640 396.000 645.000 ;
        RECT 4.400 643.600 395.600 643.640 ;
        RECT 4.000 642.240 395.600 643.600 ;
        RECT 4.000 640.920 396.000 642.240 ;
        RECT 4.400 639.560 396.000 640.920 ;
        RECT 4.400 639.520 395.600 639.560 ;
        RECT 4.000 638.160 395.600 639.520 ;
        RECT 4.000 636.840 396.000 638.160 ;
        RECT 4.400 635.480 396.000 636.840 ;
        RECT 4.400 635.440 395.600 635.480 ;
        RECT 4.000 634.080 395.600 635.440 ;
        RECT 4.000 632.760 396.000 634.080 ;
        RECT 4.400 631.400 396.000 632.760 ;
        RECT 4.400 631.360 395.600 631.400 ;
        RECT 4.000 630.000 395.600 631.360 ;
        RECT 4.000 628.680 396.000 630.000 ;
        RECT 4.400 627.320 396.000 628.680 ;
        RECT 4.400 627.280 395.600 627.320 ;
        RECT 4.000 625.920 395.600 627.280 ;
        RECT 4.000 623.920 396.000 625.920 ;
        RECT 4.400 622.520 395.600 623.920 ;
        RECT 4.000 619.840 396.000 622.520 ;
        RECT 4.400 618.440 395.600 619.840 ;
        RECT 4.000 615.760 396.000 618.440 ;
        RECT 4.400 614.360 395.600 615.760 ;
        RECT 4.000 611.680 396.000 614.360 ;
        RECT 4.400 610.280 395.600 611.680 ;
        RECT 4.000 607.600 396.000 610.280 ;
        RECT 4.400 606.200 395.600 607.600 ;
        RECT 4.000 603.520 396.000 606.200 ;
        RECT 4.400 602.120 395.600 603.520 ;
        RECT 4.000 600.120 396.000 602.120 ;
        RECT 4.000 599.440 395.600 600.120 ;
        RECT 4.400 598.720 395.600 599.440 ;
        RECT 4.400 598.040 396.000 598.720 ;
        RECT 4.000 596.040 396.000 598.040 ;
        RECT 4.000 595.360 395.600 596.040 ;
        RECT 4.400 594.640 395.600 595.360 ;
        RECT 4.400 593.960 396.000 594.640 ;
        RECT 4.000 591.960 396.000 593.960 ;
        RECT 4.000 591.280 395.600 591.960 ;
        RECT 4.400 590.560 395.600 591.280 ;
        RECT 4.400 589.880 396.000 590.560 ;
        RECT 4.000 587.880 396.000 589.880 ;
        RECT 4.000 587.200 395.600 587.880 ;
        RECT 4.400 586.480 395.600 587.200 ;
        RECT 4.400 585.800 396.000 586.480 ;
        RECT 4.000 583.800 396.000 585.800 ;
        RECT 4.000 583.120 395.600 583.800 ;
        RECT 4.400 582.400 395.600 583.120 ;
        RECT 4.400 581.720 396.000 582.400 ;
        RECT 4.000 579.720 396.000 581.720 ;
        RECT 4.000 578.360 395.600 579.720 ;
        RECT 4.400 578.320 395.600 578.360 ;
        RECT 4.400 576.960 396.000 578.320 ;
        RECT 4.000 576.320 396.000 576.960 ;
        RECT 4.000 574.920 395.600 576.320 ;
        RECT 4.000 574.280 396.000 574.920 ;
        RECT 4.400 572.880 396.000 574.280 ;
        RECT 4.000 572.240 396.000 572.880 ;
        RECT 4.000 570.840 395.600 572.240 ;
        RECT 4.000 570.200 396.000 570.840 ;
        RECT 4.400 568.800 396.000 570.200 ;
        RECT 4.000 568.160 396.000 568.800 ;
        RECT 4.000 566.760 395.600 568.160 ;
        RECT 4.000 566.120 396.000 566.760 ;
        RECT 4.400 564.720 396.000 566.120 ;
        RECT 4.000 564.080 396.000 564.720 ;
        RECT 4.000 562.680 395.600 564.080 ;
        RECT 4.000 562.040 396.000 562.680 ;
        RECT 4.400 560.640 396.000 562.040 ;
        RECT 4.000 560.000 396.000 560.640 ;
        RECT 4.000 558.600 395.600 560.000 ;
        RECT 4.000 557.960 396.000 558.600 ;
        RECT 4.400 556.600 396.000 557.960 ;
        RECT 4.400 556.560 395.600 556.600 ;
        RECT 4.000 555.200 395.600 556.560 ;
        RECT 4.000 553.880 396.000 555.200 ;
        RECT 4.400 552.520 396.000 553.880 ;
        RECT 4.400 552.480 395.600 552.520 ;
        RECT 4.000 551.120 395.600 552.480 ;
        RECT 4.000 549.800 396.000 551.120 ;
        RECT 4.400 548.440 396.000 549.800 ;
        RECT 4.400 548.400 395.600 548.440 ;
        RECT 4.000 547.040 395.600 548.400 ;
        RECT 4.000 545.720 396.000 547.040 ;
        RECT 4.400 544.360 396.000 545.720 ;
        RECT 4.400 544.320 395.600 544.360 ;
        RECT 4.000 542.960 395.600 544.320 ;
        RECT 4.000 541.640 396.000 542.960 ;
        RECT 4.400 540.280 396.000 541.640 ;
        RECT 4.400 540.240 395.600 540.280 ;
        RECT 4.000 538.880 395.600 540.240 ;
        RECT 4.000 537.560 396.000 538.880 ;
        RECT 4.400 536.200 396.000 537.560 ;
        RECT 4.400 536.160 395.600 536.200 ;
        RECT 4.000 534.800 395.600 536.160 ;
        RECT 4.000 532.800 396.000 534.800 ;
        RECT 4.400 531.400 395.600 532.800 ;
        RECT 4.000 528.720 396.000 531.400 ;
        RECT 4.400 527.320 395.600 528.720 ;
        RECT 4.000 524.640 396.000 527.320 ;
        RECT 4.400 523.240 395.600 524.640 ;
        RECT 4.000 520.560 396.000 523.240 ;
        RECT 4.400 519.160 395.600 520.560 ;
        RECT 4.000 516.480 396.000 519.160 ;
        RECT 4.400 515.080 395.600 516.480 ;
        RECT 4.000 513.080 396.000 515.080 ;
        RECT 4.000 512.400 395.600 513.080 ;
        RECT 4.400 511.680 395.600 512.400 ;
        RECT 4.400 511.000 396.000 511.680 ;
        RECT 4.000 509.000 396.000 511.000 ;
        RECT 4.000 508.320 395.600 509.000 ;
        RECT 4.400 507.600 395.600 508.320 ;
        RECT 4.400 506.920 396.000 507.600 ;
        RECT 4.000 504.920 396.000 506.920 ;
        RECT 4.000 504.240 395.600 504.920 ;
        RECT 4.400 503.520 395.600 504.240 ;
        RECT 4.400 502.840 396.000 503.520 ;
        RECT 4.000 500.840 396.000 502.840 ;
        RECT 4.000 500.160 395.600 500.840 ;
        RECT 4.400 499.440 395.600 500.160 ;
        RECT 4.400 498.760 396.000 499.440 ;
        RECT 4.000 496.760 396.000 498.760 ;
        RECT 4.000 496.080 395.600 496.760 ;
        RECT 4.400 495.360 395.600 496.080 ;
        RECT 4.400 494.680 396.000 495.360 ;
        RECT 4.000 492.680 396.000 494.680 ;
        RECT 4.000 492.000 395.600 492.680 ;
        RECT 4.400 491.280 395.600 492.000 ;
        RECT 4.400 490.600 396.000 491.280 ;
        RECT 4.000 489.280 396.000 490.600 ;
        RECT 4.000 487.880 395.600 489.280 ;
        RECT 4.000 487.240 396.000 487.880 ;
        RECT 4.400 485.840 396.000 487.240 ;
        RECT 4.000 485.200 396.000 485.840 ;
        RECT 4.000 483.800 395.600 485.200 ;
        RECT 4.000 483.160 396.000 483.800 ;
        RECT 4.400 481.760 396.000 483.160 ;
        RECT 4.000 481.120 396.000 481.760 ;
        RECT 4.000 479.720 395.600 481.120 ;
        RECT 4.000 479.080 396.000 479.720 ;
        RECT 4.400 477.680 396.000 479.080 ;
        RECT 4.000 477.040 396.000 477.680 ;
        RECT 4.000 475.640 395.600 477.040 ;
        RECT 4.000 475.000 396.000 475.640 ;
        RECT 4.400 473.600 396.000 475.000 ;
        RECT 4.000 472.960 396.000 473.600 ;
        RECT 4.000 471.560 395.600 472.960 ;
        RECT 4.000 470.920 396.000 471.560 ;
        RECT 4.400 469.520 396.000 470.920 ;
        RECT 4.000 468.880 396.000 469.520 ;
        RECT 4.000 467.480 395.600 468.880 ;
        RECT 4.000 466.840 396.000 467.480 ;
        RECT 4.400 465.480 396.000 466.840 ;
        RECT 4.400 465.440 395.600 465.480 ;
        RECT 4.000 464.080 395.600 465.440 ;
        RECT 4.000 462.760 396.000 464.080 ;
        RECT 4.400 461.400 396.000 462.760 ;
        RECT 4.400 461.360 395.600 461.400 ;
        RECT 4.000 460.000 395.600 461.360 ;
        RECT 4.000 458.680 396.000 460.000 ;
        RECT 4.400 457.320 396.000 458.680 ;
        RECT 4.400 457.280 395.600 457.320 ;
        RECT 4.000 455.920 395.600 457.280 ;
        RECT 4.000 454.600 396.000 455.920 ;
        RECT 4.400 453.240 396.000 454.600 ;
        RECT 4.400 453.200 395.600 453.240 ;
        RECT 4.000 451.840 395.600 453.200 ;
        RECT 4.000 450.520 396.000 451.840 ;
        RECT 4.400 449.160 396.000 450.520 ;
        RECT 4.400 449.120 395.600 449.160 ;
        RECT 4.000 447.760 395.600 449.120 ;
        RECT 4.000 445.760 396.000 447.760 ;
        RECT 4.400 444.360 395.600 445.760 ;
        RECT 4.000 441.680 396.000 444.360 ;
        RECT 4.400 440.280 395.600 441.680 ;
        RECT 4.000 437.600 396.000 440.280 ;
        RECT 4.400 436.200 395.600 437.600 ;
        RECT 4.000 433.520 396.000 436.200 ;
        RECT 4.400 432.120 395.600 433.520 ;
        RECT 4.000 429.440 396.000 432.120 ;
        RECT 4.400 428.040 395.600 429.440 ;
        RECT 4.000 425.360 396.000 428.040 ;
        RECT 4.400 423.960 395.600 425.360 ;
        RECT 4.000 421.960 396.000 423.960 ;
        RECT 4.000 421.280 395.600 421.960 ;
        RECT 4.400 420.560 395.600 421.280 ;
        RECT 4.400 419.880 396.000 420.560 ;
        RECT 4.000 417.880 396.000 419.880 ;
        RECT 4.000 417.200 395.600 417.880 ;
        RECT 4.400 416.480 395.600 417.200 ;
        RECT 4.400 415.800 396.000 416.480 ;
        RECT 4.000 413.800 396.000 415.800 ;
        RECT 4.000 413.120 395.600 413.800 ;
        RECT 4.400 412.400 395.600 413.120 ;
        RECT 4.400 411.720 396.000 412.400 ;
        RECT 4.000 409.720 396.000 411.720 ;
        RECT 4.000 409.040 395.600 409.720 ;
        RECT 4.400 408.320 395.600 409.040 ;
        RECT 4.400 407.640 396.000 408.320 ;
        RECT 4.000 405.640 396.000 407.640 ;
        RECT 4.000 404.960 395.600 405.640 ;
        RECT 4.400 404.240 395.600 404.960 ;
        RECT 4.400 403.560 396.000 404.240 ;
        RECT 4.000 402.240 396.000 403.560 ;
        RECT 4.000 400.840 395.600 402.240 ;
        RECT 4.000 400.200 396.000 400.840 ;
        RECT 4.400 398.800 396.000 400.200 ;
        RECT 4.000 398.160 396.000 398.800 ;
        RECT 4.000 396.760 395.600 398.160 ;
        RECT 4.000 396.120 396.000 396.760 ;
        RECT 4.400 394.720 396.000 396.120 ;
        RECT 4.000 394.080 396.000 394.720 ;
        RECT 4.000 392.680 395.600 394.080 ;
        RECT 4.000 392.040 396.000 392.680 ;
        RECT 4.400 390.640 396.000 392.040 ;
        RECT 4.000 390.000 396.000 390.640 ;
        RECT 4.000 388.600 395.600 390.000 ;
        RECT 4.000 387.960 396.000 388.600 ;
        RECT 4.400 386.560 396.000 387.960 ;
        RECT 4.000 385.920 396.000 386.560 ;
        RECT 4.000 384.520 395.600 385.920 ;
        RECT 4.000 383.880 396.000 384.520 ;
        RECT 4.400 382.480 396.000 383.880 ;
        RECT 4.000 381.840 396.000 382.480 ;
        RECT 4.000 380.440 395.600 381.840 ;
        RECT 4.000 379.800 396.000 380.440 ;
        RECT 4.400 378.440 396.000 379.800 ;
        RECT 4.400 378.400 395.600 378.440 ;
        RECT 4.000 377.040 395.600 378.400 ;
        RECT 4.000 375.720 396.000 377.040 ;
        RECT 4.400 374.360 396.000 375.720 ;
        RECT 4.400 374.320 395.600 374.360 ;
        RECT 4.000 372.960 395.600 374.320 ;
        RECT 4.000 371.640 396.000 372.960 ;
        RECT 4.400 370.280 396.000 371.640 ;
        RECT 4.400 370.240 395.600 370.280 ;
        RECT 4.000 368.880 395.600 370.240 ;
        RECT 4.000 367.560 396.000 368.880 ;
        RECT 4.400 366.200 396.000 367.560 ;
        RECT 4.400 366.160 395.600 366.200 ;
        RECT 4.000 364.800 395.600 366.160 ;
        RECT 4.000 363.480 396.000 364.800 ;
        RECT 4.400 362.120 396.000 363.480 ;
        RECT 4.400 362.080 395.600 362.120 ;
        RECT 4.000 360.720 395.600 362.080 ;
        RECT 4.000 359.400 396.000 360.720 ;
        RECT 4.400 358.040 396.000 359.400 ;
        RECT 4.400 358.000 395.600 358.040 ;
        RECT 4.000 356.640 395.600 358.000 ;
        RECT 4.000 354.640 396.000 356.640 ;
        RECT 4.400 353.240 395.600 354.640 ;
        RECT 4.000 350.560 396.000 353.240 ;
        RECT 4.400 349.160 395.600 350.560 ;
        RECT 4.000 346.480 396.000 349.160 ;
        RECT 4.400 345.080 395.600 346.480 ;
        RECT 4.000 342.400 396.000 345.080 ;
        RECT 4.400 341.000 395.600 342.400 ;
        RECT 4.000 338.320 396.000 341.000 ;
        RECT 4.400 336.920 395.600 338.320 ;
        RECT 4.000 334.920 396.000 336.920 ;
        RECT 4.000 334.240 395.600 334.920 ;
        RECT 4.400 333.520 395.600 334.240 ;
        RECT 4.400 332.840 396.000 333.520 ;
        RECT 4.000 330.840 396.000 332.840 ;
        RECT 4.000 330.160 395.600 330.840 ;
        RECT 4.400 329.440 395.600 330.160 ;
        RECT 4.400 328.760 396.000 329.440 ;
        RECT 4.000 326.760 396.000 328.760 ;
        RECT 4.000 326.080 395.600 326.760 ;
        RECT 4.400 325.360 395.600 326.080 ;
        RECT 4.400 324.680 396.000 325.360 ;
        RECT 4.000 322.680 396.000 324.680 ;
        RECT 4.000 322.000 395.600 322.680 ;
        RECT 4.400 321.280 395.600 322.000 ;
        RECT 4.400 320.600 396.000 321.280 ;
        RECT 4.000 318.600 396.000 320.600 ;
        RECT 4.000 317.920 395.600 318.600 ;
        RECT 4.400 317.200 395.600 317.920 ;
        RECT 4.400 316.520 396.000 317.200 ;
        RECT 4.000 314.520 396.000 316.520 ;
        RECT 4.000 313.160 395.600 314.520 ;
        RECT 4.400 313.120 395.600 313.160 ;
        RECT 4.400 311.760 396.000 313.120 ;
        RECT 4.000 311.120 396.000 311.760 ;
        RECT 4.000 309.720 395.600 311.120 ;
        RECT 4.000 309.080 396.000 309.720 ;
        RECT 4.400 307.680 396.000 309.080 ;
        RECT 4.000 307.040 396.000 307.680 ;
        RECT 4.000 305.640 395.600 307.040 ;
        RECT 4.000 305.000 396.000 305.640 ;
        RECT 4.400 303.600 396.000 305.000 ;
        RECT 4.000 302.960 396.000 303.600 ;
        RECT 4.000 301.560 395.600 302.960 ;
        RECT 4.000 300.920 396.000 301.560 ;
        RECT 4.400 299.520 396.000 300.920 ;
        RECT 4.000 298.880 396.000 299.520 ;
        RECT 4.000 297.480 395.600 298.880 ;
        RECT 4.000 296.840 396.000 297.480 ;
        RECT 4.400 295.440 396.000 296.840 ;
        RECT 4.000 294.800 396.000 295.440 ;
        RECT 4.000 293.400 395.600 294.800 ;
        RECT 4.000 292.760 396.000 293.400 ;
        RECT 4.400 291.360 396.000 292.760 ;
        RECT 4.000 290.720 396.000 291.360 ;
        RECT 4.000 289.320 395.600 290.720 ;
        RECT 4.000 288.680 396.000 289.320 ;
        RECT 4.400 287.320 396.000 288.680 ;
        RECT 4.400 287.280 395.600 287.320 ;
        RECT 4.000 285.920 395.600 287.280 ;
        RECT 4.000 284.600 396.000 285.920 ;
        RECT 4.400 283.240 396.000 284.600 ;
        RECT 4.400 283.200 395.600 283.240 ;
        RECT 4.000 281.840 395.600 283.200 ;
        RECT 4.000 280.520 396.000 281.840 ;
        RECT 4.400 279.160 396.000 280.520 ;
        RECT 4.400 279.120 395.600 279.160 ;
        RECT 4.000 277.760 395.600 279.120 ;
        RECT 4.000 276.440 396.000 277.760 ;
        RECT 4.400 275.080 396.000 276.440 ;
        RECT 4.400 275.040 395.600 275.080 ;
        RECT 4.000 273.680 395.600 275.040 ;
        RECT 4.000 272.360 396.000 273.680 ;
        RECT 4.400 271.000 396.000 272.360 ;
        RECT 4.400 270.960 395.600 271.000 ;
        RECT 4.000 269.600 395.600 270.960 ;
        RECT 4.000 267.600 396.000 269.600 ;
        RECT 4.400 266.200 395.600 267.600 ;
        RECT 4.000 263.520 396.000 266.200 ;
        RECT 4.400 262.120 395.600 263.520 ;
        RECT 4.000 259.440 396.000 262.120 ;
        RECT 4.400 258.040 395.600 259.440 ;
        RECT 4.000 255.360 396.000 258.040 ;
        RECT 4.400 253.960 395.600 255.360 ;
        RECT 4.000 251.280 396.000 253.960 ;
        RECT 4.400 249.880 395.600 251.280 ;
        RECT 4.000 247.200 396.000 249.880 ;
        RECT 4.400 245.800 395.600 247.200 ;
        RECT 4.000 243.800 396.000 245.800 ;
        RECT 4.000 243.120 395.600 243.800 ;
        RECT 4.400 242.400 395.600 243.120 ;
        RECT 4.400 241.720 396.000 242.400 ;
        RECT 4.000 239.720 396.000 241.720 ;
        RECT 4.000 239.040 395.600 239.720 ;
        RECT 4.400 238.320 395.600 239.040 ;
        RECT 4.400 237.640 396.000 238.320 ;
        RECT 4.000 235.640 396.000 237.640 ;
        RECT 4.000 234.960 395.600 235.640 ;
        RECT 4.400 234.240 395.600 234.960 ;
        RECT 4.400 233.560 396.000 234.240 ;
        RECT 4.000 231.560 396.000 233.560 ;
        RECT 4.000 230.880 395.600 231.560 ;
        RECT 4.400 230.160 395.600 230.880 ;
        RECT 4.400 229.480 396.000 230.160 ;
        RECT 4.000 227.480 396.000 229.480 ;
        RECT 4.000 226.800 395.600 227.480 ;
        RECT 4.400 226.080 395.600 226.800 ;
        RECT 4.400 225.400 396.000 226.080 ;
        RECT 4.000 224.080 396.000 225.400 ;
        RECT 4.000 222.680 395.600 224.080 ;
        RECT 4.000 222.040 396.000 222.680 ;
        RECT 4.400 220.640 396.000 222.040 ;
        RECT 4.000 220.000 396.000 220.640 ;
        RECT 4.000 218.600 395.600 220.000 ;
        RECT 4.000 217.960 396.000 218.600 ;
        RECT 4.400 216.560 396.000 217.960 ;
        RECT 4.000 215.920 396.000 216.560 ;
        RECT 4.000 214.520 395.600 215.920 ;
        RECT 4.000 213.880 396.000 214.520 ;
        RECT 4.400 212.480 396.000 213.880 ;
        RECT 4.000 211.840 396.000 212.480 ;
        RECT 4.000 210.440 395.600 211.840 ;
        RECT 4.000 209.800 396.000 210.440 ;
        RECT 4.400 208.400 396.000 209.800 ;
        RECT 4.000 207.760 396.000 208.400 ;
        RECT 4.000 206.360 395.600 207.760 ;
        RECT 4.000 205.720 396.000 206.360 ;
        RECT 4.400 204.320 396.000 205.720 ;
        RECT 4.000 203.680 396.000 204.320 ;
        RECT 4.000 202.280 395.600 203.680 ;
        RECT 4.000 201.640 396.000 202.280 ;
        RECT 4.400 200.280 396.000 201.640 ;
        RECT 4.400 200.240 395.600 200.280 ;
        RECT 4.000 198.880 395.600 200.240 ;
        RECT 4.000 197.560 396.000 198.880 ;
        RECT 4.400 196.200 396.000 197.560 ;
        RECT 4.400 196.160 395.600 196.200 ;
        RECT 4.000 194.800 395.600 196.160 ;
        RECT 4.000 193.480 396.000 194.800 ;
        RECT 4.400 192.120 396.000 193.480 ;
        RECT 4.400 192.080 395.600 192.120 ;
        RECT 4.000 190.720 395.600 192.080 ;
        RECT 4.000 189.400 396.000 190.720 ;
        RECT 4.400 188.040 396.000 189.400 ;
        RECT 4.400 188.000 395.600 188.040 ;
        RECT 4.000 186.640 395.600 188.000 ;
        RECT 4.000 185.320 396.000 186.640 ;
        RECT 4.400 183.960 396.000 185.320 ;
        RECT 4.400 183.920 395.600 183.960 ;
        RECT 4.000 182.560 395.600 183.920 ;
        RECT 4.000 181.240 396.000 182.560 ;
        RECT 4.400 179.880 396.000 181.240 ;
        RECT 4.400 179.840 395.600 179.880 ;
        RECT 4.000 178.480 395.600 179.840 ;
        RECT 4.000 176.480 396.000 178.480 ;
        RECT 4.400 175.080 395.600 176.480 ;
        RECT 4.000 172.400 396.000 175.080 ;
        RECT 4.400 171.000 395.600 172.400 ;
        RECT 4.000 168.320 396.000 171.000 ;
        RECT 4.400 166.920 395.600 168.320 ;
        RECT 4.000 164.240 396.000 166.920 ;
        RECT 4.400 162.840 395.600 164.240 ;
        RECT 4.000 160.160 396.000 162.840 ;
        RECT 4.400 158.760 395.600 160.160 ;
        RECT 4.000 156.760 396.000 158.760 ;
        RECT 4.000 156.080 395.600 156.760 ;
        RECT 4.400 155.360 395.600 156.080 ;
        RECT 4.400 154.680 396.000 155.360 ;
        RECT 4.000 152.680 396.000 154.680 ;
        RECT 4.000 152.000 395.600 152.680 ;
        RECT 4.400 151.280 395.600 152.000 ;
        RECT 4.400 150.600 396.000 151.280 ;
        RECT 4.000 148.600 396.000 150.600 ;
        RECT 4.000 147.920 395.600 148.600 ;
        RECT 4.400 147.200 395.600 147.920 ;
        RECT 4.400 146.520 396.000 147.200 ;
        RECT 4.000 144.520 396.000 146.520 ;
        RECT 4.000 143.840 395.600 144.520 ;
        RECT 4.400 143.120 395.600 143.840 ;
        RECT 4.400 142.440 396.000 143.120 ;
        RECT 4.000 140.440 396.000 142.440 ;
        RECT 4.000 139.760 395.600 140.440 ;
        RECT 4.400 139.040 395.600 139.760 ;
        RECT 4.400 138.360 396.000 139.040 ;
        RECT 4.000 136.360 396.000 138.360 ;
        RECT 4.000 135.000 395.600 136.360 ;
        RECT 4.400 134.960 395.600 135.000 ;
        RECT 4.400 133.600 396.000 134.960 ;
        RECT 4.000 132.960 396.000 133.600 ;
        RECT 4.000 131.560 395.600 132.960 ;
        RECT 4.000 130.920 396.000 131.560 ;
        RECT 4.400 129.520 396.000 130.920 ;
        RECT 4.000 128.880 396.000 129.520 ;
        RECT 4.000 127.480 395.600 128.880 ;
        RECT 4.000 126.840 396.000 127.480 ;
        RECT 4.400 125.440 396.000 126.840 ;
        RECT 4.000 124.800 396.000 125.440 ;
        RECT 4.000 123.400 395.600 124.800 ;
        RECT 4.000 122.760 396.000 123.400 ;
        RECT 4.400 121.360 396.000 122.760 ;
        RECT 4.000 120.720 396.000 121.360 ;
        RECT 4.000 119.320 395.600 120.720 ;
        RECT 4.000 118.680 396.000 119.320 ;
        RECT 4.400 117.280 396.000 118.680 ;
        RECT 4.000 116.640 396.000 117.280 ;
        RECT 4.000 115.240 395.600 116.640 ;
        RECT 4.000 114.600 396.000 115.240 ;
        RECT 4.400 113.240 396.000 114.600 ;
        RECT 4.400 113.200 395.600 113.240 ;
        RECT 4.000 111.840 395.600 113.200 ;
        RECT 4.000 110.520 396.000 111.840 ;
        RECT 4.400 109.160 396.000 110.520 ;
        RECT 4.400 109.120 395.600 109.160 ;
        RECT 4.000 107.760 395.600 109.120 ;
        RECT 4.000 106.440 396.000 107.760 ;
        RECT 4.400 105.080 396.000 106.440 ;
        RECT 4.400 105.040 395.600 105.080 ;
        RECT 4.000 103.680 395.600 105.040 ;
        RECT 4.000 102.360 396.000 103.680 ;
        RECT 4.400 101.000 396.000 102.360 ;
        RECT 4.400 100.960 395.600 101.000 ;
        RECT 4.000 99.600 395.600 100.960 ;
        RECT 4.000 98.280 396.000 99.600 ;
        RECT 4.400 96.920 396.000 98.280 ;
        RECT 4.400 96.880 395.600 96.920 ;
        RECT 4.000 95.520 395.600 96.880 ;
        RECT 4.000 94.200 396.000 95.520 ;
        RECT 4.400 92.840 396.000 94.200 ;
        RECT 4.400 92.800 395.600 92.840 ;
        RECT 4.000 91.440 395.600 92.800 ;
        RECT 4.000 89.440 396.000 91.440 ;
        RECT 4.400 88.040 395.600 89.440 ;
        RECT 4.000 85.360 396.000 88.040 ;
        RECT 4.400 83.960 395.600 85.360 ;
        RECT 4.000 81.280 396.000 83.960 ;
        RECT 4.400 79.880 395.600 81.280 ;
        RECT 4.000 77.200 396.000 79.880 ;
        RECT 4.400 75.800 395.600 77.200 ;
        RECT 4.000 73.120 396.000 75.800 ;
        RECT 4.400 71.720 395.600 73.120 ;
        RECT 4.000 69.040 396.000 71.720 ;
        RECT 4.400 67.640 395.600 69.040 ;
        RECT 4.000 65.640 396.000 67.640 ;
        RECT 4.000 64.960 395.600 65.640 ;
        RECT 4.400 64.240 395.600 64.960 ;
        RECT 4.400 63.560 396.000 64.240 ;
        RECT 4.000 61.560 396.000 63.560 ;
        RECT 4.000 60.880 395.600 61.560 ;
        RECT 4.400 60.160 395.600 60.880 ;
        RECT 4.400 59.480 396.000 60.160 ;
        RECT 4.000 57.480 396.000 59.480 ;
        RECT 4.000 56.800 395.600 57.480 ;
        RECT 4.400 56.080 395.600 56.800 ;
        RECT 4.400 55.400 396.000 56.080 ;
        RECT 4.000 53.400 396.000 55.400 ;
        RECT 4.000 52.720 395.600 53.400 ;
        RECT 4.400 52.000 395.600 52.720 ;
        RECT 4.400 51.320 396.000 52.000 ;
        RECT 4.000 49.320 396.000 51.320 ;
        RECT 4.000 48.640 395.600 49.320 ;
        RECT 4.400 47.920 395.600 48.640 ;
        RECT 4.400 47.240 396.000 47.920 ;
        RECT 4.000 45.920 396.000 47.240 ;
        RECT 4.000 44.520 395.600 45.920 ;
        RECT 4.000 43.880 396.000 44.520 ;
        RECT 4.400 42.480 396.000 43.880 ;
        RECT 4.000 41.840 396.000 42.480 ;
        RECT 4.000 40.440 395.600 41.840 ;
        RECT 4.000 39.800 396.000 40.440 ;
        RECT 4.400 38.400 396.000 39.800 ;
        RECT 4.000 37.760 396.000 38.400 ;
        RECT 4.000 36.360 395.600 37.760 ;
        RECT 4.000 35.720 396.000 36.360 ;
        RECT 4.400 34.320 396.000 35.720 ;
        RECT 4.000 33.680 396.000 34.320 ;
        RECT 4.000 32.280 395.600 33.680 ;
        RECT 4.000 31.640 396.000 32.280 ;
        RECT 4.400 30.240 396.000 31.640 ;
        RECT 4.000 29.600 396.000 30.240 ;
        RECT 4.000 28.200 395.600 29.600 ;
        RECT 4.000 27.560 396.000 28.200 ;
        RECT 4.400 26.160 396.000 27.560 ;
        RECT 4.000 25.520 396.000 26.160 ;
        RECT 4.000 24.120 395.600 25.520 ;
        RECT 4.000 23.480 396.000 24.120 ;
        RECT 4.400 22.120 396.000 23.480 ;
        RECT 4.400 22.080 395.600 22.120 ;
        RECT 4.000 20.720 395.600 22.080 ;
        RECT 4.000 19.400 396.000 20.720 ;
        RECT 4.400 18.040 396.000 19.400 ;
        RECT 4.400 18.000 395.600 18.040 ;
        RECT 4.000 16.640 395.600 18.000 ;
        RECT 4.000 15.320 396.000 16.640 ;
        RECT 4.400 13.960 396.000 15.320 ;
        RECT 4.400 13.920 395.600 13.960 ;
        RECT 4.000 12.560 395.600 13.920 ;
        RECT 4.000 11.240 396.000 12.560 ;
        RECT 4.400 9.880 396.000 11.240 ;
        RECT 4.400 9.840 395.600 9.880 ;
        RECT 4.000 8.480 395.600 9.840 ;
        RECT 4.000 7.160 396.000 8.480 ;
        RECT 4.400 5.800 396.000 7.160 ;
        RECT 4.400 5.760 395.600 5.800 ;
        RECT 4.000 4.400 395.600 5.760 ;
        RECT 4.000 3.080 396.000 4.400 ;
        RECT 4.400 2.400 396.000 3.080 ;
        RECT 4.400 1.680 395.600 2.400 ;
        RECT 4.000 1.535 395.600 1.680 ;
      LAYER met4 ;
        RECT 176.935 553.695 177.265 623.385 ;
  END
END ExperiarCore
END LIBRARY

