* NGSPICE file created from Peripherals.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt Peripherals flash_csb flash_io0_read flash_io0_we flash_io0_write flash_io1_read
+ flash_io1_we flash_io1_write flash_sck internal_uart_rx internal_uart_tx io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms probe_blink[0] probe_blink[1] vccd1 vga_b[0] vga_b[1] vga_g[0] vga_g[1]
+ vga_hsync vga_r[0] vga_r[1] vga_vsync vssd1 wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11]
+ wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18]
+ wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[2]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_data_i[0] wb_data_i[10] wb_data_i[11] wb_data_i[12] wb_data_i[13]
+ wb_data_i[14] wb_data_i[15] wb_data_i[16] wb_data_i[17] wb_data_i[18] wb_data_i[19]
+ wb_data_i[1] wb_data_i[20] wb_data_i[21] wb_data_i[22] wb_data_i[23] wb_data_i[24]
+ wb_data_i[25] wb_data_i[26] wb_data_i[27] wb_data_i[28] wb_data_i[29] wb_data_i[2]
+ wb_data_i[30] wb_data_i[31] wb_data_i[3] wb_data_i[4] wb_data_i[5] wb_data_i[6]
+ wb_data_i[7] wb_data_i[8] wb_data_i[9] wb_data_o[0] wb_data_o[10] wb_data_o[11]
+ wb_data_o[12] wb_data_o[13] wb_data_o[14] wb_data_o[15] wb_data_o[16] wb_data_o[17]
+ wb_data_o[18] wb_data_o[19] wb_data_o[1] wb_data_o[20] wb_data_o[21] wb_data_o[22]
+ wb_data_o[23] wb_data_o[24] wb_data_o[25] wb_data_o[26] wb_data_o[27] wb_data_o[28]
+ wb_data_o[29] wb_data_o[2] wb_data_o[30] wb_data_o[31] wb_data_o[3] wb_data_o[4]
+ wb_data_o[5] wb_data_o[6] wb_data_o[7] wb_data_o[8] wb_data_o[9] wb_error_o wb_rst_i
+ wb_sel_i[0] wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stall_o wb_stb_i wb_we_i
XFILLER_246_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09671_ _09671_/A vssd1 vssd1 vccd1 vccd1 _18907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18869_ _18869_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15756__1040 _15758__1042/A vssd1 vssd1 vccd1 vccd1 _18757_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09105_ _19191_/Q _09104_/X _09105_/S vssd1 vssd1 vccd1 vccd1 _09106_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09036_ _09035_/X _19209_/Q _09044_/S vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15122__838 _15122__838/A vssd1 vssd1 vccd1 vccd1 _18514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ _10274_/A _10620_/A vssd1 vssd1 vccd1 vccd1 _09968_/S sky130_fd_sc_hd__nor2_2
XFILLER_237_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09869_ _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09874_/A sky130_fd_sc_hd__and2_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11900_ _19250_/Q _19251_/Q _11956_/S vssd1 vssd1 vccd1 vccd1 _11900_/X sky130_fd_sc_hd__mux2_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12880_ _12877_/X _12880_/B vssd1 vssd1 vccd1 vccd1 _12881_/A sky130_fd_sc_hd__and2b_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11831_ _17722_/Q input18/X _11831_/C vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__and3b_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14550_ _14572_/A vssd1 vssd1 vccd1 vccd1 _14729_/S sky130_fd_sc_hd__buf_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11762_ _17864_/Q _17686_/Q _18001_/Q vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ _13281_/X _13500_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _13501_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10713_ _10713_/A vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__buf_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14481_ _14487_/A vssd1 vssd1 vccd1 vccd1 _14481_/X sky130_fd_sc_hd__buf_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11693_ _19040_/Q _18411_/Q _16620_/B vssd1 vssd1 vccd1 vccd1 _11694_/C sky130_fd_sc_hd__and3_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ _18597_/Q _18613_/Q _18739_/Q _18520_/Q _16195_/X _16138_/X vssd1 vssd1 vccd1
+ vccd1 _16221_/B sky130_fd_sc_hd__mux4_1
XFILLER_224_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13432_ _13430_/Y _13493_/A _13432_/S vssd1 vssd1 vccd1 vccd1 _13433_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10644_ _09265_/X _18434_/Q _10648_/S vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _18712_/Q _18720_/Q _18728_/Q _18493_/Q _16149_/X _16150_/X vssd1 vssd1 vccd1
+ vccd1 _16151_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13400_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _13363_/Y sky130_fd_sc_hd__nor2_1
X_10575_ _10575_/A vssd1 vssd1 vccd1 vccd1 _18495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12314_ _17548_/Q _12180_/X _12298_/X _17562_/Q _12313_/X vssd1 vssd1 vccd1 vccd1
+ _12315_/B sky130_fd_sc_hd__a221o_1
X_13294_ _13237_/X _13288_/X _13293_/X vssd1 vssd1 vccd1 vccd1 _13294_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15033_ _18465_/Q _14967_/X _15032_/Y _15026_/X vssd1 vssd1 vccd1 vccd1 _15034_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03410_ clkbuf_0__03410_/X vssd1 vssd1 vccd1 vccd1 _14818__747/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12176_ _17530_/Q _18030_/Q _12176_/S vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11127_ _11127_/A vssd1 vssd1 vccd1 vccd1 _18226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16984_ _16984_/A _16984_/B vssd1 vssd1 vccd1 vccd1 _16984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18723_ _18723_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_1
X_15935_ _15935_/A _15935_/B _15935_/C _15934_/X vssd1 vssd1 vccd1 vccd1 _15936_/D
+ sky130_fd_sc_hd__or4b_1
X_11058_ _11058_/A vssd1 vssd1 vccd1 vccd1 _18254_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18001_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_237_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10009_ _10009_/A vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18654_ _18654_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17605_ _17609_/CLK _17605_/D vssd1 vssd1 vccd1 vccd1 _17605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18585_ _18585_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17536_ _17536_/CLK _17536_/D vssd1 vssd1 vccd1 vccd1 _17536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17467_ _17467_/A vssd1 vssd1 vccd1 vccd1 _19336_/D sky130_fd_sc_hd__clkbuf_1
X_14679_ _14679_/A _14679_/B vssd1 vssd1 vccd1 vccd1 _14679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19206_ _19206_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
X_16418_ _16418_/A _16418_/B _16418_/C vssd1 vssd1 vccd1 vccd1 _16419_/D sky130_fd_sc_hd__or3_1
XFILLER_220_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19137_ _19143_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14375__555 _14378__558/A vssd1 vssd1 vccd1 vccd1 _18190_/CLK sky130_fd_sc_hd__inv_2
XFILLER_195_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19068_ _19068_/CLK _19068_/D vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18019_ _18021_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _10695_/A vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__buf_4
XFILLER_234_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _10138_/C vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09585_ _18941_/Q _09486_/X _09591_/S vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__mux2_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _18590_/Q _09726_/X _10364_/S vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13111__415 _13111__415/A vssd1 vssd1 vccd1 vccd1 _17711_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14276__475 _14277__476/A vssd1 vssd1 vccd1 vccd1 _18110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_164_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _10583_/B _09894_/A _10583_/A vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__or3_4
X_10291_ _10291_/A vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__clkbuf_1
X_12030_ _12023_/X _12024_/X _12026_/X _12028_/X _11907_/S _12075_/A vssd1 vssd1 vccd1
+ vccd1 _12030_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307__209 _16307__209/A vssd1 vssd1 vccd1 vccd1 _18925_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13981_ _13786_/X _13973_/X _13978_/X vssd1 vssd1 vccd1 vccd1 _13981_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _12932_/A vssd1 vssd1 vccd1 vccd1 _12932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12863_ _18002_/Q _13024_/B vssd1 vssd1 vccd1 vccd1 _12915_/S sky130_fd_sc_hd__and2_2
XFILLER_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14662_/S vssd1 vssd1 vccd1 vccd1 _14726_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11814_ _17931_/Q _11785_/X _11800_/X _11813_/X vssd1 vssd1 vccd1 vccd1 _11814_/X
+ sky130_fd_sc_hd__o211a_4
X_18370_ _18370_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15579_/X _15580_/Y _15581_/X vssd1 vssd1 vccd1 vccd1 _18650_/D sky130_fd_sc_hd__a21oi_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12794_/A vssd1 vssd1 vccd1 vccd1 _17640_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17304_/X _17321_/B vssd1 vssd1 vccd1 vccd1 _17322_/A sky130_fd_sc_hd__and2b_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11745_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17252_/A _17252_/B vssd1 vssd1 vccd1 vccd1 _17253_/C sky130_fd_sc_hd__or2_1
Xclkbuf_0__03990_ _15787_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03990_/X sky130_fd_sc_hd__clkbuf_16
X_11676_ _12828_/A vssd1 vssd1 vccd1 vccd1 _13892_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_186_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _16191_/X _16193_/Y _16197_/Y _16200_/Y _16202_/Y vssd1 vssd1 vccd1 vccd1
+ _16203_/X sky130_fd_sc_hd__o32a_2
XFILLER_224_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13415_ _17789_/Q _13405_/B _13414_/Y _13376_/X vssd1 vssd1 vccd1 vccd1 _17789_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17183_ _17183_/A vssd1 vssd1 vccd1 vccd1 _19237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _10627_/A vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16134_ _10391_/X _16121_/X _16214_/A _16133_/Y vssd1 vssd1 vccd1 vccd1 _16134_/Y
+ sky130_fd_sc_hd__o211ai_2
X_13346_ _13330_/A _13346_/B vssd1 vssd1 vccd1 vccd1 _13346_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10558_ _18502_/Q _10129_/A _10562_/S vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15402__903 _15403__904/A vssd1 vssd1 vccd1 vccd1 _18590_/CLK sky130_fd_sc_hd__inv_2
XFILLER_127_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16065_ _16065_/A vssd1 vssd1 vccd1 vccd1 _18888_/D sky130_fd_sc_hd__clkbuf_1
X_13277_ _17752_/Q _13253_/X _13276_/Y vssd1 vssd1 vccd1 vccd1 _17752_/D sky130_fd_sc_hd__o21a_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10489_ _10489_/A vssd1 vssd1 vccd1 vccd1 _18533_/D sky130_fd_sc_hd__clkbuf_1
X_15016_ _15020_/B _15057_/A _15016_/C vssd1 vssd1 vccd1 vccd1 _15016_/X sky130_fd_sc_hd__and3b_1
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12159_ _12159_/A vssd1 vssd1 vccd1 vccd1 _17524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__04373_ clkbuf_0__04373_/X vssd1 vssd1 vccd1 vccd1 _16718_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03424_ _14889_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03424_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_209_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16967_ _16986_/A _16967_/B vssd1 vssd1 vccd1 vccd1 _16967_/Y sky130_fd_sc_hd__nor2_1
XFILLER_209_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18706_ _18706_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_1
X_15918_ _15917_/B _15917_/C _18866_/Q vssd1 vssd1 vccd1 vccd1 _15935_/C sky130_fd_sc_hd__a21oi_1
X_16898_ _19207_/Q _19159_/Q _18270_/Q _18262_/Q _16882_/A _16868_/X vssd1 vssd1 vccd1
+ vccd1 _16898_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15849_ _15855_/A vssd1 vssd1 vccd1 vccd1 _15849_/X sky130_fd_sc_hd__buf_1
X_18637_ _18637_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03186_ clkbuf_0__03186_/X vssd1 vssd1 vccd1 vccd1 _14472__633/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _09370_/A vssd1 vssd1 vccd1 vccd1 _19078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18568_ _18568_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17519_ _17737_/CLK _17519_/D vssd1 vssd1 vccd1 vccd1 _17519_/Q sky130_fd_sc_hd__dfxtp_1
X_18499_ _18499_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_4 _16559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09706_ _09682_/X _18895_/Q _09710_/S vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ _10219_/A _09636_/Y _09616_/X vssd1 vssd1 vccd1 vccd1 _09637_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_216_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09568_ _18948_/Q _09489_/X _09572_/S vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03413_ clkbuf_0__03413_/X vssd1 vssd1 vccd1 vccd1 _14838__764/A sky130_fd_sc_hd__clkbuf_16
XFILLER_54_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _19007_/Q _09498_/X _09505_/S vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11530_ _11545_/S vssd1 vssd1 vccd1 vccd1 _11539_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464__952 _15464__952/A vssd1 vssd1 vccd1 vccd1 _18639_/CLK sky130_fd_sc_hd__inv_2
XFILLER_221_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11461_ _11326_/X _18062_/Q _11467_/S vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16313__213 _16313__213/A vssd1 vssd1 vccd1 vccd1 _18929_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ input66/X _13446_/B vssd1 vssd1 vccd1 vccd1 _13374_/A sky130_fd_sc_hd__nand2_1
X_10412_ _10406_/X _10412_/B _10433_/C vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__and3b_1
XFILLER_171_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11392_ _11332_/X _18119_/Q _11394_/S vssd1 vssd1 vccd1 vccd1 _11393_/A sky130_fd_sc_hd__mux2_1
X_14180_ _13128_/A _11779_/A _16690_/A vssd1 vssd1 vccd1 vccd1 _14249_/A sky130_fd_sc_hd__a21o_2
XFILLER_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17005__354 _17005__354/A vssd1 vssd1 vccd1 vccd1 _19153_/CLK sky130_fd_sc_hd__inv_2
XFILLER_164_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13131_ _13873_/A _11826_/A _13873_/C vssd1 vssd1 vccd1 vccd1 _13132_/B sky130_fd_sc_hd__a21o_1
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10343_ _18596_/Q _10342_/X _10343_/S vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13062_ _13062_/A vssd1 vssd1 vccd1 vccd1 _17697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10274_ _10274_/A _10528_/B vssd1 vssd1 vccd1 vccd1 _10290_/S sky130_fd_sc_hd__nor2_2
XFILLER_140_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12013_ _11903_/X _12012_/X _12109_/S vssd1 vssd1 vccd1 vccd1 _12103_/A sky130_fd_sc_hd__mux2_1
X_17870_ _18031_/CLK _17870_/D vssd1 vssd1 vccd1 vccd1 _17870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15851__151 _15851__151/A vssd1 vssd1 vccd1 vccd1 _18826_/CLK sky130_fd_sc_hd__inv_2
XFILLER_239_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16821_ _16900_/A vssd1 vssd1 vccd1 vccd1 _16986_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16752_ _16786_/B vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13964_ _17967_/Q _13964_/B vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12915_ _17968_/Q _17668_/Q _12915_/S vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16683_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16683_/X sky130_fd_sc_hd__buf_1
XFILLER_206_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13895_ _13786_/X _13885_/X _13894_/X vssd1 vssd1 vccd1 vccd1 _13895_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_235_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15135__848 _15136__849/A vssd1 vssd1 vccd1 vccd1 _18524_/CLK sky130_fd_sc_hd__inv_2
X_18422_ _18422_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
X_15634_ _16054_/A _15638_/B vssd1 vssd1 vccd1 vccd1 _18661_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ _17648_/Q _12846_/B vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__xnor2_1
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18353_ _18353_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15565_ _15563_/X _15564_/Y _15553_/X vssd1 vssd1 vccd1 vccd1 _18647_/D sky130_fd_sc_hd__a21oi_1
XFILLER_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _18003_/Q _13024_/B vssd1 vssd1 vccd1 vccd1 _12831_/S sky130_fd_sc_hd__nand2_2
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17304_ _17437_/A vssd1 vssd1 vccd1 vccd1 _17304_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11728_/A vssd1 vssd1 vccd1 vccd1 _11728_/X sky130_fd_sc_hd__clkbuf_1
X_18284_ _18284_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ _18650_/Q vssd1 vssd1 vccd1 vccd1 _15585_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_230_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17235_ _17240_/B _17235_/B _17235_/C vssd1 vssd1 vccd1 vccd1 _17236_/A sky130_fd_sc_hd__and3b_1
Xclkbuf_0__03973_ _15705_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03973_/X sky130_fd_sc_hd__clkbuf_16
X_11659_ _17513_/Q _09679_/A _11665_/S vssd1 vssd1 vccd1 vccd1 _11660_/A sky130_fd_sc_hd__mux2_1
X_17166_ _17169_/C _17166_/B vssd1 vssd1 vccd1 vccd1 _19232_/D sky130_fd_sc_hd__nor2_1
XFILLER_174_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _16117_/A vssd1 vssd1 vccd1 vccd1 _16117_/X sky130_fd_sc_hd__buf_2
XFILLER_115_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13329_ _13330_/A vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__clkbuf_2
X_17097_ _17776_/Q _17774_/Q _17101_/C _17096_/Y vssd1 vssd1 vccd1 vccd1 _17097_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_192_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16048_ _16044_/A _16044_/B _18879_/Q vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__a21oi_1
XFILLER_157_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08870_ _08870_/A vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17999_ _18014_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03407_ _14802_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03407_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ _08925_/X _19055_/Q _09424_/S vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03169_ clkbuf_0__03169_/X vssd1 vssd1 vccd1 vccd1 _14449_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_164_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09353_ _09353_/A vssd1 vssd1 vccd1 vccd1 _19085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409__909 _15409__909/A vssd1 vssd1 vccd1 vccd1 _18596_/CLK sky130_fd_sc_hd__inv_2
XFILLER_240_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _09299_/S vssd1 vssd1 vccd1 vccd1 _09293_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03962_ clkbuf_0__03962_/X vssd1 vssd1 vccd1 vccd1 _15654__959/A sky130_fd_sc_hd__clkbuf_16
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ _08728_/X _08998_/Y input74/X vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__a21oi_4
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _08880_/X _18293_/Q hold9/X vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12700_ _12700_/A _12700_/B vssd1 vssd1 vccd1 vccd1 _17617_/D sky130_fd_sc_hd__nor2_1
XFILLER_232_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13680_ _17870_/Q _13660_/X _13679_/Y vssd1 vssd1 vccd1 vccd1 _17870_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10892_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _10892_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_231_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _12631_/A _12631_/B vssd1 vssd1 vccd1 vccd1 _12632_/C sky130_fd_sc_hd__or2_1
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _18574_/Q _15207_/A _15270_/X _15349_/X vssd1 vssd1 vccd1 vccd1 _18574_/D
+ sky130_fd_sc_hd__o211a_1
X_12562_ _12552_/Y _13085_/B _12828_/A vssd1 vssd1 vccd1 vccd1 _12563_/D sky130_fd_sc_hd__a21oi_1
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04376_ clkbuf_0__04376_/X vssd1 vssd1 vccd1 vccd1 _16349__241/A sky130_fd_sc_hd__clkbuf_16
XFILLER_184_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11513_ _18039_/Q _11321_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__mux2_1
X_15281_ _15281_/A vssd1 vssd1 vccd1 vccd1 _15281_/X sky130_fd_sc_hd__clkbuf_4
X_12493_ _12638_/B _12638_/A _12383_/X _17602_/Q _12443_/X _12390_/S vssd1 vssd1 vccd1
+ vccd1 _12493_/X sky130_fd_sc_hd__mux4_1
X_14232_ _18086_/Q input44/X _16997_/S vssd1 vssd1 vccd1 vccd1 _14233_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11444_ _18096_/Q _11267_/X _11448_/S vssd1 vssd1 vccd1 vccd1 _11445_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11375_ _11335_/X _18126_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _11376_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03189_ clkbuf_0__03189_/X vssd1 vssd1 vccd1 vccd1 _14484__642/A sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10326_ _09697_/X _18601_/Q _10326_/S vssd1 vssd1 vccd1 vccd1 _10327_/A sky130_fd_sc_hd__mux2_1
X_14094_ _18014_/Q _14091_/X _14093_/Y vssd1 vssd1 vccd1 vccd1 _18014_/D sky130_fd_sc_hd__o21a_1
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332__520 _14334__522/A vssd1 vssd1 vccd1 vccd1 _18155_/CLK sky130_fd_sc_hd__inv_2
X_18971_ _18971_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13045_/A vssd1 vssd1 vccd1 vccd1 _17692_/D sky130_fd_sc_hd__clkbuf_1
X_17922_ _17922_/CLK _17922_/D vssd1 vssd1 vccd1 vccd1 _17922_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10257_ _10272_/S vssd1 vssd1 vccd1 vccd1 _10266_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17853_ _17953_/CLK _17853_/D vssd1 vssd1 vccd1 vccd1 _17853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10188_ _10188_/A vssd1 vssd1 vccd1 vccd1 _18691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16804_ _16894_/A vssd1 vssd1 vccd1 vccd1 _16804_/X sky130_fd_sc_hd__clkbuf_2
X_14996_ _14996_/A vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__clkbuf_1
X_17784_ _17922_/CLK _17784_/D vssd1 vssd1 vccd1 vccd1 _17784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13947_ _13964_/B vssd1 vssd1 vccd1 vccd1 _13950_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _13885_/A vssd1 vssd1 vccd1 vccd1 _13878_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15617_ _15617_/A vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__clkbuf_1
X_18405_ _18405_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12829_ _17303_/A vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__buf_2
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19385_ input23/X vssd1 vssd1 vccd1 vccd1 _19385_/X sky130_fd_sc_hd__buf_6
X_16597_ _19027_/Q _16595_/B _16596_/Y vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__o21a_1
XFILLER_201_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ _15545_/X _15547_/Y _15624_/A vssd1 vssd1 vccd1 vccd1 _18644_/D sky130_fd_sc_hd__a21oi_1
X_18336_ _18336_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18267_ _18267_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
X_15479_ _17830_/Q _17829_/Q _15489_/B vssd1 vssd1 vccd1 vccd1 _15529_/B sky130_fd_sc_hd__or3_1
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17218_ _17225_/D _17235_/B _17218_/C vssd1 vssd1 vccd1 vccd1 _17219_/A sky130_fd_sc_hd__and3b_1
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18198_ _18198_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15858__157 _15859__158/A vssd1 vssd1 vccd1 vccd1 _18832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17149_ _19227_/Q _19226_/Q _17149_/C _17149_/D vssd1 vssd1 vccd1 vccd1 _17162_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_144_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _09971_/A _18557_/Q _09971_/C vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__and3_1
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08922_ _08921_/X _19297_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08853_ _08853_/A _08853_/B _08853_/C vssd1 vssd1 vccd1 vccd1 _09084_/C sky130_fd_sc_hd__or3_2
XFILLER_112_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _19348_/Q _08724_/X _08796_/S vssd1 vssd1 vccd1 vccd1 _08785_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_213_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09405_ _09405_/A vssd1 vssd1 vccd1 vccd1 _19063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09336_ _19092_/Q _08967_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09337_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09267_ _09267_/A vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _19158_/Q _09139_/X _09202_/S vssd1 vssd1 vccd1 vccd1 _09199_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11160_ _11159_/X _18213_/Q _11166_/S vssd1 vssd1 vccd1 vccd1 _11161_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10111_ _10111_/A vssd1 vssd1 vccd1 vccd1 _18719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ _11091_/A vssd1 vssd1 vccd1 vccd1 _18242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _18745_/Q _09959_/X _10046_/S vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _17910_/Q _13796_/X _13800_/Y vssd1 vssd1 vccd1 vccd1 _17910_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11993_ _19251_/Q _17237_/B _12025_/S vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__mux2_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16520_ _16520_/A _16530_/B vssd1 vssd1 vccd1 vccd1 _16521_/A sky130_fd_sc_hd__and2_1
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13732_ _13732_/A vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10944_ _10944_/A vssd1 vssd1 vccd1 vccd1 _18301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ _16464_/A _16451_/B vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__nor2_1
X_13663_ _17863_/Q _13659_/X _13662_/Y vssd1 vssd1 vccd1 vccd1 _17863_/D sky130_fd_sc_hd__o21a_1
XFILLER_147_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10875_ _18336_/Q _10797_/X _10879_/S vssd1 vssd1 vccd1 vccd1 _10876_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12614_ _17594_/Q _17593_/Q _17592_/Q _12614_/D vssd1 vssd1 vccd1 vccd1 _12630_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19170_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _17797_/Q _16382_/B vssd1 vssd1 vccd1 vccd1 _16383_/B sky130_fd_sc_hd__nand2_1
XFILLER_197_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13594_ _11714_/B _13425_/A _13597_/S vssd1 vssd1 vccd1 vccd1 _13595_/B sky130_fd_sc_hd__mux2_1
XFILLER_185_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18654_/CLK sky130_fd_sc_hd__clkbuf_16
X_18121_ _18121_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ _18573_/Q _15207_/X _15270_/X _15332_/X vssd1 vssd1 vccd1 vccd1 _18573_/D
+ sky130_fd_sc_hd__o211a_1
X_12545_ _17632_/Q vssd1 vssd1 vccd1 vccd1 _12746_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19135_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052_ _18052_/CLK _18052_/D vssd1 vssd1 vccd1 vccd1 _18052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ _15264_/A _15307_/A vssd1 vssd1 vccd1 vccd1 _15264_/X sky130_fd_sc_hd__or2b_1
X_12476_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12476_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ _14215_/A vssd1 vssd1 vccd1 vccd1 _18078_/D sky130_fd_sc_hd__clkbuf_1
X_11427_ _11427_/A vssd1 vssd1 vccd1 vccd1 _18104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11358_ _11358_/A vssd1 vssd1 vccd1 vccd1 _18134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10309_ _10309_/A vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__clkbuf_1
X_14077_ _12560_/S _13529_/A _14077_/S vssd1 vssd1 vccd1 vccd1 _14078_/B sky130_fd_sc_hd__mux2_1
X_18954_ _18954_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11289_ _18161_/Q _11264_/X _11295_/S vssd1 vssd1 vccd1 vccd1 _11290_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13028_ _13028_/A vssd1 vssd1 vccd1 vccd1 _17687_/D sky130_fd_sc_hd__clkbuf_1
X_17905_ _17922_/CLK _17905_/D vssd1 vssd1 vccd1 vccd1 _17905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18885_ _18996_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17836_ _18919_/CLK _17836_/D vssd1 vssd1 vccd1 vccd1 _17836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17767_ _19340_/CLK _17767_/D vssd1 vssd1 vccd1 vccd1 _17767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14979_ _18456_/Q _18455_/Q _14979_/C vssd1 vssd1 vccd1 vccd1 _14986_/B sky130_fd_sc_hd__and3_1
X_16718_ _16718_/A vssd1 vssd1 vccd1 vccd1 _16718_/X sky130_fd_sc_hd__buf_1
X_17698_ _17951_/CLK _17698_/D vssd1 vssd1 vccd1 vccd1 _17698_/Q sky130_fd_sc_hd__dfxtp_1
X_15864__161 _15867__164/A vssd1 vssd1 vccd1 vccd1 _18836_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _09894_/A _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__or3b_4
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16710__332 _16710__332/A vssd1 vssd1 vccd1 vccd1 _19107_/CLK sky130_fd_sc_hd__inv_2
X_18319_ _18319_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19299_ _19299_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
X_14339__526 _14339__526/A vssd1 vssd1 vccd1 vccd1 _18161_/CLK sky130_fd_sc_hd__inv_2
X_09052_ _09051_/X _19205_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_5_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09954_ _18476_/Q vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08905_ _19301_/Q _08801_/X _08907_/S vssd1 vssd1 vccd1 vccd1 _08906_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ hold22/X vssd1 vssd1 vccd1 vccd1 _11383_/B sky130_fd_sc_hd__inv_2
XFILLER_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ hold20/A _09148_/B vssd1 vssd1 vccd1 vccd1 _08838_/A sky130_fd_sc_hd__nand2_1
XFILLER_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _09612_/B _09611_/B _09612_/A vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03592_ clkbuf_0__03592_/X vssd1 vssd1 vccd1 vccd1 _15123__839/A sky130_fd_sc_hd__clkbuf_16
XFILLER_81_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10660_ _18426_/Q _09726_/X _10662_/S vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09319_ _09319_/A vssd1 vssd1 vccd1 vccd1 _19100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10591_ _10591_/A vssd1 vssd1 vccd1 vccd1 _18489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17394__87 _17395__88/A vssd1 vssd1 vccd1 vccd1 _19300_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12261_ _12261_/A vssd1 vssd1 vccd1 vccd1 _17553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _13750_/A _13995_/X _13992_/X vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11212_ _18191_/Q _11053_/X _11214_/S vssd1 vssd1 vccd1 vccd1 _11213_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12192_ _12192_/A _12192_/B _12191_/X vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__or3b_1
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11143_ _11223_/A hold18/X vssd1 vssd1 vccd1 vccd1 _11166_/S sky130_fd_sc_hd__or2_2
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput86 _11765_/X vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__buf_2
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput97 _11870_/X vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__buf_2
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11074_ _11074_/A vssd1 vssd1 vccd1 vccd1 _18249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15951_ _15951_/A _15951_/B vssd1 vssd1 vccd1 vccd1 _15951_/Y sky130_fd_sc_hd__nor2_1
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14902_ _14922_/B _17847_/Q _17846_/Q _14907_/A vssd1 vssd1 vccd1 vccd1 _14913_/B
+ sky130_fd_sc_hd__or4_2
X_10025_ _10025_/A vssd1 vssd1 vccd1 vccd1 _18753_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18670_ _18670_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17621_ _17621_/CLK _17621_/D vssd1 vssd1 vccd1 vccd1 _17621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14444__610 _14448__614/A vssd1 vssd1 vccd1 vccd1 _18245_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14833_ _14833_/A vssd1 vssd1 vccd1 vccd1 _14833_/X sky130_fd_sc_hd__buf_1
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17552_ _17776_/CLK _17552_/D vssd1 vssd1 vccd1 vccd1 _17552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _19241_/Q _19242_/Q _12007_/S vssd1 vssd1 vccd1 vccd1 _11976_/X sky130_fd_sc_hd__mux2_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ _13735_/B vssd1 vssd1 vccd1 vccd1 _13715_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16503_ _16503_/A _16503_/B vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__nor2_1
X_17483_ _19328_/Q _12206_/A _12199_/A _19335_/Q _17482_/Y vssd1 vssd1 vccd1 vccd1
+ _17483_/X sky130_fd_sc_hd__o221a_1
XFILLER_17_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10927_ _18308_/Q _10907_/X _10929_/S vssd1 vssd1 vccd1 vccd1 _10928_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14695_ _19080_/Q _18344_/Q _17578_/Q _18796_/Q _14568_/X _14569_/X vssd1 vssd1 vccd1
+ vccd1 _14696_/B sky130_fd_sc_hd__mux4_2
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19222_ _19266_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13646_ _13759_/A _13874_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__and3_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16434_ _18969_/Q _16440_/A _16433_/Y _16427_/X vssd1 vssd1 vccd1 vccd1 _16435_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_10858_ _10858_/A vssd1 vssd1 vccd1 vccd1 _18344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19153_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _18967_/Q _16464_/A _16364_/Y vssd1 vssd1 vccd1 vccd1 _18967_/D sky130_fd_sc_hd__a21o_1
X_13577_ _17837_/Q _16530_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13578_/B sky130_fd_sc_hd__mux2_1
X_10789_ _18994_/Q vssd1 vssd1 vccd1 vccd1 _10789_/X sky130_fd_sc_hd__buf_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18104_ _18104_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__04842_ _17031_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04842_/X sky130_fd_sc_hd__clkbuf_16
X_15316_ _18572_/Q _15207_/X _15270_/X _15315_/X vssd1 vssd1 vccd1 vccd1 _18572_/D
+ sky130_fd_sc_hd__o211a_1
X_12528_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12528_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19084_ _19084_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_1
X_16296_ _17810_/Q _08773_/X _13681_/A _16061_/B vssd1 vssd1 vccd1 vccd1 _18923_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18035_ _18035_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
X_15247_ _18998_/Q _18960_/Q _18952_/Q _17541_/Q _15209_/X _15218_/X vssd1 vssd1 vccd1
+ vccd1 _15247_/X sky130_fd_sc_hd__mux4_1
X_12459_ _12707_/A _17619_/Q _12706_/A _17621_/Q _12436_/S _12359_/A vssd1 vssd1 vccd1
+ vccd1 _12459_/X sky130_fd_sc_hd__mux4_2
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__07492_ _12235_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07492_/X sky130_fd_sc_hd__clkbuf_16
X_15178_ _18670_/Q vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ _18027_/Q _14115_/X _14128_/Y vssd1 vssd1 vccd1 vccd1 _18027_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03586_ _15092_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03586_/X sky130_fd_sc_hd__clkbuf_16
X_18937_ _18937_/CLK _18937_/D vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09670_ _18907_/Q _09277_/X _09672_/S vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18868_ _18869_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17819_ _17819_/CLK _17819_/D vssd1 vssd1 vccd1 vccd1 _17819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18799_ _19144_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16669__304 _16669__304/A vssd1 vssd1 vccd1 vccd1 _19078_/CLK sky130_fd_sc_hd__inv_2
XFILLER_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09104_ _10704_/A vssd1 vssd1 vccd1 vccd1 _09104_/X sky130_fd_sc_hd__buf_2
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09035_ _11329_/A vssd1 vssd1 vccd1 vccd1 _09035_/X sky130_fd_sc_hd__buf_4
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09937_ _10602_/B vssd1 vssd1 vccd1 vccd1 _10620_/A sky130_fd_sc_hd__buf_4
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17300__76 _17302__78/A vssd1 vssd1 vccd1 vccd1 _19272_/CLK sky130_fd_sc_hd__inv_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _16826_/A vssd1 vssd1 vccd1 vccd1 _09868_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _08819_/A vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A vssd1 vssd1 vccd1 vccd1 _18832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508__662 _14509__663/A vssd1 vssd1 vccd1 vccd1 _18297_/CLK sky130_fd_sc_hd__inv_2
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _17927_/Q _11815_/X _11824_/X _11848_/A vssd1 vssd1 vccd1 vccd1 _11830_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11761_ _11761_/A vssd1 vssd1 vccd1 vccd1 _11761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_242_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13507_/S vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10712_ _10712_/A vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14511_/A vssd1 vssd1 vccd1 vccd1 _14480_/X sky130_fd_sc_hd__buf_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _19040_/Q _16620_/B _18411_/Q vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__a21oi_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13431_ input62/X _13431_/B vssd1 vssd1 vccd1 vccd1 _13493_/A sky130_fd_sc_hd__nand2_2
XFILLER_139_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10643_ _10643_/A vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16150_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16150_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13362_ _13362_/A vssd1 vssd1 vccd1 vccd1 _13400_/A sky130_fd_sc_hd__buf_4
X_14851__774 _14851__774/A vssd1 vssd1 vccd1 vccd1 _18419_/CLK sky130_fd_sc_hd__inv_2
X_10574_ _10126_/X _18495_/Q _10574_/S vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _17553_/Q _17478_/B vssd1 vssd1 vccd1 vccd1 _12313_/X sky130_fd_sc_hd__xor2_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13293_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ _15032_/A _15043_/C vssd1 vssd1 vccd1 vccd1 _15032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ _12244_/A vssd1 vssd1 vccd1 vccd1 _17548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12175_ _12175_/A vssd1 vssd1 vccd1 vccd1 _17529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11126_ _18226_/Q _11042_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16983_ _18210_/Q _18130_/Q _19187_/Q _18258_/Q _16822_/X _16823_/X vssd1 vssd1 vccd1
+ vccd1 _16984_/B sky130_fd_sc_hd__mux4_1
XFILLER_110_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18722_ _18722_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15934_ _15922_/Y _15923_/X _15928_/Y _15931_/Y _15933_/Y vssd1 vssd1 vccd1 vccd1
+ _15934_/X sky130_fd_sc_hd__o2111a_1
X_11057_ _18254_/Q _11056_/X _11057_/S vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__mux2_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ _18760_/Q _09963_/X _10010_/S vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _18654_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17604_ _17611_/CLK _17604_/D vssd1 vssd1 vccd1 vccd1 _17604_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18584_ _18584_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409__582 _14410__583/A vssd1 vssd1 vccd1 vccd1 _18217_/CLK sky130_fd_sc_hd__inv_2
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _17535_/CLK _17535_/D vssd1 vssd1 vccd1 vccd1 _17535_/Q sky130_fd_sc_hd__dfxtp_1
X_11959_ _11953_/X _11957_/X _12091_/A vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__mux2_1
X_14747_ _14759_/A vssd1 vssd1 vccd1 vccd1 _14747_/X sky130_fd_sc_hd__buf_1
XFILLER_178_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17070__56 _17071__57/A vssd1 vssd1 vccd1 vccd1 _19205_/CLK sky130_fd_sc_hd__inv_2
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _17454_/X _17466_/B vssd1 vssd1 vccd1 vccd1 _17467_/A sky130_fd_sc_hd__and2b_1
X_14678_ _17585_/Q _18383_/Q _18391_/Q _18425_/Q _14574_/X _14637_/X vssd1 vssd1 vccd1
+ vccd1 _14679_/B sky130_fd_sc_hd__mux4_1
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19205_ _19205_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
X_13629_ _13629_/A _13629_/B vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__or2_1
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16417_ _16417_/A _16417_/B _16417_/C _16416_/Y vssd1 vssd1 vccd1 vccd1 _16418_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _17415_/A vssd1 vssd1 vccd1 vccd1 _17397_/X sky130_fd_sc_hd__buf_1
XFILLER_192_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19136_ _19136_/CLK _19136_/D vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14752__694 _14752__694/A vssd1 vssd1 vccd1 vccd1 _18337_/CLK sky130_fd_sc_hd__inv_2
XFILLER_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19067_ _19067_/CLK _19067_/D vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfxtp_1
X_16279_ _18444_/Q _18694_/Q _18702_/Q _18710_/Q _16198_/X _16102_/X vssd1 vssd1 vccd1
+ vccd1 _16280_/B sky130_fd_sc_hd__mux4_1
XFILLER_173_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18018_ _18021_/CLK _18018_/D vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04587_ clkbuf_0__04587_/X vssd1 vssd1 vccd1 vccd1 _16717__334/A sky130_fd_sc_hd__clkbuf_16
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09722_ _09722_/A vssd1 vssd1 vccd1 vccd1 _18860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09653_ _10075_/B vssd1 vssd1 vccd1 vccd1 _10138_/C sky130_fd_sc_hd__buf_2
XFILLER_227_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09584_ _09584_/A vssd1 vssd1 vccd1 vccd1 _18942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14794__728 _14795__729/A vssd1 vssd1 vccd1 vccd1 _18371_/CLK sky130_fd_sc_hd__inv_2
XFILLER_224_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09018_ _09861_/A _09879_/A vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__nand2_1
XFILLER_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10290_ _18617_/Q _10198_/X _10290_/S vssd1 vssd1 vccd1 vccd1 _10291_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13980_ _17972_/Q _13967_/X _13979_/Y vssd1 vssd1 vccd1 vccd1 _17972_/D sky130_fd_sc_hd__o21a_1
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12931_ _12931_/A _12931_/B _12931_/C _12931_/D vssd1 vssd1 vccd1 vccd1 _12931_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12862_ _16578_/A _12862_/B _12862_/C vssd1 vssd1 vccd1 vccd1 _17652_/D sky130_fd_sc_hd__nor3_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _17912_/Q _11812_/X _11809_/Y input13/X _11802_/X vssd1 vssd1 vccd1 vccd1
+ _11813_/X sky130_fd_sc_hd__a221o_1
X_14601_ _18854_/Q _18348_/Q _19189_/Q _18356_/Q _14599_/X _14600_/X vssd1 vssd1 vccd1
+ vccd1 _14601_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15581_/A vssd1 vssd1 vccd1 vccd1 _15581_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12761_/X _12793_/B vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__and2b_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17764_/Q _19279_/Q _17333_/S vssd1 vssd1 vccd1 vccd1 _17321_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11744_ _17770_/Q _17879_/Q vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__and2b_4
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _17262_/D vssd1 vssd1 vccd1 vccd1 _17258_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11675_ _11675_/A vssd1 vssd1 vccd1 vccd1 _12828_/A sky130_fd_sc_hd__buf_8
XFILLER_105_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13414_ _13414_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _13414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16202_ _16143_/X _16201_/X _16119_/X vssd1 vssd1 vccd1 vccd1 _16202_/Y sky130_fd_sc_hd__o21ai_1
X_17182_ _17184_/B _17189_/B _17182_/C vssd1 vssd1 vccd1 vccd1 _17183_/A sky130_fd_sc_hd__and3b_1
X_10626_ _18442_/Q _10120_/A _10630_/S vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14394_ _14400_/A vssd1 vssd1 vccd1 vccd1 _14394_/X sky130_fd_sc_hd__buf_1
XFILLER_167_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ _16234_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13345_ _17774_/Q vssd1 vssd1 vccd1 vccd1 _13346_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10557_ _10557_/A vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16064_ _16064_/A _16064_/B _16064_/C vssd1 vssd1 vccd1 vccd1 _16065_/A sky130_fd_sc_hd__and3_1
XFILLER_170_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13276_ _13274_/X _13259_/A _13275_/X vssd1 vssd1 vccd1 vccd1 _13276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10488_ _18533_/Q _10348_/X _10490_/S vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15015_ _18461_/Q _15005_/A _15005_/B _18462_/Q vssd1 vssd1 vccd1 vccd1 _15016_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _12149_/X _12158_/B vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__and2b_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04372_ clkbuf_0__04372_/X vssd1 vssd1 vccd1 vccd1 _16337__233/A sky130_fd_sc_hd__clkbuf_16
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03423_ _14883_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03423_/X sky130_fd_sc_hd__clkbuf_16
X_11109_ _11109_/A vssd1 vssd1 vccd1 vccd1 _18234_/D sky130_fd_sc_hd__clkbuf_1
X_12089_ _12082_/Y _12083_/Y _12084_/Y _12088_/Y _12034_/A _12020_/A vssd1 vssd1 vccd1
+ vccd1 _12184_/A sky130_fd_sc_hd__mux4_2
X_16966_ _18185_/Q _18177_/Q _18169_/Q _18161_/Q _16881_/X _16882_/X vssd1 vssd1 vccd1
+ vccd1 _16967_/B sky130_fd_sc_hd__mux4_1
XFILLER_110_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18705_ _18705_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15917_ _18866_/Q _15917_/B _15917_/C vssd1 vssd1 vccd1 vccd1 _15935_/B sky130_fd_sc_hd__and3_1
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16897_ _16895_/X _16896_/X _16982_/A vssd1 vssd1 vccd1 vccd1 _16897_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ _18636_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03185_ clkbuf_0__03185_/X vssd1 vssd1 vccd1 vccd1 _14463__625/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14381__560 _14382__561/A vssd1 vssd1 vccd1 vccd1 _18195_/CLK sky130_fd_sc_hd__inv_2
X_18567_ _18567_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_1
X_15779_ _15779_/A vssd1 vssd1 vccd1 vccd1 _15779_/X sky130_fd_sc_hd__buf_1
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17518_ _19339_/CLK _17518_/D vssd1 vssd1 vccd1 vccd1 _17518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18498_ _18498_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17449_ _17437_/X _17449_/B vssd1 vssd1 vccd1 vccd1 _17450_/A sky130_fd_sc_hd__and2b_1
XFILLER_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14457__620 _14460__623/A vssd1 vssd1 vccd1 vccd1 _18255_/CLK sky130_fd_sc_hd__inv_2
XFILLER_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19119_ _19119_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_5 _08874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _09705_/A vssd1 vssd1 vccd1 vccd1 _18896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236__380 _12239__383/A vssd1 vssd1 vccd1 vccd1 _17544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ _09639_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__04530_ clkbuf_0__04530_/X vssd1 vssd1 vccd1 vccd1 _16558__266/A sky130_fd_sc_hd__clkbuf_16
XFILLER_243_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _09567_/A vssd1 vssd1 vccd1 vccd1 _18949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14282__480 _14284__482/A vssd1 vssd1 vccd1 vccd1 _18115_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03412_ clkbuf_0__03412_/X vssd1 vssd1 vccd1 vccd1 _14832__759/A sky130_fd_sc_hd__clkbuf_16
XFILLER_54_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09498_ _18882_/Q vssd1 vssd1 vccd1 vccd1 _09498_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_223_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11460_ _11460_/A vssd1 vssd1 vccd1 vccd1 _18063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _15174_/B vssd1 vssd1 vccd1 vccd1 _10433_/C sky130_fd_sc_hd__clkbuf_2
X_11391_ _11391_/A vssd1 vssd1 vccd1 vccd1 _18120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _13540_/A _13130_/B _18068_/Q vssd1 vssd1 vccd1 vccd1 _13873_/C sky130_fd_sc_hd__or3b_2
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10342_ _18476_/Q vssd1 vssd1 vccd1 vccd1 _10342_/X sky130_fd_sc_hd__buf_2
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13061_ _13049_/X _13061_/B vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ _10273_/A vssd1 vssd1 vccd1 vccd1 _18625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12012_ _19254_/Q _19255_/Q _19256_/Q _19257_/Q _11995_/X _11938_/A vssd1 vssd1 vccd1
+ vccd1 _12012_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19288_/CLK sky130_fd_sc_hd__clkbuf_16
X_16820_ _16820_/A vssd1 vssd1 vccd1 vccd1 _16900_/A sky130_fd_sc_hd__buf_2
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16751_ _16775_/A _16751_/B vssd1 vssd1 vccd1 vccd1 _19128_/D sky130_fd_sc_hd__nor2_1
X_13963_ _16055_/A _13950_/B _13962_/Y _11697_/X vssd1 vssd1 vccd1 vccd1 _17966_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12914_ _12914_/A vssd1 vssd1 vccd1 vccd1 _17667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13894_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18421_ _18421_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12845_ _12845_/A vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__clkbuf_4
X_15633_ _15641_/B vssd1 vssd1 vccd1 vccd1 _15638_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18352_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12776_/A _12776_/B vssd1 vssd1 vccd1 vccd1 _13024_/B sky130_fd_sc_hd__nand2_4
XFILLER_199_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15564_ _18647_/Q _15569_/B vssd1 vssd1 vccd1 vccd1 _15564_/Y sky130_fd_sc_hd__nand2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/A vssd1 vssd1 vccd1 vccd1 _17437_/A sky130_fd_sc_hd__buf_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _17912_/Q _19128_/Q _11869_/B vssd1 vssd1 vccd1 vccd1 _11728_/A sky130_fd_sc_hd__mux2_8
X_15495_ _15494_/B _15494_/C _18651_/Q vssd1 vssd1 vccd1 vccd1 _15527_/C sky130_fd_sc_hd__a21oi_1
X_18283_ _18283_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ _17237_/C _17233_/C _17237_/B vssd1 vssd1 vccd1 vccd1 _17235_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_0__03972_ _15699_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03972_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_174_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11658_ _11658_/A vssd1 vssd1 vccd1 vccd1 _17514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10609_ _10609_/A vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__clkbuf_1
X_17165_ _19232_/Q _17158_/X _17164_/X vssd1 vssd1 vccd1 vccd1 _17166_/B sky130_fd_sc_hd__o21ai_1
XFILLER_128_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ _17578_/Q _10698_/A _11593_/S vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13328_ _14090_/A _14113_/B _14076_/B vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__and3_2
X_16116_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16117_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_171_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17096_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17096_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13259_ _13259_/A vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16047_ _16044_/A _16050_/A _16046_/Y _15242_/X vssd1 vssd1 vccd1 vccd1 _18878_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17998_ _18014_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03406_ _14796_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03406_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16949_ _18216_/Q _18200_/Q _18489_/Q _18192_/Q _09852_/A _09858_/A vssd1 vssd1 vccd1
+ vccd1 _16949_/X sky130_fd_sc_hd__mux4_2
XFILLER_226_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17016__12 _17016__12/A vssd1 vssd1 vccd1 vccd1 _19161_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _09421_/A vssd1 vssd1 vccd1 vccd1 _19056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _18619_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03168_ clkbuf_0__03168_/X vssd1 vssd1 vccd1 vccd1 _14385__564/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09352_ _19085_/Q _09274_/X _09356_/S vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03199_ _14536_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03199_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _10310_/A _09508_/A vssd1 vssd1 vccd1 vccd1 _09299_/S sky130_fd_sc_hd__nor2_2
XFILLER_240_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16078__193 _16079__194/A vssd1 vssd1 vccd1 vccd1 _18898_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08998_ _13645_/B _08998_/B vssd1 vssd1 vccd1 vccd1 _08998_/Y sky130_fd_sc_hd__nor2_4
XFILLER_248_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10960_ _10960_/A vssd1 vssd1 vccd1 vccd1 _18294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _18933_/Q vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ _10891_/A vssd1 vssd1 vccd1 vccd1 _18322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12630_ _17596_/Q _17595_/Q _12630_/C _12630_/D vssd1 vssd1 vccd1 vccd1 _12641_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_19_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12561_ _12561_/A vssd1 vssd1 vccd1 vccd1 _13085_/B sky130_fd_sc_hd__buf_4
XFILLER_240_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__04375_ clkbuf_0__04375_/X vssd1 vssd1 vccd1 vccd1 _16346__239/A sky130_fd_sc_hd__clkbuf_16
XFILLER_129_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ hold24/A vssd1 vssd1 vccd1 vccd1 _11521_/S sky130_fd_sc_hd__buf_2
X_14300_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__buf_1
XFILLER_211_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15280_ _15220_/X _15277_/X _15279_/X _15222_/X vssd1 vssd1 vccd1 vccd1 _15280_/X
+ sky130_fd_sc_hd__o211a_1
X_12492_ _12485_/X _12486_/X _12487_/X _12489_/X _12768_/S _12502_/A vssd1 vssd1 vccd1
+ vccd1 _12492_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14231_ _14231_/A vssd1 vssd1 vccd1 vccd1 _16997_/S sky130_fd_sc_hd__clkbuf_4
X_11443_ _11443_/A vssd1 vssd1 vccd1 vccd1 _18097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11374_ _11374_/A vssd1 vssd1 vccd1 vccd1 _18127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03188_ clkbuf_0__03188_/X vssd1 vssd1 vccd1 vccd1 _14505_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_153_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10325_ _10325_/A vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__clkbuf_1
X_14093_ _13717_/A _14092_/X _14060_/X vssd1 vssd1 vccd1 vccd1 _14093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18970_ _18971_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13032_/X _13044_/B vssd1 vssd1 vccd1 vccd1 _13045_/A sky130_fd_sc_hd__and2b_1
X_17921_ _17923_/CLK _17921_/D vssd1 vssd1 vccd1 vccd1 _17921_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _10546_/B _10620_/A vssd1 vssd1 vccd1 vccd1 _10272_/S sky130_fd_sc_hd__nor2_2
XFILLER_140_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15141__853 _15142__854/A vssd1 vssd1 vccd1 vccd1 _18529_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17852_ _18462_/CLK _17852_/D vssd1 vssd1 vccd1 vccd1 _17852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10187_ _18691_/Q _10186_/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _16893_/A vssd1 vssd1 vccd1 vccd1 _16803_/X sky130_fd_sc_hd__buf_2
XFILLER_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17783_ _19128_/CLK _17783_/D vssd1 vssd1 vccd1 vccd1 _17783_/Q sky130_fd_sc_hd__dfxtp_1
X_14289__486 _14290__487/A vssd1 vssd1 vccd1 vccd1 _18121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _15001_/A _14995_/B vssd1 vssd1 vccd1 vccd1 _14996_/A sky130_fd_sc_hd__and2_1
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13946_ _13964_/B vssd1 vssd1 vccd1 vccd1 _13946_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13877_ _14090_/A _16516_/D _14076_/C vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__and3_1
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18404_ _18404_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _15616_/A _15616_/B _15616_/C vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__and3_1
XFILLER_34_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ _12828_/A vssd1 vssd1 vccd1 vccd1 _17303_/A sky130_fd_sc_hd__buf_6
X_16596_ _16602_/A _16596_/B vssd1 vssd1 vccd1 vccd1 _16596_/Y sky130_fd_sc_hd__nor2_1
X_18335_ _18335_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15547_ _18644_/Q _15569_/B vssd1 vssd1 vccd1 vccd1 _15547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12759_/A _12759_/B _12759_/C vssd1 vssd1 vccd1 vccd1 _12760_/A sky130_fd_sc_hd__and3_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18266_ _18266_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15478_ _17831_/Q _15486_/B vssd1 vssd1 vccd1 vccd1 _15489_/B sky130_fd_sc_hd__or2_1
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17217_ _17216_/B _17216_/C _17216_/D _19247_/Q vssd1 vssd1 vccd1 vccd1 _17218_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_163_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18197_ _18197_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17148_ _19229_/Q _19228_/Q vssd1 vssd1 vccd1 vccd1 _17149_/D sky130_fd_sc_hd__and2_1
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09970_ _09970_/A vssd1 vssd1 vccd1 vccd1 _15174_/B sky130_fd_sc_hd__buf_4
XFILLER_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ _09682_/A vssd1 vssd1 vccd1 vccd1 _08921_/X sky130_fd_sc_hd__buf_2
XFILLER_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08852_ _08844_/Y _08846_/X _08847_/X _08851_/X vssd1 vssd1 vccd1 vccd1 _08853_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17088__70 _17297__74/A vssd1 vssd1 vccd1 vccd1 _19219_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08783_ _08805_/S vssd1 vssd1 vccd1 vccd1 _08796_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415__914 _15415__914/A vssd1 vssd1 vccd1 vccd1 _18601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__04369_ _16315_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04369_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09404_ _08925_/X _19063_/Q _09406_/S vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14502__657 _14503__658/A vssd1 vssd1 vccd1 vccd1 _18292_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _09335_/A vssd1 vssd1 vccd1 vccd1 _19093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09266_ _19125_/Q _09265_/X _09272_/S vssd1 vssd1 vccd1 vccd1 _09267_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09197_ _09197_/A vssd1 vssd1 vccd1 vccd1 _19159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10110_ _18719_/Q _10072_/X _10110_/S vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11090_ _08991_/X _18242_/Q _11098_/S vssd1 vssd1 vccd1 vccd1 _11091_/A sky130_fd_sc_hd__mux2_1
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _10041_/A vssd1 vssd1 vccd1 vccd1 _18746_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_216_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540__252 _16541__253/A vssd1 vssd1 vccd1 vccd1 _18998_/CLK sky130_fd_sc_hd__inv_2
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _13256_/X _13797_/X _13789_/X vssd1 vssd1 vccd1 vccd1 _13800_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11992_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__inv_2
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13731_ _17887_/Q _13719_/B _13730_/Y _13726_/X vssd1 vssd1 vccd1 vccd1 _17887_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ _18301_/Q _10904_/X hold16/A vssd1 vssd1 vccd1 vccd1 _10944_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16450_ _16453_/B _16440_/A _16449_/Y _16427_/X vssd1 vssd1 vccd1 vccd1 _16451_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13662_ _13281_/X _13660_/X _13661_/X vssd1 vssd1 vccd1 vccd1 _13662_/Y sky130_fd_sc_hd__a21oi_1
X_10874_ _10874_/A vssd1 vssd1 vccd1 vccd1 _18337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12613_ _12613_/A vssd1 vssd1 vccd1 vccd1 _17593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _13761_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13597_/S sky130_fd_sc_hd__nor2_1
X_16381_ _18980_/Q _16381_/B vssd1 vssd1 vccd1 vccd1 _16421_/A sky130_fd_sc_hd__xnor2_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14403__577 _14403__577/A vssd1 vssd1 vccd1 vccd1 _18212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_212_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18120_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_1
X_12544_ _12511_/X _18004_/Q _12845_/A _12543_/X vssd1 vssd1 vccd1 vccd1 _12563_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15332_ _15244_/X _15321_/X _15331_/X _15267_/X vssd1 vssd1 vccd1 vccd1 _15332_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_223_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18051_ _18051_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ _12369_/X _12473_/X _12547_/S vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__mux2_1
X_15263_ _18672_/Q _18578_/Q _17533_/Q _17508_/Q _15262_/X _09631_/A vssd1 vssd1 vccd1
+ vccd1 _15264_/A sky130_fd_sc_hd__mux4_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14214_ _18078_/Q input36/X _14218_/S vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__mux2_1
X_11426_ _18104_/Q _11267_/X _11430_/S vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295__490 _14297__492/A vssd1 vssd1 vccd1 vccd1 _18125_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_54_wb_clk_i clkbuf_leaf_54_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17629_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14145_ _14151_/A vssd1 vssd1 vccd1 vccd1 _14145_/X sky130_fd_sc_hd__buf_1
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11357_ _18134_/Q _11273_/X _11357_/S vssd1 vssd1 vccd1 vccd1 _11358_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10308_ _18609_/Q _10198_/X _10308_/S vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__mux2_1
X_14076_ _16689_/A _14076_/B _14076_/C vssd1 vssd1 vccd1 vccd1 _14077_/S sky130_fd_sc_hd__and3_4
XFILLER_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18953_ _18953_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11288_ _11288_/A vssd1 vssd1 vccd1 vccd1 _18162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13027_ _12992_/X _13027_/B vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__and2b_1
X_17904_ _17922_/CLK _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/Q sky130_fd_sc_hd__dfxtp_1
X_10239_ _10254_/S vssd1 vssd1 vccd1 vccd1 _10248_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_239_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18884_ _18886_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_2
X_16326__224 _16326__224/A vssd1 vssd1 vccd1 vccd1 _18940_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17835_ _18919_/CLK _17835_/D vssd1 vssd1 vccd1 vccd1 _17835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ _19290_/CLK _17766_/D vssd1 vssd1 vccd1 vccd1 _17766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ _14991_/A vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _17953_/Q _13929_/B vssd1 vssd1 vccd1 vccd1 _13929_/Y sky130_fd_sc_hd__nor2_1
X_17697_ _17951_/CLK _17697_/D vssd1 vssd1 vccd1 vccd1 _17697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16579_ _16579_/A vssd1 vssd1 vccd1 vccd1 _16585_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ _11222_/A _11068_/B _10987_/B vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__or3_2
X_18318_ _18318_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19298_ _19298_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _11341_/A vssd1 vssd1 vccd1 vccd1 _09051_/X sky130_fd_sc_hd__buf_2
XFILLER_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18249_ _18249_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15148__859 _15148__859/A vssd1 vssd1 vccd1 vccd1 _18535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15675__975 _15677__977/A vssd1 vssd1 vccd1 vccd1 _18692_/CLK sky130_fd_sc_hd__inv_2
X_09953_ _09953_/A vssd1 vssd1 vccd1 vccd1 _18779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08904_ _08904_/A vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _11068_/B vssd1 vssd1 vccd1 vccd1 _11456_/B sky130_fd_sc_hd__inv_2
XFILLER_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ hold21/X vssd1 vssd1 vccd1 vccd1 _09148_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _18930_/Q _18925_/Q vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__and2b_1
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03591_ clkbuf_0__03591_/X vssd1 vssd1 vccd1 vccd1 _15114__831/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _08941_/X _19100_/Q _09318_/S vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10590_ _09035_/X _18489_/Q _10594_/S vssd1 vssd1 vccd1 vccd1 _10591_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09249_ _18557_/Q _09971_/C vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__and2_1
XFILLER_193_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ _12245_/X _12260_/B vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__and2b_1
XFILLER_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _11211_/A vssd1 vssd1 vccd1 vccd1 _18192_/D sky130_fd_sc_hd__clkbuf_1
X_12191_ _17529_/Q _12298_/A _12182_/A _17518_/Q _12190_/Y vssd1 vssd1 vccd1 vccd1
+ _12191_/X sky130_fd_sc_hd__o221a_1
X_16726__340 _16728__342/A vssd1 vssd1 vccd1 vccd1 _19119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11142_ _11321_/A vssd1 vssd1 vccd1 vccd1 _11142_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_218_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 _11761_/X vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__buf_2
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11073_ _09031_/X _18249_/Q _11079_/S vssd1 vssd1 vccd1 vccd1 _11074_/A sky130_fd_sc_hd__mux2_1
X_15950_ _15949_/Y _17811_/Q _18876_/Q vssd1 vssd1 vccd1 vccd1 _15951_/B sky130_fd_sc_hd__a21oi_1
Xoutput98 _11719_/X vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__buf_2
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ _17851_/Q _17850_/Q _17849_/Q _14938_/A vssd1 vssd1 vccd1 vccd1 _14907_/A
+ sky130_fd_sc_hd__or4_1
X_10024_ _18753_/Q _09959_/X _10028_/S vssd1 vssd1 vccd1 vccd1 _10025_/A sky130_fd_sc_hd__mux2_1
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _17621_/CLK _17620_/D vssd1 vssd1 vccd1 vccd1 _17620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _17772_/CLK _17551_/D vssd1 vssd1 vccd1 vccd1 _17551_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_101_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18996_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ _19239_/Q _19240_/Q _11975_/S vssd1 vssd1 vccd1 vccd1 _11975_/X sky130_fd_sc_hd__mux2_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17082__65 _17083__66/A vssd1 vssd1 vccd1 vccd1 _19214_/CLK sky130_fd_sc_hd__inv_2
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _18983_/Q _16429_/Y _16498_/C _16426_/A _16362_/A vssd1 vssd1 vccd1 vccd1
+ _16503_/B sky130_fd_sc_hd__a311o_1
XFILLER_232_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _13769_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13735_/B sky130_fd_sc_hd__or2_2
XFILLER_45_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17482_ _19328_/Q _12206_/A _12212_/A _19332_/Q _17481_/X vssd1 vssd1 vccd1 vccd1
+ _17482_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _10926_/A vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14694_ _14732_/A _14694_/B vssd1 vssd1 vccd1 vccd1 _14694_/Y sky130_fd_sc_hd__nor2_1
X_19221_ _19281_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16433_ _18969_/Q _16437_/C vssd1 vssd1 vccd1 vccd1 _16433_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13645_ _13645_/A _13645_/B vssd1 vssd1 vccd1 vccd1 _16688_/B sky130_fd_sc_hd__nor2_1
X_10857_ _18344_/Q _10797_/X _10861_/S vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19152_ _19152_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16426_/A _16469_/A vssd1 vssd1 vccd1 vccd1 _16364_/Y sky130_fd_sc_hd__nor2_1
X_13576_ _17454_/A vssd1 vssd1 vccd1 vccd1 _13629_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10788_ _10788_/A vssd1 vssd1 vccd1 vccd1 _18371_/D sky130_fd_sc_hd__clkbuf_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18103_ _18103_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__04841_ _17025_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04841_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15315_ _15244_/X _15297_/X _15314_/X _15267_/X vssd1 vssd1 vccd1 vccd1 _15315_/X
+ sky130_fd_sc_hd__a211o_1
X_12527_ _14067_/B _12452_/X _12510_/X _12526_/X vssd1 vssd1 vccd1 vccd1 _12527_/X
+ sky130_fd_sc_hd__o211a_1
X_19083_ _19083_/CLK _19083_/D vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfxtp_1
X_16295_ _16295_/A vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _18034_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__07560_ _12345_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07560_/X sky130_fd_sc_hd__clkbuf_16
X_15246_ _19113_/Q _18944_/Q _18602_/Q _19342_/Q _15245_/X _09626_/A vssd1 vssd1 vccd1
+ vccd1 _15246_/X sky130_fd_sc_hd__mux4_1
X_12458_ _12378_/X _12353_/X _12464_/S vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14451__615 _14451__615/A vssd1 vssd1 vccd1 vccd1 _18250_/CLK sky130_fd_sc_hd__inv_2
X_11409_ _11409_/A vssd1 vssd1 vccd1 vccd1 _18112_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__07491_ _12229_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07491_/X sky130_fd_sc_hd__clkbuf_16
X_12389_ _17606_/Q _17607_/Q _12435_/A vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
X_15177_ _15177_/A _15177_/B vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__nor2_1
XFILLER_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547__258 _16547__258/A vssd1 vssd1 vccd1 vccd1 _19004_/CLK sky130_fd_sc_hd__inv_2
XFILLER_158_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14128_ _13414_/A _14120_/X _14123_/X vssd1 vssd1 vccd1 vccd1 _14128_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03585_ _15086_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03585_/X sky130_fd_sc_hd__clkbuf_16
X_14059_ _18001_/Q _14054_/X _14058_/Y vssd1 vssd1 vccd1 vccd1 _18001_/D sky130_fd_sc_hd__o21a_1
X_18936_ _18936_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18867_ _18889_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _19339_/CLK _17818_/D vssd1 vssd1 vccd1 vccd1 _17818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18798_ _18798_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17749_ _19327_/CLK _17749_/D vssd1 vssd1 vccd1 vccd1 _17749_/Q sky130_fd_sc_hd__dfxtp_1
X_14345__531 _14347__533/A vssd1 vssd1 vccd1 vccd1 _18166_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230__375 _12230__375/A vssd1 vssd1 vccd1 vccd1 _17539_/CLK sky130_fd_sc_hd__inv_2
XFILLER_196_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16634__275 _16635__276/A vssd1 vssd1 vccd1 vccd1 _19049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09103_ _18990_/Q vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__buf_2
XFILLER_248_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09034_ _18666_/Q vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_191_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _10432_/A _09971_/A _09936_/C vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__or3_4
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _09867_/A vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _19321_/Q _08789_/X _08822_/S vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _18832_/Q _09755_/X _09800_/S vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__mux2_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _13541_/A _13759_/B _09253_/A vssd1 vssd1 vccd1 vccd1 _08749_/X sky130_fd_sc_hd__and3b_1
XFILLER_22_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11760_ _18001_/Q _17883_/Q vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__and2b_2
XFILLER_42_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _18404_/Q _10710_/X _10714_/S vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__mux2_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11691_ _19039_/Q _16619_/B vssd1 vssd1 vccd1 vccd1 _16620_/B sky130_fd_sc_hd__and2_1
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13430_ _17793_/Q vssd1 vssd1 vccd1 vccd1 _13430_/Y sky130_fd_sc_hd__inv_2
X_10642_ _09262_/X _18435_/Q _10648_/S vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__mux2_1
X_15428__924 _15428__924/A vssd1 vssd1 vccd1 vccd1 _18611_/CLK sky130_fd_sc_hd__inv_2
XFILLER_220_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13361_ _17776_/Q vssd1 vssd1 vccd1 vccd1 _13361_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10573_ _10573_/A vssd1 vssd1 vccd1 vccd1 _18496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15100_ _15100_/A vssd1 vssd1 vccd1 vccd1 _15100_/X sky130_fd_sc_hd__buf_1
X_12312_ _17549_/Q _12187_/X _12199_/X _17559_/Q vssd1 vssd1 vccd1 vccd1 _12315_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_13292_ _17756_/Q _13280_/X _13291_/Y vssd1 vssd1 vccd1 vccd1 _17756_/D sky130_fd_sc_hd__o21a_1
X_16080_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16080_/X sky130_fd_sc_hd__buf_1
XFILLER_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12243_ _12166_/X _12243_/B vssd1 vssd1 vccd1 vccd1 _12244_/A sky130_fd_sc_hd__and2b_1
X_15031_ _18465_/Q _18464_/Q _15031_/C vssd1 vssd1 vccd1 vccd1 _15043_/C sky130_fd_sc_hd__and3_1
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14515__667 _14517__669/A vssd1 vssd1 vccd1 vccd1 _18302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12174_ _12166_/X _12174_/B vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__and2b_1
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11125_ _11140_/S vssd1 vssd1 vccd1 vccd1 _11134_/S sky130_fd_sc_hd__buf_2
XFILLER_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16982_ _16982_/A _16982_/B vssd1 vssd1 vccd1 vccd1 _16982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15097__817 _15099__819/A vssd1 vssd1 vccd1 vccd1 _18493_/CLK sky130_fd_sc_hd__inv_2
X_18721_ _18721_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15933_ _18865_/Q _15933_/B vssd1 vssd1 vccd1 vccd1 _15933_/Y sky130_fd_sc_hd__xnor2_1
X_11056_ _18664_/Q vssd1 vssd1 vccd1 vccd1 _11056_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _10007_/A vssd1 vssd1 vccd1 vccd1 _18761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _18654_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17603_ _17611_/CLK _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14815_/X sky130_fd_sc_hd__buf_1
XFILLER_236_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _18583_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17534_/CLK _17534_/D vssd1 vssd1 vccd1 vccd1 _17534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14808_/A vssd1 vssd1 vccd1 vccd1 _14746_/X sky130_fd_sc_hd__buf_1
XFILLER_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11958_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17465_ _17740_/Q _19336_/Q _17468_/S vssd1 vssd1 vccd1 vccd1 _17466_/B sky130_fd_sc_hd__mux2_1
X_10909_ _10909_/A vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14677_ _14696_/A _14677_/B vssd1 vssd1 vccd1 vccd1 _14677_/Y sky130_fd_sc_hd__nor2_1
X_11889_ _19246_/Q vssd1 vssd1 vccd1 vccd1 _17216_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19204_ _19204_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16553__262 _16555__264/A vssd1 vssd1 vccd1 vccd1 _19008_/CLK sky130_fd_sc_hd__inv_2
X_16416_ _16453_/B _16416_/B vssd1 vssd1 vccd1 vccd1 _16416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13628_ _17854_/Q _16530_/A _13635_/B vssd1 vssd1 vccd1 vccd1 _13629_/B sky130_fd_sc_hd__mux2_1
XFILLER_193_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19135_ _19135_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ _16543_/A vssd1 vssd1 vccd1 vccd1 _16347_/X sky130_fd_sc_hd__buf_1
X_13559_ _17831_/Q _13446_/X _13559_/S vssd1 vssd1 vccd1 vccd1 _13560_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19066_ _19066_/CLK _19066_/D vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16278_ _16278_/A _16278_/B vssd1 vssd1 vccd1 vccd1 _16278_/Y sky130_fd_sc_hd__nor2_1
X_18017_ _18021_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ _15220_/X _15226_/X _15228_/X _15222_/X vssd1 vssd1 vccd1 vccd1 _15229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16072__188 _16073__189/A vssd1 vssd1 vccd1 vccd1 _18893_/CLK sky130_fd_sc_hd__inv_2
XFILLER_154_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04586_ clkbuf_0__04586_/X vssd1 vssd1 vccd1 vccd1 _16704__327/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14828__755 _14829__756/A vssd1 vssd1 vccd1 vccd1 _18398_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09721_ _18860_/Q _09718_/X _09733_/S vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__mux2_1
X_18919_ _18919_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _10437_/B vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__03399_ clkbuf_0__03399_/X vssd1 vssd1 vccd1 vccd1 _14763__703/A sky130_fd_sc_hd__clkbuf_16
XFILLER_227_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09583_ _18942_/Q _09481_/X _09591_/S vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__mux2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15877__172 _15879__174/A vssd1 vssd1 vccd1 vccd1 _18847_/CLK sky130_fd_sc_hd__inv_2
XFILLER_163_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ _09016_/X _18800_/Q vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__and2b_4
XFILLER_191_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09919_ _09919_/A vssd1 vssd1 vccd1 vccd1 _18790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12930_ _17660_/Q _12921_/X _12838_/X _17668_/Q _12929_/X vssd1 vssd1 vccd1 vccd1
+ _12931_/D sky130_fd_sc_hd__a221oi_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12861_ _12836_/X _12860_/X _17652_/Q vssd1 vssd1 vccd1 vccd1 _12862_/C sky130_fd_sc_hd__o21ba_1
XFILLER_206_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14627_/A vssd1 vssd1 vccd1 vccd1 _14600_/X sky130_fd_sc_hd__buf_2
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11812_/A vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15585_/B _15597_/B vssd1 vssd1 vccd1 vccd1 _15580_/Y sky130_fd_sc_hd__nand2_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _17640_/Q _17995_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12793_/B sky130_fd_sc_hd__mux2_1
XFILLER_199_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A vssd1 vssd1 vccd1 vccd1 _11743_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_242_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17250_ _17252_/A _17250_/B _17250_/C _17250_/D vssd1 vssd1 vccd1 vccd1 _17262_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14474_/A vssd1 vssd1 vccd1 vccd1 _14462_/X sky130_fd_sc_hd__buf_1
XFILLER_175_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11674_ input2/X vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__inv_8
XFILLER_70_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16201_ _18448_/Q _19086_/Q _19123_/Q _18432_/Q _16144_/X _10420_/X vssd1 vssd1 vccd1
+ vccd1 _16201_/X sky130_fd_sc_hd__mux4_2
X_13413_ _17788_/Q _13393_/X _13412_/Y vssd1 vssd1 vccd1 vccd1 _17788_/D sky130_fd_sc_hd__o21a_1
X_17181_ _17179_/B _17180_/A _19237_/Q vssd1 vssd1 vccd1 vccd1 _17182_/C sky130_fd_sc_hd__a21o_1
X_10625_ _10625_/A vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16132_ _16125_/X _16130_/X _16162_/S vssd1 vssd1 vccd1 vccd1 _16133_/B sky130_fd_sc_hd__mux2_1
X_13344_ input73/X _16518_/B _13329_/X _13342_/X _13343_/X vssd1 vssd1 vccd1 vccd1
+ _17773_/D sky130_fd_sc_hd__a311o_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ _18503_/Q _10126_/A _10556_/S vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16063_ _16063_/A _16063_/B vssd1 vssd1 vccd1 vccd1 _16064_/C sky130_fd_sc_hd__nand2_1
X_13275_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__clkbuf_2
X_10487_ _10487_/A vssd1 vssd1 vccd1 vccd1 _18534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _18462_/Q _18461_/Q _15014_/C vssd1 vssd1 vccd1 vccd1 _15020_/B sky130_fd_sc_hd__and3_1
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105__824 _15105__824/A vssd1 vssd1 vccd1 vccd1 _18500_/CLK sky130_fd_sc_hd__inv_2
XFILLER_151_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ _17524_/Q _17727_/Q _12170_/S vssd1 vssd1 vccd1 vccd1 _12158_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04371_ clkbuf_0__04371_/X vssd1 vssd1 vccd1 vccd1 _16329__226/A sky130_fd_sc_hd__clkbuf_16
XFILLER_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11108_ _18234_/Q _11042_/X _11116_/S vssd1 vssd1 vccd1 vccd1 _11109_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03422_ _14877_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03422_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12088_ _12088_/A vssd1 vssd1 vccd1 vccd1 _12088_/Y sky130_fd_sc_hd__inv_2
X_16965_ _16984_/A _16965_/B vssd1 vssd1 vccd1 vccd1 _16965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15916_ _17821_/Q _15932_/B _17820_/Q vssd1 vssd1 vccd1 vccd1 _15917_/C sky130_fd_sc_hd__o21ai_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ _11039_/A vssd1 vssd1 vccd1 vccd1 _18260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _18704_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16896_ _18150_/Q _18142_/Q _18134_/Q _18278_/Q _16803_/X _16804_/X vssd1 vssd1 vccd1
+ vccd1 _16896_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18635_ _18635_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14149__433 _14149__433/A vssd1 vssd1 vccd1 vccd1 _18041_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03184_ clkbuf_0__03184_/X vssd1 vssd1 vccd1 vccd1 _14460__623/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18566_ _18566_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17517_ _19339_/CLK _17517_/D vssd1 vssd1 vccd1 vccd1 _17517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14729_ _14727_/X _14728_/X _14729_/S vssd1 vssd1 vccd1 vccd1 _14729_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18497_ _18497_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _17745_/Q _19331_/Q _17451_/S vssd1 vssd1 vccd1 vccd1 _17449_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17379_ _19289_/Q _12298_/X _12182_/X _19278_/Q _17378_/X vssd1 vssd1 vccd1 vccd1
+ _17379_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18922_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19118_ _19118_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19049_ _19049_/CLK _19049_/D vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_238_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04569_ clkbuf_0__04569_/X vssd1 vssd1 vccd1 vccd1 _16635__276/A sky130_fd_sc_hd__clkbuf_16
XFILLER_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_6 _09016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09704_ _09679_/X _18896_/Q _09710_/S vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09635_ _09635_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09643_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ _18949_/Q _09486_/X _09572_/S vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03411_ clkbuf_0__03411_/X vssd1 vssd1 vccd1 vccd1 _14826__754/A sky130_fd_sc_hd__clkbuf_16
XFILLER_230_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ _09497_/A vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358__541 _14358__541/A vssd1 vssd1 vccd1 vccd1 _18176_/CLK sky130_fd_sc_hd__inv_2
X_10410_ _10406_/B _10405_/A _10405_/B _10406_/A vssd1 vssd1 vccd1 vccd1 _10412_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__05012_ clkbuf_0__05012_/X vssd1 vssd1 vccd1 vccd1 _17302__78/A sky130_fd_sc_hd__clkbuf_16
X_11390_ _11329_/X _18120_/Q _11394_/S vssd1 vssd1 vccd1 vccd1 _11391_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _10341_/A vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13060_ _17941_/Q _17697_/Q _13070_/S vssd1 vssd1 vccd1 vccd1 _13061_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16647__285 _16649__287/A vssd1 vssd1 vccd1 vccd1 _19059_/CLK sky130_fd_sc_hd__inv_2
X_10272_ _18625_/Q _10198_/X _10272_/S vssd1 vssd1 vccd1 vccd1 _10273_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17489_/B sky130_fd_sc_hd__buf_4
XFILLER_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17411__101 _17412__102/A vssd1 vssd1 vccd1 vccd1 _19314_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16750_ _16762_/A _16740_/Y _16749_/Y _16687_/B vssd1 vssd1 vccd1 vccd1 _16751_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13962_ _17966_/Q _13962_/B vssd1 vssd1 vccd1 vccd1 _13962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17618_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12913_ _12911_/X _12913_/B vssd1 vssd1 vccd1 vccd1 _12914_/A sky130_fd_sc_hd__and2b_1
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13893_ _14095_/A vssd1 vssd1 vccd1 vccd1 _13992_/A sky130_fd_sc_hd__clkbuf_2
X_16320__219 _16320__219/A vssd1 vssd1 vccd1 vccd1 _18935_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18420_ _18420_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15632_ _08998_/B _15808_/B _16052_/C vssd1 vssd1 vccd1 vccd1 _15641_/B sky130_fd_sc_hd__nand3b_4
X_12844_ _17641_/Q _13095_/B vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__xor2_1
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18351_ _18351_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15579_/A _15563_/B _15572_/C vssd1 vssd1 vccd1 vccd1 _15563_/X sky130_fd_sc_hd__or3_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12561_/A _12775_/B _12775_/C _12775_/D vssd1 vssd1 vccd1 vccd1 _12776_/B
+ sky130_fd_sc_hd__and4b_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04589_ clkbuf_0__04589_/X vssd1 vssd1 vccd1 vccd1 _17000_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_203_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11726_/A vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18282_ _18282_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15494_ _18651_/Q _15494_/B _15494_/C vssd1 vssd1 vccd1 vccd1 _15527_/B sky130_fd_sc_hd__and3_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17233_ _17237_/B _17237_/C _17233_/C vssd1 vssd1 vccd1 vccd1 _17240_/B sky130_fd_sc_hd__and3_1
XFILLER_35_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03971_ _15693_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03971_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_202_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11657_ _17514_/Q _09674_/A _11665_/S vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17164_ _17191_/A vssd1 vssd1 vccd1 vccd1 _17164_/X sky130_fd_sc_hd__clkbuf_2
X_10608_ _10120_/X _18450_/Q _10612_/S vssd1 vssd1 vccd1 vccd1 _10609_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11588_ _11588_/A vssd1 vssd1 vccd1 vccd1 _17579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16115_ _18565_/Q vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__buf_2
XFILLER_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _14053_/B vssd1 vssd1 vccd1 vccd1 _14076_/B sky130_fd_sc_hd__buf_2
XFILLER_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17095_ _17091_/X _17094_/X _17101_/C vssd1 vssd1 vccd1 vccd1 _17109_/A sky130_fd_sc_hd__a21o_1
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10539_ _10539_/A vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16044_/Y _16045_/X _16050_/A vssd1 vssd1 vccd1 vccd1 _16046_/Y sky130_fd_sc_hd__o21ai_1
X_13258_ _17746_/Q _13252_/X _13257_/Y vssd1 vssd1 vccd1 vccd1 _17746_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12209_ _17519_/Q _12206_/A _12212_/A _17523_/Q _12208_/X vssd1 vssd1 vccd1 vccd1
+ _12209_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13189_ _13216_/B vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17997_ _18014_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03405_ _14790_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03405_/X sky130_fd_sc_hd__clkbuf_16
X_16948_ _16986_/A _16948_/B vssd1 vssd1 vccd1 vccd1 _16948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_237_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16879_ _18205_/Q _18125_/Q _19182_/Q _18253_/Q _16827_/X _16828_/X vssd1 vssd1 vccd1
+ vccd1 _16880_/B sky130_fd_sc_hd__mux4_1
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ _08921_/X _19056_/Q _09424_/S vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15828__133 _15829__134/A vssd1 vssd1 vccd1 vccd1 _18808_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _18618_/CLK _18618_/D vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03167_ clkbuf_0__03167_/X vssd1 vssd1 vccd1 vccd1 _14379__559/A sky130_fd_sc_hd__clkbuf_16
XFILLER_213_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03198_ _14530_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03198_/X sky130_fd_sc_hd__clkbuf_16
X_09351_ _09351_/A vssd1 vssd1 vccd1 vccd1 _19086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18549_ _18549_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03098_ clkbuf_0__03098_/X vssd1 vssd1 vccd1 vccd1 _14255__459/A sky130_fd_sc_hd__clkbuf_16
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14162__441 _14162__441/A vssd1 vssd1 vccd1 vccd1 _18049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_221_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09282_ _09282_/A vssd1 vssd1 vccd1 vccd1 _19120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16720__335 _16723__338/A vssd1 vssd1 vccd1 vccd1 _19114_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08997_ _13540_/B _13520_/B _08997_/C vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__or3_4
XFILLER_68_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09618_ _09600_/X _09615_/X _09617_/Y vssd1 vssd1 vccd1 vccd1 _18934_/D sky130_fd_sc_hd__o21a_1
XFILLER_189_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _18322_/Q _10887_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10891_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09549_ _09549_/A vssd1 vssd1 vccd1 vccd1 _18957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12560_ _12558_/X _12559_/X _12560_/S vssd1 vssd1 vccd1 vccd1 _12561_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04374_ clkbuf_0__04374_/X vssd1 vssd1 vccd1 vccd1 _16359_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_240_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11511_/A hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__nor2_2
XFILLER_54_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12491_ _12538_/A vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__clkbuf_2
X_14230_ _14230_/A vssd1 vssd1 vccd1 vccd1 _18085_/D sky130_fd_sc_hd__clkbuf_1
X_11442_ _18097_/Q _11264_/X _11448_/S vssd1 vssd1 vccd1 vccd1 _11443_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15769__1051 _15771__1053/A vssd1 vssd1 vccd1 vccd1 _18768_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _11332_/X _18127_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _11374_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03187_ clkbuf_0__03187_/X vssd1 vssd1 vccd1 vccd1 _14479__639/A sky130_fd_sc_hd__clkbuf_16
X_10324_ _09694_/X _18602_/Q _10326_/S vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__mux2_1
X_14092_ _14099_/A vssd1 vssd1 vccd1 vccd1 _14092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13043_ _17946_/Q _17692_/Q _13053_/S vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__mux2_1
X_17920_ _17923_/CLK _17920_/D vssd1 vssd1 vccd1 vccd1 _17920_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10255_/A vssd1 vssd1 vccd1 vccd1 _18633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17851_ _18462_/CLK _17851_/D vssd1 vssd1 vccd1 vccd1 _17851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ _18477_/Q vssd1 vssd1 vccd1 vccd1 _10186_/X sky130_fd_sc_hd__buf_4
XFILLER_65_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16802_ _18115_/Q _18107_/Q _18099_/Q _18091_/Q _16799_/X _16801_/X vssd1 vssd1 vccd1
+ vccd1 _16802_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17782_ _19281_/CLK _17782_/D vssd1 vssd1 vccd1 vccd1 _17782_/Q sky130_fd_sc_hd__dfxtp_1
X_14994_ _18458_/Q _14991_/X _14992_/X _14993_/X vssd1 vssd1 vccd1 vccd1 _14995_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13945_ _14113_/A _13945_/B vssd1 vssd1 vccd1 vccd1 _13964_/B sky130_fd_sc_hd__and2_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16664_ _16670_/A vssd1 vssd1 vccd1 vccd1 _16664_/X sky130_fd_sc_hd__buf_1
XFILLER_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13876_ _14053_/C vssd1 vssd1 vccd1 vccd1 _14076_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15615_ _18657_/Q _15615_/B _15615_/C vssd1 vssd1 vccd1 vccd1 _15616_/C sky130_fd_sc_hd__nand3_1
X_18403_ _18403_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ _12827_/A vssd1 vssd1 vccd1 vccd1 _17650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16595_ _16613_/A _16595_/B _16595_/C vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__nor3_1
XFILLER_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _18334_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15546_ _15612_/B vssd1 vssd1 vccd1 vccd1 _15569_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _17635_/Q _12758_/B _12758_/C _12758_/D vssd1 vssd1 vccd1 vccd1 _12759_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11709_ _17843_/Q vssd1 vssd1 vccd1 vccd1 _11714_/B sky130_fd_sc_hd__inv_2
X_18265_ _18265_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15477_ _17832_/Q _15494_/B vssd1 vssd1 vccd1 vccd1 _15486_/B sky130_fd_sc_hd__or2_1
X_12689_ _12687_/X _12709_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12690_/A sky130_fd_sc_hd__and3b_1
XFILLER_175_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17216_ _19247_/Q _17216_/B _17216_/C _17216_/D vssd1 vssd1 vccd1 vccd1 _17225_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18196_ _18196_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17147_ _11978_/X _17142_/X _17146_/Y vssd1 vssd1 vccd1 vccd1 _19228_/D sky130_fd_sc_hd__a21oi_1
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17418__107 _17419__108/A vssd1 vssd1 vccd1 vccd1 _19320_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08920_ _18885_/Q vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__buf_4
X_16029_ _18874_/Q _16024_/C _16028_/X _15242_/X vssd1 vssd1 vccd1 vccd1 _18874_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08851_ _09440_/A _09440_/B _09441_/C vssd1 vssd1 vccd1 vccd1 _08851_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08782_ _09745_/A _10310_/A vssd1 vssd1 vccd1 vccd1 _08805_/S sky130_fd_sc_hd__nor2_1
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04368_ _16309_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04368_/X sky130_fd_sc_hd__clkbuf_16
X_14309__502 _14310__503/A vssd1 vssd1 vccd1 vccd1 _18137_/CLK sky130_fd_sc_hd__inv_2
XFILLER_225_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _09403_/A vssd1 vssd1 vccd1 vccd1 _19064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09334_ _19093_/Q _08964_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09265_ _18478_/Q vssd1 vssd1 vccd1 vccd1 _09265_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09196_ _19159_/Q _09136_/X _09196_/S vssd1 vssd1 vccd1 vccd1 _09197_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15084__808 _15085__809/A vssd1 vssd1 vccd1 vccd1 _18484_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15422__919 _15422__919/A vssd1 vssd1 vccd1 vccd1 _18606_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _18746_/Q _09955_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__mux2_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14169__447 _14171__449/A vssd1 vssd1 vccd1 vccd1 _18055_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11991_ _11945_/X _11970_/X _11990_/X vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__o21ai_2
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13730_ _13786_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10942_ _10942_/A vssd1 vssd1 vccd1 vccd1 _18302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13661_ _13689_/A vssd1 vssd1 vccd1 vccd1 _13661_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_232_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10873_ _18337_/Q _10794_/X _10879_/S vssd1 vssd1 vccd1 vccd1 _10874_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12612_ _12610_/X _12612_/B _12709_/B vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__and3b_1
XFILLER_188_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _17796_/Q _16383_/A vssd1 vssd1 vccd1 vccd1 _16381_/B sky130_fd_sc_hd__xor2_1
XFILLER_197_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _09250_/A _11826_/A _13541_/A _09252_/B _14069_/B vssd1 vssd1 vccd1 vccd1
+ _13623_/B sky130_fd_sc_hd__a2111o_4
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15331_ _15325_/X _15330_/X _09620_/A vssd1 vssd1 vccd1 vccd1 _15331_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _18004_/Q _12351_/X _12835_/A vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__a21o_1
XFILLER_196_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18050_ _18050_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15262_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _15262_/X sky130_fd_sc_hd__buf_2
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12474_ _12474_/A vssd1 vssd1 vccd1 vccd1 _12547_/S sky130_fd_sc_hd__buf_2
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14213_ _14213_/A vssd1 vssd1 vccd1 vccd1 _18077_/D sky130_fd_sc_hd__clkbuf_1
X_11425_ _11425_/A vssd1 vssd1 vccd1 vccd1 _18105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15193_ _15199_/A vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__buf_1
XFILLER_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11356_ _11356_/A vssd1 vssd1 vccd1 vccd1 _18135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10307_ _10307_/A vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__clkbuf_1
X_14075_ _18007_/Q _14070_/X _14074_/Y _13868_/X vssd1 vssd1 vccd1 vccd1 _18007_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18952_ _18952_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ _18162_/Q _11259_/X _11295_/S vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__mux2_1
X_13026_ _17951_/Q _17687_/Q _13099_/B vssd1 vssd1 vccd1 vccd1 _13027_/B sky130_fd_sc_hd__mux2_1
X_17903_ _17922_/CLK _17903_/D vssd1 vssd1 vccd1 vccd1 _17903_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_opt_3_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _14157_/A
+ sky130_fd_sc_hd__clkbuf_16
X_10238_ _10456_/A _10274_/A vssd1 vssd1 vccd1 vccd1 _10254_/S sky130_fd_sc_hd__nor2_2
X_18883_ _18886_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _17878_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17834_ _18482_/CLK _17834_/D vssd1 vssd1 vccd1 vccd1 _17834_/Q sky130_fd_sc_hd__dfxtp_1
X_10169_ _18697_/Q _10066_/X _10173_/S vssd1 vssd1 vccd1 vccd1 _10170_/A sky130_fd_sc_hd__mux2_1
X_17765_ _19290_/CLK _17765_/D vssd1 vssd1 vccd1 vccd1 _17765_/Q sky130_fd_sc_hd__dfxtp_1
X_14977_ _15059_/A _14977_/B vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__nor2_1
XFILLER_130_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ _13434_/X _13925_/X _13927_/Y _13636_/X vssd1 vssd1 vccd1 vccd1 _17952_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17696_ _17951_/CLK _17696_/D vssd1 vssd1 vccd1 vccd1 _17696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13859_ input69/X _13867_/B vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__and2_1
XFILLER_63_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16578_ _16578_/A _16578_/B _16578_/C vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__nor3_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15529_ _17828_/Q _15529_/B vssd1 vssd1 vccd1 vccd1 _15530_/B sky130_fd_sc_hd__or2_1
X_18317_ _18317_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
X_19297_ _19297_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304__498 _14305__499/A vssd1 vssd1 vccd1 vccd1 _18133_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ _18662_/Q vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__buf_2
XFILLER_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _18248_/CLK _18248_/D vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_opt_12_0_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_82_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_148_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ _18179_/CLK _18179_/D vssd1 vssd1 vccd1 vccd1 _18179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09952_ _18779_/Q _09951_/X _09956_/S vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03799_ _15416_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03799_/X sky130_fd_sc_hd__clkbuf_16
X_15871__167 _15872__168/A vssd1 vssd1 vccd1 vccd1 _18842_/CLK sky130_fd_sc_hd__inv_2
X_08903_ _19302_/Q _08798_/X _08907_/S vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _11024_/A _09892_/B _09882_/X _09870_/X vssd1 vssd1 vccd1 vccd1 _18806_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _09358_/B _09770_/B _09770_/A vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__or3b_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08765_ _18931_/Q hold14/A vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15768__1050 _15772__1054/A vssd1 vssd1 vccd1 vccd1 _18767_/CLK sky130_fd_sc_hd__inv_2
XFILLER_246_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03590_ clkbuf_0__03590_/X vssd1 vssd1 vccd1 vccd1 _15111__829/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09317_ _09317_/A vssd1 vssd1 vccd1 vccd1 _19101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09248_ _09231_/X _10403_/A _09247_/X vssd1 vssd1 vccd1 vccd1 _09971_/C sky130_fd_sc_hd__o21bai_4
XFILLER_167_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09179_ _09179_/A vssd1 vssd1 vccd1 vccd1 _19167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11210_ _18192_/Q _11050_/X _11214_/S vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__mux2_1
X_12190_ _17524_/Q _17487_/B vssd1 vssd1 vccd1 vccd1 _12190_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11141_ _11141_/A vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11072_ _11072_/A vssd1 vssd1 vccd1 vccd1 _18250_/D sky130_fd_sc_hd__clkbuf_1
Xoutput88 _11757_/X vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__buf_2
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput99 _11868_/X vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__buf_2
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _17853_/Q _17852_/Q _14930_/A vssd1 vssd1 vccd1 vccd1 _14938_/A sky130_fd_sc_hd__or3_2
X_10023_ _10023_/A vssd1 vssd1 vccd1 vccd1 _18754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15880_ _15880_/A vssd1 vssd1 vccd1 vccd1 _15880_/X sky130_fd_sc_hd__buf_1
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _18027_/CLK _17550_/D vssd1 vssd1 vccd1 vccd1 _17550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11974_ _19235_/Q _17179_/B _19237_/Q _17186_/B _11961_/X _11977_/S vssd1 vssd1 vccd1
+ vccd1 _11974_/X sky130_fd_sc_hd__mux4_2
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16501_ _16429_/Y _16498_/C _18983_/Q vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__a21oi_1
XFILLER_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13713_ _17881_/Q _13709_/B _13712_/Y _13710_/X vssd1 vssd1 vccd1 vccd1 _17881_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _19339_/Q _12185_/A _12204_/A _19331_/Q vssd1 vssd1 vccd1 vccd1 _17481_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _18309_/Q _10904_/X _10929_/S vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14693_ _19153_/Q _18418_/Q _18312_/Q _18296_/Q _14563_/X _14564_/X vssd1 vssd1 vccd1
+ vccd1 _14694_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19220_ _19281_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_1
X_16432_ _16475_/A vssd1 vssd1 vccd1 vccd1 _16440_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13644_ _13644_/A vssd1 vssd1 vccd1 vccd1 _17859_/D sky130_fd_sc_hd__clkbuf_1
X_14143__428 _14144__429/A vssd1 vssd1 vccd1 vccd1 _18036_/CLK sky130_fd_sc_hd__inv_2
X_10856_ _10856_/A vssd1 vssd1 vccd1 vccd1 _18345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19151_ _19151_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16469_/A vssd1 vssd1 vccd1 vccd1 _16464_/A sky130_fd_sc_hd__clkbuf_2
X_13575_ _16061_/A _13574_/B _13574_/Y _13569_/X vssd1 vssd1 vccd1 vccd1 _17836_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_73_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ _18371_/Q _10713_/X _10787_/S vssd1 vssd1 vccd1 vccd1 _10788_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18102_ _18102_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__04840_ _17019_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04840_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _15306_/X _15313_/X _09615_/A vssd1 vssd1 vccd1 vccd1 _15314_/X sky130_fd_sc_hd__o21a_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _18007_/Q _12511_/X _12924_/A _12525_/X vssd1 vssd1 vccd1 vccd1 _12526_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19082_ _19082_/CLK _19082_/D vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16294_ _18852_/Q _16294_/B _16294_/C _17809_/Q vssd1 vssd1 vccd1 vccd1 _16295_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18033_ _18033_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _15273_/A vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__clkbuf_2
X_12457_ _12727_/A _17627_/Q _12737_/B _12737_/A _12396_/X _12397_/X vssd1 vssd1 vccd1
+ vccd1 _12457_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11408_ _11329_/X _18112_/Q _11412_/S vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__07490_ _12223_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07490_/X sky130_fd_sc_hd__clkbuf_16
X_15176_ _13596_/Y _09971_/C _11816_/X vssd1 vssd1 vccd1 vccd1 _15177_/B sky130_fd_sc_hd__o21ai_1
X_12388_ _17604_/Q _12387_/X _12426_/S vssd1 vssd1 vccd1 vccd1 _12388_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _18026_/Q _14114_/X _14126_/Y vssd1 vssd1 vccd1 vccd1 _18026_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11339_ _11338_/X _18141_/Q _11345_/S vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ _13724_/A _14055_/X _14046_/X vssd1 vssd1 vccd1 vccd1 _14058_/Y sky130_fd_sc_hd__a21oi_1
X_18935_ _18935_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13009_ _17677_/Q _12921_/X _12838_/X _17685_/Q _13008_/X vssd1 vssd1 vccd1 vccd1
+ _13010_/D sky130_fd_sc_hd__a221oi_1
XFILLER_122_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18866_ _18889_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17817_ _19339_/CLK _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18797_ _18797_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17748_ _19327_/CLK _17748_/D vssd1 vssd1 vccd1 vccd1 _17748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15154__864 _15154__864/A vssd1 vssd1 vccd1 vccd1 _18540_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17679_ _17963_/CLK _17679_/D vssd1 vssd1 vccd1 vccd1 _17679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15681__980 _15682__981/A vssd1 vssd1 vccd1 vccd1 _18697_/CLK sky130_fd_sc_hd__inv_2
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09102_ _09102_/A vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09033_ _09033_/A vssd1 vssd1 vccd1 vccd1 _19210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14764__704 _14764__704/A vssd1 vssd1 vccd1 vccd1 _18347_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09935_ _10112_/A vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__clkbuf_2
X_17297__74 _17297__74/A vssd1 vssd1 vccd1 vccd1 _19270_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _09860_/X _09866_/B _09895_/C vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__and3b_1
X_15202__887 _15203__888/A vssd1 vssd1 vccd1 vccd1 _18566_/CLK sky130_fd_sc_hd__inv_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08817_ _08817_/A vssd1 vssd1 vccd1 vccd1 _19322_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _09797_/A vssd1 vssd1 vccd1 vccd1 _18833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08995_/A vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_233_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11690_ _19038_/Q _19037_/Q _16614_/B vssd1 vssd1 vccd1 vccd1 _16619_/B sky130_fd_sc_hd__and3_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10641_ _10641_/A vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13360_ _17101_/A _13355_/X _13358_/Y _13359_/X vssd1 vssd1 vccd1 vccd1 _17775_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10572_ _10123_/X _18496_/Q _10574_/S vssd1 vssd1 vccd1 vccd1 _10573_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _17554_/Q _12202_/X _12212_/X _17556_/Q vssd1 vssd1 vccd1 vccd1 _12316_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13291_ _13146_/X _13288_/X _13275_/X vssd1 vssd1 vccd1 vccd1 _13291_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15030_ _18464_/Q _15031_/C _18465_/Q vssd1 vssd1 vccd1 vccd1 _15032_/A sky130_fd_sc_hd__a21oi_1
XFILLER_154_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12242_ _17548_/Q _18029_/Q _12318_/B vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__mux2_1
XFILLER_120_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12173_ _17529_/Q _18031_/Q _12176_/S vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _11204_/B _11124_/B vssd1 vssd1 vccd1 vccd1 _11140_/S sky130_fd_sc_hd__nor2_2
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16981_ _18250_/Q _18242_/Q _18234_/Q _18226_/Q _16799_/X _16801_/X vssd1 vssd1 vccd1
+ vccd1 _16982_/B sky130_fd_sc_hd__mux4_2
XFILLER_231_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18720_ _18720_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15932_ _17821_/Q _15932_/B vssd1 vssd1 vccd1 vccd1 _15933_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11055_ _11055_/A vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _18761_/Q _09959_/X _10010_/S vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18651_ _18654_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _17602_/CLK _17602_/D vssd1 vssd1 vccd1 vccd1 _17602_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17055__44 _17055__44/A vssd1 vssd1 vccd1 vccd1 _19193_/CLK sky130_fd_sc_hd__inv_2
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _18582_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17533_/CLK _17533_/D vssd1 vssd1 vccd1 vccd1 _17533_/Q sky130_fd_sc_hd__dfxtp_1
X_14745_ _15447_/A vssd1 vssd1 vccd1 vccd1 _14745_/X sky130_fd_sc_hd__buf_1
X_11957_ _11954_/X _11956_/X _11957_/S vssd1 vssd1 vccd1 vccd1 _11957_/X sky130_fd_sc_hd__mux2_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17464_ _17464_/A vssd1 vssd1 vccd1 vccd1 _19335_/D sky130_fd_sc_hd__clkbuf_1
X_10908_ _18316_/Q _10907_/X _10911_/S vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__mux2_1
X_14676_ _19079_/Q _18343_/Q _17577_/Q _18795_/Q _14568_/X _14580_/X vssd1 vssd1 vccd1
+ vccd1 _14677_/B sky130_fd_sc_hd__mux4_2
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ _12245_/A vssd1 vssd1 vccd1 vccd1 _11888_/X sky130_fd_sc_hd__buf_4
XFILLER_232_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19203_ _19203_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
X_16415_ _18972_/Q vssd1 vssd1 vccd1 vccd1 _16453_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13627_ _13173_/X _13626_/B _13626_/Y _13619_/X vssd1 vssd1 vccd1 vccd1 _17853_/D
+ sky130_fd_sc_hd__a211oi_1
X_15822__128 _15823__129/A vssd1 vssd1 vccd1 vccd1 _18803_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10839_ _18352_/Q _10797_/X _10843_/S vssd1 vssd1 vccd1 vccd1 _10840_/A sky130_fd_sc_hd__mux2_1
X_19134_ _19135_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13558_ _13140_/X _13549_/X _13557_/Y _13555_/X vssd1 vssd1 vccd1 vccd1 _17830_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12509_ _12772_/C vssd1 vssd1 vccd1 vccd1 _12920_/A sky130_fd_sc_hd__buf_2
X_19065_ _19065_/CLK _19065_/D vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ _18600_/Q _18616_/Q _18742_/Q _18523_/Q _16195_/X _16112_/X vssd1 vssd1 vccd1
+ vccd1 _16278_/B sky130_fd_sc_hd__mux4_1
X_13489_ _13520_/A _13541_/A _14069_/B vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__or3_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18016_ _18021_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
X_15228_ _15228_/A _15307_/A vssd1 vssd1 vccd1 vccd1 _15228_/X sky130_fd_sc_hd__or2b_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04585_ clkbuf_0__04585_/X vssd1 vssd1 vccd1 vccd1 _16697__321/A sky130_fd_sc_hd__clkbuf_16
X_14416__588 _14417__589/A vssd1 vssd1 vccd1 vccd1 _18223_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09720_ _09742_/S vssd1 vssd1 vccd1 vccd1 _09733_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_113_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18918_ _18919_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16640__280 _16643__283/A vssd1 vssd1 vccd1 vccd1 _19054_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_opt_1_1_wb_clk_i clkbuf_opt_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _10049_/A vssd1 vssd1 vccd1 vccd1 _09975_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_228_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18849_ _18849_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03398_ clkbuf_0__03398_/X vssd1 vssd1 vccd1 vccd1 _14757__698/A sky130_fd_sc_hd__clkbuf_16
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _09597_/S vssd1 vssd1 vccd1 vccd1 _09591_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_227_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__04019_ clkbuf_0__04019_/X vssd1 vssd1 vccd1 vccd1 _15895__184/A sky130_fd_sc_hd__clkbuf_16
XFILLER_211_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_223_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16682__314 _16682__314/A vssd1 vssd1 vccd1 vccd1 _19088_/CLK sky130_fd_sc_hd__inv_2
X_09016_ _09009_/X _09016_/B _09016_/C _09016_/D vssd1 vssd1 vccd1 vccd1 _09016_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_145_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16346__239 _16346__239/A vssd1 vssd1 vccd1 vccd1 _18955_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09918_ _18790_/Q _09223_/X _09926_/S vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ _16826_/A vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _12860_/A _12860_/B _12860_/C _12860_/D vssd1 vssd1 vccd1 vccd1 _12860_/X
+ sky130_fd_sc_hd__or4_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _17932_/Q _11785_/X _11800_/X _11810_/X vssd1 vssd1 vccd1 vccd1 _11811_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688__986 _15689__987/A vssd1 vssd1 vccd1 vccd1 _18703_/CLK sky130_fd_sc_hd__inv_2
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12831_/S vssd1 vssd1 vccd1 vccd1 _12805_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14530_ _14536_/A vssd1 vssd1 vccd1 vccd1 _14530_/X sky130_fd_sc_hd__buf_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11742_ _17916_/Q _11742_/B vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__and2_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14521__672 _14523__674/A vssd1 vssd1 vccd1 vccd1 _18307_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ input4/X vssd1 vssd1 vccd1 vccd1 _11772_/A sky130_fd_sc_hd__inv_8
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16223_/A _16200_/B vssd1 vssd1 vccd1 vccd1 _16200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_224_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13412_ _13411_/X _13395_/X _13408_/X vssd1 vssd1 vccd1 vccd1 _13412_/Y sky130_fd_sc_hd__a21oi_1
X_17180_ _17180_/A _17186_/D vssd1 vssd1 vccd1 vccd1 _17184_/B sky130_fd_sc_hd__and2_1
X_10624_ _18443_/Q _10117_/A _10630_/S vssd1 vssd1 vccd1 vccd1 _10625_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _18567_/Q vssd1 vssd1 vccd1 vccd1 _16162_/S sky130_fd_sc_hd__buf_2
X_13343_ _16584_/A vssd1 vssd1 vccd1 vccd1 _13343_/X sky130_fd_sc_hd__clkbuf_4
X_10555_ _10555_/A vssd1 vssd1 vccd1 vccd1 _18504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12324__388 _12325__389/A vssd1 vssd1 vccd1 vccd1 _17569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _15958_/B _16049_/C _16063_/A _15207_/A vssd1 vssd1 vccd1 vccd1 _16064_/B
+ sky130_fd_sc_hd__a211o_1
X_13274_ _13815_/A vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10486_ _18534_/Q _10345_/X _10490_/S vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15013_ _15013_/A vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ _12176_/S vssd1 vssd1 vccd1 vccd1 _12170_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_123_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__04370_ clkbuf_0__04370_/X vssd1 vssd1 vccd1 vccd1 _16323__221/A sky130_fd_sc_hd__clkbuf_16
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03421_ _14871_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03421_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_150_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _11122_/S vssd1 vssd1 vccd1 vccd1 _11116_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_231_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12087_ _12085_/X _12086_/X _12087_/S vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16964_ _18209_/Q _18129_/Q _19186_/Q _18257_/Q _16822_/X _16823_/X vssd1 vssd1 vccd1
+ vccd1 _16965_/B sky130_fd_sc_hd__mux4_1
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18703_ _18703_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_1
X_15915_ _18867_/Q _15915_/B vssd1 vssd1 vccd1 vccd1 _15935_/A sky130_fd_sc_hd__xnor2_1
X_11038_ _18260_/Q _09142_/X _11040_/S vssd1 vssd1 vccd1 vccd1 _11039_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16895_ _18118_/Q _18110_/Q _18102_/Q _18094_/Q _16893_/X _16894_/X vssd1 vssd1 vccd1
+ vccd1 _16895_/X sky130_fd_sc_hd__mux4_1
X_17028__22 _17028__22/A vssd1 vssd1 vccd1 vccd1 _19171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_237_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _18634_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03183_ clkbuf_0__03183_/X vssd1 vssd1 vccd1 vccd1 _14451__615/A sky130_fd_sc_hd__clkbuf_16
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18565_ _18565_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_2
X_12989_ _17955_/Q _17682_/Q _12993_/S vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__mux2_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ _17737_/CLK _17516_/D vssd1 vssd1 vccd1 vccd1 _17516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14728_ _18860_/Q _18354_/Q _19195_/Q _18362_/Q _14553_/X _14554_/X vssd1 vssd1 vccd1
+ vccd1 _14728_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18496_ _18496_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17447_ _17447_/A vssd1 vssd1 vccd1 vccd1 _19330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14659_ _14657_/X _14658_/X _14729_/S vssd1 vssd1 vccd1 vccd1 _14659_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14422__592 _14423__593/A vssd1 vssd1 vccd1 vccd1 _18227_/CLK sky130_fd_sc_hd__inv_2
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17378_ _17378_/A _17378_/B _17378_/C _17378_/D vssd1 vssd1 vccd1 vccd1 _17378_/X
+ sky130_fd_sc_hd__and4_1
X_14834__760 _14835__761/A vssd1 vssd1 vccd1 vccd1 _18403_/CLK sky130_fd_sc_hd__inv_2
XFILLER_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19117_ _19117_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _19048_/CLK _19048_/D vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__04568_ clkbuf_0__04568_/X vssd1 vssd1 vccd1 vccd1 _16631__273/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_7 _09679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03619_ _15193_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03619_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09703_/A vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14464__626 _14467__629/A vssd1 vssd1 vccd1 vccd1 _18261_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09634_ _09634_/A vssd1 vssd1 vccd1 vccd1 _18930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09565_ _09565_/A vssd1 vssd1 vccd1 vccd1 _18950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03410_ clkbuf_0__03410_/X vssd1 vssd1 vccd1 vccd1 _14820__749/A sky130_fd_sc_hd__clkbuf_16
X_09496_ _19008_/Q _09495_/X _09496_/S vssd1 vssd1 vccd1 vccd1 _09497_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15167__874 _15167__874/A vssd1 vssd1 vccd1 vccd1 _18550_/CLK sky130_fd_sc_hd__inv_2
X_10340_ _18597_/Q _10339_/X _10343_/S vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _10271_/A vssd1 vssd1 vccd1 vccd1 _18626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12003_/X _12009_/X _12022_/A vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15694__990 _15696__992/A vssd1 vssd1 vccd1 vccd1 _18707_/CLK sky130_fd_sc_hd__inv_2
XFILLER_155_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ _16056_/A _13950_/B _13960_/Y _13951_/X vssd1 vssd1 vccd1 vccd1 _17965_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_24_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12912_ _17969_/Q _17667_/Q _12915_/S vssd1 vssd1 vccd1 vccd1 _12913_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _13892_/A vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__buf_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12843_ _12843_/A _12843_/B _12842_/X vssd1 vssd1 vccd1 vccd1 _12860_/A sky130_fd_sc_hd__or3b_1
X_15631_ _16915_/A _15642_/B _15630_/Y _15616_/A _18660_/Q vssd1 vssd1 vccd1 vccd1
+ _18660_/D sky130_fd_sc_hd__a32o_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ _18647_/Q _18646_/Q _15562_/C vssd1 vssd1 vccd1 vccd1 _15572_/C sky130_fd_sc_hd__and3_1
X_18350_ _18350_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
X_12330__392 _12332__394/A vssd1 vssd1 vccd1 vccd1 _17573_/CLK sky130_fd_sc_hd__inv_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12470_/A _12845_/A _12774_/C _12774_/D vssd1 vssd1 vccd1 vccd1 _12775_/C
+ sky130_fd_sc_hd__and4b_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_48_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18021_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11725_ _11717_/X _17931_/Q vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__and2b_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _17834_/Q _15501_/A _17833_/Q vssd1 vssd1 vccd1 vccd1 _15494_/C sky130_fd_sc_hd__o21ai_1
X_18281_ _18281_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17232_ _17237_/C _17233_/C _17231_/Y vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__a21oi_1
XFILLER_187_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03970_ _15692_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03970_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11656_ _11671_/S vssd1 vssd1 vccd1 vccd1 _11665_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17163_ _17173_/D vssd1 vssd1 vccd1 vccd1 _17169_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10607_ _10607_/A vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11587_ _17579_/Q _10695_/A _11593_/S vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14259__462 _14260__463/A vssd1 vssd1 vccd1 vccd1 _18097_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16114_ _16223_/A _16114_/B vssd1 vssd1 vccd1 vccd1 _16114_/Y sky130_fd_sc_hd__nor2_1
X_13326_ _13645_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _14053_/B sky130_fd_sc_hd__nor2_2
X_17094_ _13361_/X _12204_/A _12212_/A _17093_/X _12121_/D vssd1 vssd1 vccd1 vccd1
+ _17094_/X sky130_fd_sc_hd__o2111a_1
X_10538_ _18511_/Q _10342_/X _10538_/S vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16045_ _16044_/A _16044_/B _16049_/A _16063_/A vssd1 vssd1 vccd1 vccd1 _16045_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _13256_/X _13253_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _13257_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10469_ _10469_/A vssd1 vssd1 vccd1 vccd1 _18542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12208_ _17530_/Q _12185_/A _12204_/A _17522_/Q vssd1 vssd1 vccd1 vccd1 _12208_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13188_ _13170_/X _13184_/X _13186_/Y _13187_/X vssd1 vssd1 vccd1 vccd1 _17731_/D
+ sky130_fd_sc_hd__a211oi_1
X_12139_ _12176_/S vssd1 vssd1 vccd1 vccd1 _12153_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17996_ _18014_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03404_ _14784_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03404_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__07172_ _11883_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07172_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16947_ _18184_/Q _18176_/Q _18168_/Q _18160_/Q _16881_/X _16882_/X vssd1 vssd1 vccd1
+ vccd1 _16948_/B sky130_fd_sc_hd__mux4_2
XFILLER_81_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14528__678 _14529__679/A vssd1 vssd1 vccd1 vccd1 _18313_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16878_ _16963_/A _16878_/B vssd1 vssd1 vccd1 vccd1 _16878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18617_ _18617_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03166_ clkbuf_0__03166_/X vssd1 vssd1 vccd1 vccd1 _14370__551/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09350_ _19086_/Q _09271_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _09351_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03197_ _14524_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03197_/X sky130_fd_sc_hd__clkbuf_16
X_18548_ _18548_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03097_ clkbuf_0__03097_/X vssd1 vssd1 vccd1 vccd1 _14173__450/A sky130_fd_sc_hd__clkbuf_16
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09281_ _19120_/Q _09280_/X _09281_/S vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18479_ _15785_/A _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835__138 _15836__139/A vssd1 vssd1 vccd1 vccd1 _18813_/CLK sky130_fd_sc_hd__inv_2
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08996_ _18077_/Q vssd1 vssd1 vccd1 vccd1 _13540_/B sky130_fd_sc_hd__inv_2
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16085__199 _16085__199/A vssd1 vssd1 vccd1 vccd1 _18904_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09617_ _09600_/X _09615_/X _09616_/X vssd1 vssd1 vccd1 vccd1 _09617_/Y sky130_fd_sc_hd__a21boi_1
X_14429__598 _14430__599/A vssd1 vssd1 vccd1 vccd1 _18233_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09548_ _08917_/X _18957_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17022__17 _17022__17/A vssd1 vssd1 vccd1 vccd1 _19166_/CLK sky130_fd_sc_hd__inv_2
XFILLER_212_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09479_ _09148_/B _08860_/A _09477_/C vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__o21ai_1
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16653__290 _16655__292/A vssd1 vssd1 vccd1 vccd1 _19064_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__04373_ clkbuf_0__04373_/X vssd1 vssd1 vccd1 vccd1 _16549_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_200_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11510_/A vssd1 vssd1 vccd1 vccd1 _18040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12490_ _18009_/Q vssd1 vssd1 vccd1 vccd1 _12538_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11441_ _11441_/A vssd1 vssd1 vccd1 vccd1 _18098_/D sky130_fd_sc_hd__clkbuf_1
X_14160_ _14166_/A vssd1 vssd1 vccd1 vccd1 _14160_/X sky130_fd_sc_hd__buf_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11372_ _11372_/A vssd1 vssd1 vccd1 vccd1 _18128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03186_ clkbuf_0__03186_/X vssd1 vssd1 vccd1 vccd1 _14473__634/A sky130_fd_sc_hd__clkbuf_16
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10323_ _10323_/A vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__clkbuf_1
X_14091_ _14099_/A vssd1 vssd1 vccd1 vccd1 _14091_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13042_ _13042_/A vssd1 vssd1 vccd1 vccd1 _17691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10254_ _18633_/Q _10198_/X _10254_/S vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17850_ _17850_/CLK _17850_/D vssd1 vssd1 vccd1 vccd1 _17850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10185_ _10185_/A vssd1 vssd1 vccd1 vccd1 _18692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16801_ _16894_/A vssd1 vssd1 vccd1 vccd1 _16801_/X sky130_fd_sc_hd__buf_4
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17781_ _19281_/CLK _17781_/D vssd1 vssd1 vccd1 vccd1 _17781_/Q sky130_fd_sc_hd__dfxtp_1
X_14993_ _15026_/A vssd1 vssd1 vccd1 vccd1 _14993_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13944_ _13165_/X _13929_/B _13943_/Y _13937_/X vssd1 vssd1 vccd1 vccd1 _17959_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_207_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _13923_/B vssd1 vssd1 vccd1 vccd1 _14053_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_235_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18402_ _18402_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12826_ _12812_/X _12826_/B vssd1 vssd1 vccd1 vccd1 _12827_/A sky130_fd_sc_hd__and2b_1
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15614_ _15615_/B _15615_/C _18657_/Q vssd1 vssd1 vccd1 vccd1 _15616_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16594_ _19025_/Q _16593_/C _19026_/Q vssd1 vssd1 vccd1 vccd1 _16595_/C sky130_fd_sc_hd__a21oi_1
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18333_ _18333_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12757_ _12758_/B _17633_/Q _12747_/A _17635_/Q vssd1 vssd1 vccd1 vccd1 _12759_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_199_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15545_ _15551_/A _15557_/C _15545_/C vssd1 vssd1 vccd1 vccd1 _15545_/X sky130_fd_sc_hd__or3_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A vssd1 vssd1 vccd1 vccd1 _11708_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15476_ _17834_/Q _17833_/Q _15501_/A vssd1 vssd1 vccd1 vccd1 _15494_/B sky130_fd_sc_hd__or3_1
X_18264_ _18264_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
X_12688_ _12686_/B _12687_/A _17614_/Q vssd1 vssd1 vccd1 vccd1 _12689_/C sky130_fd_sc_hd__a21o_1
XFILLER_187_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17215_ _17216_/B _17210_/X _17214_/Y vssd1 vssd1 vccd1 vccd1 _19246_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _08724_/X _17539_/Q _11647_/S vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18195_ _18195_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17146_ _11978_/X _17142_/X _17126_/X vssd1 vssd1 vccd1 vccd1 _17146_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ _13256_/X _13304_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _13309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ _15963_/X _16031_/B _18874_/Q _16025_/B vssd1 vssd1 vccd1 vccd1 _16028_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ _19047_/Q hold20/A vssd1 vssd1 vccd1 vccd1 _09441_/C sky130_fd_sc_hd__xor2_1
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _10219_/A _10219_/B _10219_/C vssd1 vssd1 vccd1 vccd1 _10310_/A sky130_fd_sc_hd__or3_4
XFILLER_245_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17979_ _18001_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
X_12337__398 _12338__399/A vssd1 vssd1 vccd1 vccd1 _17579_/CLK sky130_fd_sc_hd__inv_2
XFILLER_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04367_ _16308_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04367_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09402_ _08921_/X _19064_/Q _09406_/S vssd1 vssd1 vccd1 vccd1 _09403_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03149_ clkbuf_0__03149_/X vssd1 vssd1 vccd1 vccd1 _14284__482/A sky130_fd_sc_hd__clkbuf_16
XFILLER_240_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09333_ _09333_/A vssd1 vssd1 vccd1 vccd1 _19094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _09264_/A vssd1 vssd1 vccd1 vccd1 _19126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09195_ _09195_/A vssd1 vssd1 vccd1 vccd1 _19160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14847__770 _14850__773/A vssd1 vssd1 vccd1 vccd1 _18415_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_248_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08979_ _08979_/A vssd1 vssd1 vccd1 vccd1 _19217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _12020_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11990_/X sky130_fd_sc_hd__or2_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _18302_/Q _10901_/X _10941_/S vssd1 vssd1 vccd1 vccd1 _10942_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13660_ _13666_/A vssd1 vssd1 vccd1 vccd1 _13660_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_231_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _10872_/A vssd1 vssd1 vccd1 vccd1 _18338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12611_ _12610_/B _12610_/C _12610_/A vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__a21o_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13591_/A vssd1 vssd1 vccd1 vccd1 _17842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15307_/X _15326_/X _15329_/Y vssd1 vssd1 vccd1 vccd1 _15330_/X sky130_fd_sc_hd__o21a_2
X_12542_ _12774_/C vssd1 vssd1 vccd1 vccd1 _12835_/A sky130_fd_sc_hd__buf_2
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _18829_/Q _18821_/Q _18813_/Q _18680_/Q _15214_/X _15225_/X vssd1 vssd1 vccd1
+ vccd1 _15261_/X sky130_fd_sc_hd__mux4_1
X_12473_ _12727_/C _12727_/B _12727_/A _17627_/Q _12366_/X _12368_/X vssd1 vssd1 vccd1
+ vccd1 _12473_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ _09250_/A input35/X _14218_/S vssd1 vssd1 vccd1 vccd1 _14213_/A sky130_fd_sc_hd__mux2_1
X_17000_ _17000_/A vssd1 vssd1 vccd1 vccd1 _17000_/X sky130_fd_sc_hd__buf_1
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11424_ _18105_/Q _11264_/X _11430_/S vssd1 vssd1 vccd1 vccd1 _11425_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _15535_/A _15190_/B _16915_/A _15191_/X vssd1 vssd1 vccd1 vccd1 _18558_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11355_ _18135_/Q _11270_/X _11357_/S vssd1 vssd1 vccd1 vccd1 _11356_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03169_ clkbuf_0__03169_/X vssd1 vssd1 vccd1 vccd1 _14511_/A sky130_fd_sc_hd__clkbuf_16
X_10306_ _18610_/Q _10195_/X _10308_/S vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__mux2_1
X_14074_ _14074_/A _14083_/B vssd1 vssd1 vccd1 vccd1 _14074_/Y sky130_fd_sc_hd__nor2_1
X_18951_ _18951_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _11301_/S vssd1 vssd1 vccd1 vccd1 _11295_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ _13076_/S vssd1 vssd1 vccd1 vccd1 _13099_/B sky130_fd_sc_hd__clkbuf_2
X_17902_ _17922_/CLK _17902_/D vssd1 vssd1 vccd1 vccd1 _17902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _10237_/A vssd1 vssd1 vccd1 vccd1 _18671_/D sky130_fd_sc_hd__clkbuf_1
X_18882_ _18886_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748__690 _14749__691/A vssd1 vssd1 vccd1 vccd1 _18333_/CLK sky130_fd_sc_hd__inv_2
X_17833_ _18482_/CLK _17833_/D vssd1 vssd1 vccd1 vccd1 _17833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _10168_/A vssd1 vssd1 vccd1 vccd1 _18698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17764_ _19288_/CLK _17764_/D vssd1 vssd1 vccd1 vccd1 _17764_/Q sky130_fd_sc_hd__dfxtp_1
X_14976_ _14973_/Y _14975_/X _18455_/Q vssd1 vssd1 vccd1 vccd1 _14977_/B sky130_fd_sc_hd__mux2_1
X_10099_ _10099_/A vssd1 vssd1 vccd1 vccd1 _18725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_63_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _17945_/CLK sky130_fd_sc_hd__clkbuf_16
X_16715_ _19109_/Q _16715_/B _19111_/Q vssd1 vssd1 vccd1 vccd1 _19111_/D sky130_fd_sc_hd__nor3b_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13927_ _17952_/Q _13929_/B vssd1 vssd1 vccd1 vccd1 _13927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_207_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17695_ _17703_/CLK _17695_/D vssd1 vssd1 vccd1 vccd1 _17695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16646_ _16658_/A vssd1 vssd1 vccd1 vccd1 _16646_/X sky130_fd_sc_hd__buf_1
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13858_ _17929_/Q _13850_/X _13856_/X _13857_/X vssd1 vssd1 vccd1 vccd1 _17929_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _17645_/Q _17990_/Q _12822_/S vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__mux2_1
XFILLER_204_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16577_ _19019_/Q _16576_/C _19020_/Q vssd1 vssd1 vccd1 vccd1 _16578_/C sky130_fd_sc_hd__a21oi_1
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13789_ _13880_/A vssd1 vssd1 vccd1 vccd1 _13789_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18316_ _18316_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
X_15528_ _15528_/A _15528_/B _15528_/C _15528_/D vssd1 vssd1 vccd1 vccd1 _15528_/X
+ sky130_fd_sc_hd__or4_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19296_ _19296_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18247_ _18247_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ _18178_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _17129_/A _17129_/B _17129_/C vssd1 vssd1 vccd1 vccd1 _17135_/B sky130_fd_sc_hd__and3_1
XFILLER_190_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ _10123_/A vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__03798_ _15410_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03798_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ _08902_/A vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__clkbuf_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _11383_/A _09011_/A _09894_/B _09025_/A vssd1 vssd1 vccd1 vccd1 _09882_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ hold15/X vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _18925_/Q _18930_/Q vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__and2b_1
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15090__813 _15091__814/A vssd1 vssd1 vccd1 vccd1 _18489_/CLK sky130_fd_sc_hd__inv_2
XFILLER_241_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09316_ _08937_/X _19101_/Q _09318_/S vssd1 vssd1 vccd1 vccd1 _09317_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _09247_/A _09247_/B _09247_/C _09247_/D vssd1 vssd1 vccd1 vccd1 _09247_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_31_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _19167_/Q _09104_/X _09178_/S vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14175__452 _14177__454/A vssd1 vssd1 vccd1 vccd1 _18060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11140_ _18219_/Q _11065_/X _11140_/S vssd1 vssd1 vccd1 vccd1 _11141_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11071_ _08991_/X _18250_/Q _11079_/S vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__mux2_1
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput89 _11753_/X vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__buf_2
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10022_ _18754_/Q _09955_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11973_ _19238_/Q vssd1 vssd1 vccd1 vccd1 _17186_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _16498_/X _16499_/Y _16469_/A vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__a21oi_1
X_13712_ _13712_/A _13712_/B vssd1 vssd1 vccd1 vccd1 _13712_/Y sky130_fd_sc_hd__nor2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ _10924_/A vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__clkbuf_1
X_17480_ _19335_/Q _12199_/X _12187_/X _19325_/Q vssd1 vssd1 vccd1 vccd1 _17485_/C
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14692_ _14688_/X _14691_/X _14730_/S vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__mux2_2
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16733__346 _16999__349/A vssd1 vssd1 vccd1 vccd1 _19125_/CLK sky130_fd_sc_hd__inv_2
X_16431_ _16464_/A _16431_/B vssd1 vssd1 vccd1 vccd1 _18968_/D sky130_fd_sc_hd__nor2_1
X_13643_ _13710_/A _13643_/B vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__or2_1
X_10855_ _18345_/Q _10794_/X _10861_/S vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19150_ _19150_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13574_ _17836_/Q _13574_/B vssd1 vssd1 vccd1 vccd1 _13574_/Y sky130_fd_sc_hd__nor2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _16362_/A vssd1 vssd1 vccd1 vccd1 _16469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10786_ _10786_/A vssd1 vssd1 vccd1 vccd1 _18372_/D sky130_fd_sc_hd__clkbuf_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _18101_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12574_/B _12511_/X _12524_/X vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__a21bo_1
X_15313_ _15307_/X _15309_/X _15312_/Y vssd1 vssd1 vccd1 vccd1 _15313_/X sky130_fd_sc_hd__o21a_2
X_16293_ _18921_/Q _16164_/X _16292_/Y _16216_/X vssd1 vssd1 vccd1 vccd1 _18921_/D
+ sky130_fd_sc_hd__o211a_1
X_19081_ _19081_/CLK _19081_/D vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17504__2 _11876_/A vssd1 vssd1 vccd1 vccd1 _19346_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18032_ _18032_/CLK _18032_/D vssd1 vssd1 vccd1 vccd1 _18032_/Q sky130_fd_sc_hd__dfxtp_1
X_12456_ _17629_/Q vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _15244_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _11407_/A vssd1 vssd1 vccd1 vccd1 _18113_/D sky130_fd_sc_hd__clkbuf_1
X_15175_ _15175_/A vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__clkbuf_1
X_12387_ _17605_/Q vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14126_ _13750_/A _14120_/X _14123_/X vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__a21oi_1
X_11338_ _11338_/A vssd1 vssd1 vccd1 vccd1 _11338_/X sky130_fd_sc_hd__buf_2
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14057_ _18000_/Q _14054_/X _14056_/Y vssd1 vssd1 vccd1 vccd1 _18000_/D sky130_fd_sc_hd__o21a_1
XFILLER_140_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18934_ _18934_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_1
X_11269_ _11269_/A vssd1 vssd1 vccd1 vccd1 _18168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13008_ _17680_/Q _13085_/B vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__xor2_1
XFILLER_234_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18865_ _18889_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17816_ _19339_/CLK _17816_/D vssd1 vssd1 vccd1 vccd1 _17816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18796_ _18796_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17747_ _19327_/CLK _17747_/D vssd1 vssd1 vccd1 vccd1 _17747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14959_ _18482_/Q vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__inv_2
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17678_ _17963_/CLK _17678_/D vssd1 vssd1 vccd1 vccd1 _17678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_220 _09223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19348_ _19348_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09101_ _19192_/Q _09100_/X _09105_/S vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19279_ _19281_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09032_ _09031_/X _19210_/Q _09044_/S vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14352__537 _14352__537/A vssd1 vssd1 vccd1 vccd1 _18172_/CLK sky130_fd_sc_hd__inv_2
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15161__869 _15161__869/A vssd1 vssd1 vccd1 vccd1 _18545_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _18480_/Q vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__buf_4
XFILLER_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09865_ _16875_/S _09872_/A vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__or2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08816_ _19322_/Q _08786_/X _08822_/S vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__mux2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09796_ _18833_/Q _09752_/X _09800_/S vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08747_ _18067_/Q _08747_/B _13873_/B vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__nor3_1
XFILLER_172_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10640_ _09223_/X _18436_/Q _10648_/S vssd1 vssd1 vccd1 vccd1 _10641_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10571_ _10571_/A vssd1 vssd1 vccd1 vccd1 _18497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12310_ _17554_/Q _12202_/X _12204_/X _17555_/Q _12309_/X vssd1 vssd1 vccd1 vccd1
+ _12316_/B sky130_fd_sc_hd__o221a_1
XFILLER_194_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13290_ _17755_/Q _13280_/X _13289_/Y vssd1 vssd1 vccd1 vccd1 _17755_/D sky130_fd_sc_hd__o21a_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12241_ _12293_/S vssd1 vssd1 vccd1 vccd1 _12318_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _12172_/A vssd1 vssd1 vccd1 vccd1 _17528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14253__457 _14255__459/A vssd1 vssd1 vccd1 vccd1 _18092_/CLK sky130_fd_sc_hd__inv_2
X_11123_ _11123_/A vssd1 vssd1 vccd1 vccd1 _18227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16980_ _16976_/X _16979_/X _16980_/S vssd1 vssd1 vccd1 vccd1 _16980_/X sky130_fd_sc_hd__mux2_2
XFILLER_104_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15931_ _18864_/Q _15931_/B vssd1 vssd1 vccd1 vccd1 _15931_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11054_ _18255_/Q _11053_/X _11057_/S vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10005_ _10005_/A vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _18654_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15862_ _15880_/A vssd1 vssd1 vccd1 vccd1 _15862_/X sky130_fd_sc_hd__buf_1
XFILLER_236_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17601_ _17602_/CLK _17601_/D vssd1 vssd1 vccd1 vccd1 _17601_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _18581_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _15799_/A vssd1 vssd1 vccd1 vccd1 _15793_/X sky130_fd_sc_hd__buf_1
XFILLER_217_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17532_ _17532_/CLK _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ _17225_/B _19250_/Q _11956_/S vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__mux2_1
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_4_0_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_233_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17463_ _17454_/X _17463_/B vssd1 vssd1 vccd1 vccd1 _17464_/A sky130_fd_sc_hd__and2b_1
X_10907_ _18988_/Q vssd1 vssd1 vccd1 vccd1 _10907_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11887_ _12918_/A vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__clkbuf_2
X_14675_ _14732_/A _14675_/B vssd1 vssd1 vccd1 vccd1 _14675_/Y sky130_fd_sc_hd__nor2_1
XFILLER_233_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19202_ _19202_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16414_ _18972_/Q _16416_/B vssd1 vssd1 vccd1 vccd1 _16417_/C sky130_fd_sc_hd__nor2_1
X_13626_ _17853_/Q _13626_/B vssd1 vssd1 vccd1 vccd1 _13626_/Y sky130_fd_sc_hd__nor2_1
X_10838_ _10838_/A vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19133_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13557_ _17830_/Q _13557_/B vssd1 vssd1 vccd1 vccd1 _13557_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ _10769_/A vssd1 vssd1 vccd1 vccd1 _18379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12508_ _12469_/S _12501_/X _12504_/Y _12507_/Y vssd1 vssd1 vccd1 vccd1 _12772_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_19064_ _19064_/CLK _19064_/D vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfxtp_1
X_16276_ _16276_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16276_/Y sky130_fd_sc_hd__nor2_1
X_13488_ _13488_/A _13540_/B _14186_/D _08741_/D vssd1 vssd1 vccd1 vccd1 _13520_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_185_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18015_ _18021_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
X_12439_ _17605_/Q _17606_/Q _12440_/S vssd1 vssd1 vccd1 vccd1 _12439_/X sky130_fd_sc_hd__mux2_1
X_15227_ _18671_/Q _18577_/Q _17532_/Q _17507_/Q _09605_/A _09631_/A vssd1 vssd1 vccd1
+ vccd1 _15228_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ _13733_/A _14099_/X _14108_/X vssd1 vssd1 vccd1 vccd1 _14109_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18917_ _18919_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09650_ _09650_/A vssd1 vssd1 vccd1 vccd1 _18925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18848_ _18848_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03397_ clkbuf_0__03397_/X vssd1 vssd1 vccd1 vccd1 _14749__691/A sky130_fd_sc_hd__clkbuf_16
XFILLER_228_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ _10220_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09597_/S sky130_fd_sc_hd__nor2_2
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18779_ _18779_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09015_ hold26/A _09880_/B _09856_/C vssd1 vssd1 vccd1 vccd1 _09016_/D sky130_fd_sc_hd__a21o_1
XFILLER_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09917_ _09932_/S vssd1 vssd1 vccd1 vccd1 _09926_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_59_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09848_ _18809_/Q vssd1 vssd1 vccd1 vccd1 _16826_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09779_ _08874_/X _18840_/Q _09781_/S vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__mux2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _17913_/Q _11793_/X _11809_/Y input12/X _11802_/X vssd1 vssd1 vccd1 vccd1
+ _11810_/X sky130_fd_sc_hd__a221o_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A vssd1 vssd1 vccd1 vccd1 _17639_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11741_/A vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11672_/A vssd1 vssd1 vccd1 vccd1 _17507_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13411_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10623_ _10623_/A vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13342_ _13330_/A _17101_/C vssd1 vssd1 vccd1 vccd1 _13342_/X sky130_fd_sc_hd__and2b_1
X_16130_ _16126_/X _16129_/X _16194_/A vssd1 vssd1 vccd1 vccd1 _16130_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _18504_/Q _10123_/A _10556_/S vssd1 vssd1 vccd1 vccd1 _10555_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13273_ _17751_/Q _13253_/X _13272_/Y vssd1 vssd1 vccd1 vccd1 _17751_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ _16061_/A _16061_/B vssd1 vssd1 vccd1 vccd1 _18887_/D sky130_fd_sc_hd__nor2_1
X_10485_ _10485_/A vssd1 vssd1 vccd1 vccd1 _18535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ _15034_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _15013_/A sky130_fd_sc_hd__and2_1
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _12155_/A vssd1 vssd1 vccd1 vccd1 _17523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03420_ _14870_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03420_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11106_ _11260_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11122_/S sky130_fd_sc_hd__nor2_2
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12086_ _19263_/Q _19264_/Q _19265_/Q _19266_/Q _11980_/X _11981_/X vssd1 vssd1 vccd1
+ vccd1 _12086_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16698__322 _16700__324/A vssd1 vssd1 vccd1 vccd1 _19097_/CLK sky130_fd_sc_hd__inv_2
X_16963_ _16963_/A _16963_/B vssd1 vssd1 vccd1 vccd1 _16963_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18702_ _18702_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ _17819_/Q _15917_/B vssd1 vssd1 vccd1 vccd1 _15915_/B sky130_fd_sc_hd__xor2_1
X_11037_ _11037_/A vssd1 vssd1 vccd1 vccd1 _18261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16894_ _16894_/A vssd1 vssd1 vccd1 vccd1 _16894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18633_ _18633_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03182_ clkbuf_0__03182_/X vssd1 vssd1 vccd1 vccd1 _14456_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18564_ _18564_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12988_ _12988_/A vssd1 vssd1 vccd1 vccd1 _17681_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17515_ _17878_/CLK _17515_/D vssd1 vssd1 vccd1 vccd1 _17515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14727_ _18370_/Q _18322_/Q _18378_/Q _17711_/Q _14599_/X _14627_/X vssd1 vssd1 vccd1
+ vccd1 _14727_/X sky130_fd_sc_hd__mux4_1
X_11939_ _11931_/X _11933_/X _11935_/X _11936_/X _12017_/S _11907_/S vssd1 vssd1 vccd1
+ vccd1 _11939_/X sky130_fd_sc_hd__mux4_1
X_18495_ _18495_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17446_ _17437_/X _17446_/B vssd1 vssd1 vccd1 vccd1 _17447_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14658_ _18406_/Q _18398_/Q _19311_/Q _17715_/Q _14580_/A _14615_/X vssd1 vssd1 vccd1
+ vccd1 _14658_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13609_ _13140_/X _13601_/X _13608_/Y _13604_/X vssd1 vssd1 vccd1 vccd1 _17847_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17377_ _17377_/A _17377_/B _17377_/C _17377_/D vssd1 vssd1 vccd1 vccd1 _17378_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_242_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14589_ _14623_/A vssd1 vssd1 vccd1 vccd1 _14589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_229_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19116_ _19116_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19047_ _19047_/CLK _19047_/D vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfxtp_2
X_16259_ _16278_/A _16259_/B vssd1 vssd1 vccd1 vccd1 _16259_/Y sky130_fd_sc_hd__nor2_1
X_14156__439 _14156__439/A vssd1 vssd1 vccd1 vccd1 _18047_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_8 _09688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09702_ _09674_/X _18897_/Q _09710_/S vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14841__765 _14843__767/A vssd1 vssd1 vccd1 vccd1 _18408_/CLK sky130_fd_sc_hd__inv_2
X_09633_ _09626_/B _09633_/B _09649_/C vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__and3b_1
XFILLER_244_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09564_ _18950_/Q _09481_/X _09572_/S vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _18883_/Q vssd1 vssd1 vccd1 vccd1 _09495_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16352__244 _16352__244/A vssd1 vssd1 vccd1 vccd1 _18960_/CLK sky130_fd_sc_hd__inv_2
XFILLER_221_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ _18626_/Q _10195_/X _10272_/S vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13960_ _17965_/Q _13962_/B vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12911_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13891_ _17940_/Q _13878_/X _13890_/Y vssd1 vssd1 vccd1 vccd1 _17940_/D sky130_fd_sc_hd__o21a_1
X_14365__547 _14367__549/A vssd1 vssd1 vccd1 vccd1 _18182_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15630_ _15630_/A _15630_/B vssd1 vssd1 vccd1 vccd1 _15630_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _17639_/Q _12932_/A _13092_/B _17650_/Q _12841_/Y vssd1 vssd1 vccd1 vccd1
+ _12842_/X sky130_fd_sc_hd__o221a_1
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _18647_/Q _15561_/B vssd1 vssd1 vccd1 vccd1 _15563_/B sky130_fd_sc_hd__nor2_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12451_/A _12773_/B _12921_/A _12773_/D vssd1 vssd1 vccd1 vccd1 _12776_/A
+ sky130_fd_sc_hd__and4b_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04587_ clkbuf_0__04587_/X vssd1 vssd1 vccd1 vccd1 _16710__332/A sky130_fd_sc_hd__clkbuf_16
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14524_/A vssd1 vssd1 vccd1 vccd1 _14512_/X sky130_fd_sc_hd__buf_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11724_/A vssd1 vssd1 vccd1 vccd1 _11724_/X sky130_fd_sc_hd__clkbuf_1
X_18280_ _18280_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15492_ _18652_/Q _15492_/B vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__xnor2_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17237_/C _17233_/C _17191_/X vssd1 vssd1 vccd1 vccd1 _17231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11655_ _11655_/A hold2/X vssd1 vssd1 vccd1 vccd1 _11671_/S sky130_fd_sc_hd__nor2_2
X_14443_ _14443_/A vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__buf_1
XFILLER_202_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17162_ _19232_/Q _19231_/Q _19230_/Q _17162_/D vssd1 vssd1 vccd1 vccd1 _17173_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_168_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18921_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10606_ _10117_/X _18451_/Q _10612_/S vssd1 vssd1 vccd1 vccd1 _10607_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11586_ _11586_/A vssd1 vssd1 vccd1 vccd1 _17580_/D sky130_fd_sc_hd__clkbuf_1
X_14374_ _14374_/A vssd1 vssd1 vccd1 vccd1 _14374_/X sky130_fd_sc_hd__buf_1
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16113_ _18437_/Q _18687_/Q _18695_/Q _18703_/Q _16112_/X _10405_/A vssd1 vssd1 vccd1
+ vccd1 _16114_/B sky130_fd_sc_hd__mux4_1
X_13325_ _14053_/A vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19132_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10537_ _10537_/A vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__clkbuf_1
X_17093_ _12202_/A _12203_/A _17092_/X _13346_/B _17101_/A vssd1 vssd1 vccd1 vccd1
+ _17093_/X sky130_fd_sc_hd__a32o_1
XFILLER_155_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15703__998 _15704__999/A vssd1 vssd1 vccd1 vccd1 _18715_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _16044_/A _16044_/B vssd1 vssd1 vccd1 vccd1 _16044_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13256_ _14074_/A vssd1 vssd1 vccd1 vccd1 _13256_/X sky130_fd_sc_hd__buf_4
X_10468_ _18542_/Q _10345_/X _10472_/S vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12207_/A vssd1 vssd1 vccd1 vccd1 _12212_/A sky130_fd_sc_hd__buf_2
XFILLER_142_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13187_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13187_/X sky130_fd_sc_hd__clkbuf_2
X_10399_ _18564_/Q vssd1 vssd1 vccd1 vccd1 _16205_/A sky130_fd_sc_hd__buf_2
XFILLER_215_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12138_ _12138_/A vssd1 vssd1 vccd1 vccd1 _17518_/D sky130_fd_sc_hd__clkbuf_1
X_17995_ _18014_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03403_ _14778_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03403_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__07171_ _11882_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07171_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12069_ _12069_/A _12069_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__or2_1
X_16946_ _16984_/A _16946_/B vssd1 vssd1 vccd1 vccd1 _16946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16877_ _18245_/Q _18237_/Q _18229_/Q _18221_/Q _16849_/X _16850_/X vssd1 vssd1 vccd1
+ vccd1 _16878_/B sky130_fd_sc_hd__mux4_1
XFILLER_226_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18616_ _18616_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14266__467 _14268__469/A vssd1 vssd1 vccd1 vccd1 _18102_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03165_ clkbuf_0__03165_/X vssd1 vssd1 vccd1 vccd1 _14367__549/A sky130_fd_sc_hd__clkbuf_16
XFILLER_93_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17406__97 _17408__99/A vssd1 vssd1 vccd1 vccd1 _19310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03196_ _14518_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03196_/X sky130_fd_sc_hd__clkbuf_16
X_18547_ _18547_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03096_ clkbuf_0__03096_/X vssd1 vssd1 vccd1 vccd1 _14171__449/A sky130_fd_sc_hd__clkbuf_16
XFILLER_205_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09280_ _18473_/Q vssd1 vssd1 vccd1 vccd1 _09280_/X sky130_fd_sc_hd__buf_2
X_18478_ _15785_/A _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17429_ _17356_/X _17429_/B vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__and2b_1
XFILLER_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14470__631 _14473__634/A vssd1 vssd1 vccd1 vccd1 _18266_/CLK sky130_fd_sc_hd__inv_2
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08995_ _08995_/A vssd1 vssd1 vccd1 vccd1 _13645_/B sky130_fd_sc_hd__clkinv_2
XFILLER_214_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _16294_/B vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09547_ _09547_/A vssd1 vssd1 vccd1 vccd1 _18958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09478_ _09478_/A vssd1 vssd1 vccd1 vccd1 _19042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04372_ clkbuf_0__04372_/X vssd1 vssd1 vccd1 vccd1 _16338__234/A sky130_fd_sc_hd__clkbuf_16
XFILLER_240_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ _18098_/Q _11259_/X _11448_/S vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11371_ _11329_/X _18128_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03185_ clkbuf_0__03185_/X vssd1 vssd1 vccd1 vccd1 _14467__629/A sky130_fd_sc_hd__clkbuf_16
X_13110_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13110_/X sky130_fd_sc_hd__buf_1
X_10322_ _09691_/X _18603_/Q _10326_/S vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__mux2_1
X_14090_ _14090_/A _14113_/B _16052_/C vssd1 vssd1 vccd1 vccd1 _14099_/A sky130_fd_sc_hd__and3_2
XFILLER_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _13032_/X _13041_/B vssd1 vssd1 vccd1 vccd1 _13042_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ _10253_/A vssd1 vssd1 vccd1 vccd1 _18634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10184_ _18692_/Q _10183_/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10185_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16800_ _18808_/Q vssd1 vssd1 vccd1 vccd1 _16894_/A sky130_fd_sc_hd__clkbuf_4
X_17780_ _19246_/CLK _17780_/D vssd1 vssd1 vccd1 vccd1 _17780_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14992_ _18458_/Q _14998_/C vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__xor2_1
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16731_ _17006_/A vssd1 vssd1 vccd1 vccd1 _16731_/X sky130_fd_sc_hd__buf_1
X_13943_ _17959_/Q _13943_/B vssd1 vssd1 vccd1 vccd1 _13943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13874_ _13759_/A _13874_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__and3b_1
XFILLER_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ _18401_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
X_15613_ _15611_/X _15612_/Y _15581_/A vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12825_ _17650_/Q _17985_/Q _12831_/S vssd1 vssd1 vccd1 vccd1 _12826_/B sky130_fd_sc_hd__mux2_1
XFILLER_216_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16593_ _19026_/Q _19025_/Q _16593_/C vssd1 vssd1 vccd1 vccd1 _16595_/B sky130_fd_sc_hd__and3_1
XFILLER_90_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18332_ _18332_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15544_ _18643_/Q _15543_/C _18644_/Q vssd1 vssd1 vccd1 vccd1 _15545_/C sky130_fd_sc_hd__a21oi_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ _12756_/A vssd1 vssd1 vccd1 vccd1 _17634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11707_ _17907_/Q _17720_/Q _11707_/S vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__mux2_8
XFILLER_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18263_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15475_ _17835_/Q _15505_/B vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__or2_1
X_12687_ _12687_/A _12694_/D vssd1 vssd1 vccd1 vccd1 _12687_/X sky130_fd_sc_hd__and2_1
XFILLER_203_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17214_ _17216_/B _17210_/X _17112_/B vssd1 vssd1 vccd1 vccd1 _17214_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11638_ _11653_/S vssd1 vssd1 vccd1 vccd1 _11647_/S sky130_fd_sc_hd__clkbuf_2
X_18194_ _18194_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17145_ _17145_/A vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11569_ _17587_/Q _10892_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__mux2_1
X_13308_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13308_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14534__683 _14535__684/A vssd1 vssd1 vccd1 vccd1 _18318_/CLK sky130_fd_sc_hd__inv_2
XFILLER_170_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16027_ _18874_/Q _18873_/Q _16027_/C vssd1 vssd1 vccd1 vccd1 _16031_/B sky130_fd_sc_hd__and3_1
XFILLER_115_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13239_ _17741_/Q _13218_/X _13238_/Y vssd1 vssd1 vccd1 vccd1 _17741_/D sky130_fd_sc_hd__o21a_1
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08780_ _09789_/A vssd1 vssd1 vccd1 vccd1 _10219_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17978_ _18001_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_1
X_15454__944 _15454__944/A vssd1 vssd1 vccd1 vccd1 _18631_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16929_ _16929_/A _16929_/B vssd1 vssd1 vccd1 vccd1 _16929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _09401_/A vssd1 vssd1 vccd1 vccd1 _19065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03148_ clkbuf_0__03148_/X vssd1 vssd1 vccd1 vccd1 _14277__476/A sky130_fd_sc_hd__clkbuf_16
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _19094_/Q _08961_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03179_ _14431_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03179_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _19126_/Q _09262_/X _09272_/S vssd1 vssd1 vccd1 vccd1 _09264_/A sky130_fd_sc_hd__mux2_1
X_15841__143 _15842__144/A vssd1 vssd1 vccd1 vccd1 _18818_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _19160_/Q _09133_/X _09196_/S vssd1 vssd1 vccd1 vccd1 _09195_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14316__508 _14317__509/A vssd1 vssd1 vccd1 vccd1 _18143_/CLK sky130_fd_sc_hd__inv_2
XFILLER_161_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08978_ _19217_/Q _08952_/X _08982_/S vssd1 vssd1 vccd1 vccd1 _08979_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _10940_/A vssd1 vssd1 vccd1 vccd1 _18303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10871_ _18338_/Q _10789_/X _10879_/S vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12610_ _12610_/A _12610_/B _12610_/C vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__and3_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13629_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__or2_1
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12586_/S _12537_/X _12539_/Y _12540_/Y vssd1 vssd1 vccd1 vccd1 _12774_/C
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14477__637 _14479__639/A vssd1 vssd1 vccd1 vccd1 _18272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15260_ _15220_/X _15255_/X _15259_/Y vssd1 vssd1 vccd1 vccd1 _15260_/X sky130_fd_sc_hd__o21a_1
X_12472_ _17625_/Q vssd1 vssd1 vccd1 vccd1 _12727_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _14211_/A vssd1 vssd1 vccd1 vccd1 _18076_/D sky130_fd_sc_hd__clkbuf_1
X_11423_ _11423_/A vssd1 vssd1 vccd1 vccd1 _18106_/D sky130_fd_sc_hd__clkbuf_1
X_15191_ _15182_/Y _15185_/X _15189_/X _15630_/A vssd1 vssd1 vccd1 vccd1 _15191_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11354_ _11354_/A vssd1 vssd1 vccd1 vccd1 _18136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03168_ clkbuf_0__03168_/X vssd1 vssd1 vccd1 vccd1 _14382__561/A sky130_fd_sc_hd__clkbuf_16
X_10305_ _10305_/A vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14073_ _12574_/B _14070_/X _14072_/Y _13868_/X vssd1 vssd1 vccd1 vccd1 _18006_/D
+ sky130_fd_sc_hd__a211o_1
X_11285_ _11511_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11301_/S sky130_fd_sc_hd__nor2_2
X_18950_ _18950_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13024_ _18000_/Q _13024_/B vssd1 vssd1 vccd1 vccd1 _13076_/S sky130_fd_sc_hd__and2_2
X_17901_ _17922_/CLK _17901_/D vssd1 vssd1 vccd1 vccd1 _17901_/Q sky130_fd_sc_hd__dfxtp_1
X_10236_ _18671_/Q _09767_/X hold3/X vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18881_ _18886_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_133_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17832_ _18482_/CLK _17832_/D vssd1 vssd1 vccd1 vccd1 _17832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10167_ _18698_/Q _10063_/X _10167_/S vssd1 vssd1 vccd1 vccd1 _10168_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _19288_/CLK _17763_/D vssd1 vssd1 vccd1 vccd1 _17763_/Q sky130_fd_sc_hd__dfxtp_1
X_14975_ _14979_/C _16097_/B _15076_/B _15080_/C vssd1 vssd1 vccd1 vccd1 _14975_/X
+ sky130_fd_sc_hd__o31a_1
X_10098_ _18725_/Q _10054_/X _10104_/S vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16714_ _19109_/Q _16715_/B _19110_/Q vssd1 vssd1 vccd1 vccd1 _19110_/D sky130_fd_sc_hd__nor3b_1
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13926_ _13943_/B vssd1 vssd1 vccd1 vccd1 _13929_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17694_ _17703_/CLK _17694_/D vssd1 vssd1 vccd1 vccd1 _17694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ _16718_/A vssd1 vssd1 vccd1 vccd1 _16645_/X sky130_fd_sc_hd__buf_1
X_13857_ _16584_/A vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12808_ _12831_/S vssd1 vssd1 vccd1 vccd1 _12822_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16576_ _19020_/Q _19019_/Q _16576_/C vssd1 vssd1 vccd1 vccd1 _16578_/B sky130_fd_sc_hd__and3_1
XFILLER_188_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13788_ _17906_/Q _13771_/X _13787_/Y vssd1 vssd1 vccd1 vccd1 _17906_/D sky130_fd_sc_hd__o21a_1
XFILLER_204_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18315_ _18315_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
X_15527_ _15527_/A _15527_/B _15527_/C _15526_/Y vssd1 vssd1 vccd1 vccd1 _15528_/D
+ sky130_fd_sc_hd__or4b_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _12746_/D _12739_/B vssd1 vssd1 vccd1 vccd1 _17629_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_32_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19290_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19295_ _19295_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18246_ _18246_/CLK _18246_/D vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18177_ _18177_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17128_ _17129_/B _17129_/C _17127_/Y vssd1 vssd1 vccd1 vccd1 _19223_/D sky130_fd_sc_hd__a21oi_1
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09950_ _18477_/Q vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__buf_4
XFILLER_239_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03797_ _15404_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03797_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _19303_/Q _08795_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _08902_/A sky130_fd_sc_hd__mux2_1
X_17001__350 _17002__351/A vssd1 vssd1 vccd1 vccd1 _19149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09881_ _10985_/B vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__inv_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08832_ hold7/X vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107__413 _13108__414/A vssd1 vssd1 vccd1 vccd1 _17709_/CLK sky130_fd_sc_hd__inv_2
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08763_ _08761_/X _08757_/X _09635_/A vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09315_ _09315_/A vssd1 vssd1 vccd1 vccd1 _19102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _09231_/X _09244_/Y _10402_/A _18564_/Q _10403_/D vssd1 vssd1 vccd1 vccd1
+ _09247_/D sky130_fd_sc_hd__a221o_1
XFILLER_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09177_ _09177_/A vssd1 vssd1 vccd1 vccd1 _19168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11070_ _11085_/S vssd1 vssd1 vccd1 vccd1 _11079_/S sky130_fd_sc_hd__clkbuf_2
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10021_ _10021_/A vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17067__54 _17067__54/A vssd1 vssd1 vccd1 vccd1 _19203_/CLK sky130_fd_sc_hd__inv_2
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483__641 _14484__642/A vssd1 vssd1 vccd1 vccd1 _18276_/CLK sky130_fd_sc_hd__inv_2
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16692__317 _16694__319/A vssd1 vssd1 vccd1 vccd1 _19092_/CLK sky130_fd_sc_hd__inv_2
X_11972_ _19236_/Q vssd1 vssd1 vccd1 vccd1 _17179_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848__149 _15848__149/A vssd1 vssd1 vccd1 vccd1 _18824_/CLK sky130_fd_sc_hd__inv_2
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13711_ _17880_/Q _13709_/B _13709_/Y _13710_/X vssd1 vssd1 vccd1 vccd1 _17880_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10923_ _18310_/Q _10901_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10924_/A sky130_fd_sc_hd__mux2_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _14689_/X _14690_/X _14726_/S vssd1 vssd1 vccd1 vccd1 _14691_/X sky130_fd_sc_hd__mux2_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16430_ _16427_/X _16429_/Y _16437_/C vssd1 vssd1 vccd1 vccd1 _16431_/B sky130_fd_sc_hd__mux2_1
X_13642_ _14940_/A _16520_/A _13642_/S vssd1 vssd1 vccd1 vccd1 _13643_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _10854_/A vssd1 vssd1 vccd1 vccd1 _18346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _08857_/X _14244_/A _17303_/A vssd1 vssd1 vccd1 vccd1 _16362_/A sky130_fd_sc_hd__a21o_1
XFILLER_197_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ _13584_/B vssd1 vssd1 vccd1 vccd1 _13574_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10785_ _18372_/Q _10710_/X _10787_/S vssd1 vssd1 vccd1 vccd1 _10786_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18100_ _18100_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _09614_/A _15311_/Y _15285_/X vssd1 vssd1 vccd1 vccd1 _15312_/Y sky130_fd_sc_hd__a21oi_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _13095_/B _12517_/A vssd1 vssd1 vccd1 vccd1 _12524_/X sky130_fd_sc_hd__or2b_1
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19080_ _19080_/CLK _19080_/D vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16190_/X _16283_/X _16291_/Y _16214_/X vssd1 vssd1 vccd1 vccd1 _16292_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18031_ _18031_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
X_15405__905 _15407__907/A vssd1 vssd1 vccd1 vccd1 _18592_/CLK sky130_fd_sc_hd__inv_2
X_15243_ _18569_/Q _15207_/X _15239_/X _15242_/X vssd1 vssd1 vccd1 vccd1 _18569_/D
+ sky130_fd_sc_hd__o211a_1
X_12455_ _17628_/Q vssd1 vssd1 vccd1 vccd1 _12737_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ _11326_/X _18113_/Q _11412_/S vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03620_ clkbuf_0__03620_/X vssd1 vssd1 vccd1 vccd1 _15204__889/A sky130_fd_sc_hd__clkbuf_16
XFILLER_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15174_ _18453_/Q _15174_/B _16097_/A _17843_/Q vssd1 vssd1 vccd1 vccd1 _15175_/A
+ sky130_fd_sc_hd__and4b_1
X_12386_ _12638_/A _12383_/X _12647_/B _12647_/A _12366_/X _12368_/X vssd1 vssd1 vccd1
+ vccd1 _12386_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14125_ _18025_/Q _14114_/X _14124_/Y vssd1 vssd1 vccd1 vccd1 _18025_/D sky130_fd_sc_hd__o21a_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11337_ _11337_/A vssd1 vssd1 vccd1 vccd1 _18142_/D sky130_fd_sc_hd__clkbuf_1
X_15790__112 _15792__114/A vssd1 vssd1 vccd1 vccd1 _18784_/CLK sky130_fd_sc_hd__inv_2
XFILLER_126_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _13777_/X _14055_/X _14046_/X vssd1 vssd1 vccd1 vccd1 _14056_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18933_ _18933_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11268_ _18168_/Q _11267_/X _11274_/S vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13007_ _17676_/Q _12924_/X _12834_/X _17671_/Q _13006_/X vssd1 vssd1 vccd1 vccd1
+ _13010_/C sky130_fd_sc_hd__o221a_1
X_10219_ _10219_/A _10219_/B _10219_/C vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__nand3_4
X_11199_ _11199_/A vssd1 vssd1 vccd1 vccd1 _18197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18864_ _18876_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17815_ _19339_/CLK _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/Q sky130_fd_sc_hd__dfxtp_1
X_18795_ _18795_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17746_ _19336_/CLK _17746_/D vssd1 vssd1 vccd1 vccd1 _17746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14958_ _16097_/B _15076_/B vssd1 vssd1 vccd1 vccd1 _15026_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__05083_ clkbuf_0__05083_/X vssd1 vssd1 vccd1 vccd1 _17501__8/A sky130_fd_sc_hd__clkbuf_16
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13909_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13909_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17677_ _17963_/CLK _17677_/D vssd1 vssd1 vccd1 vccd1 _17677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14889_ _15086_/A vssd1 vssd1 vccd1 vccd1 _14889_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_210 _11830_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_221 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19347_ _19347_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
X_16559_ _18967_/Q _16559_/B _16559_/C _17792_/Q vssd1 vssd1 vccd1 vccd1 _16560_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ _10701_/A vssd1 vssd1 vccd1 vccd1 _09100_/X sky130_fd_sc_hd__buf_2
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19278_ _19290_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09031_ _11326_/A vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18229_ _18229_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09933_ _09933_/A vssd1 vssd1 vccd1 vccd1 _18783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _09845_/X _09860_/X _09863_/Y vssd1 vssd1 vccd1 vccd1 _18811_/D sky130_fd_sc_hd__o21a_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08815_/A vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__clkbuf_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _09795_/A vssd1 vssd1 vccd1 vccd1 _18834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _18066_/Q _08746_/B vssd1 vssd1 vccd1 vccd1 _13873_/B sky130_fd_sc_hd__nand2_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15391__894 _15391__894/A vssd1 vssd1 vccd1 vccd1 _18581_/CLK sky130_fd_sc_hd__inv_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10570_ _10120_/X _18497_/Q _10574_/S vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__mux2_1
X_16316__215 _16318__217/A vssd1 vssd1 vccd1 vccd1 _18931_/CLK sky130_fd_sc_hd__inv_2
XFILLER_194_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _09972_/A vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17008__356 _17008__356/A vssd1 vssd1 vccd1 vccd1 _19155_/CLK sky130_fd_sc_hd__inv_2
XFILLER_154_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _17769_/Q _17423_/B vssd1 vssd1 vccd1 vccd1 _12293_/S sky130_fd_sc_hd__nand2_2
XFILLER_181_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12171_ _12166_/X _12171_/B vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__and2b_1
XFILLER_135_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15658__962 _15660__964/A vssd1 vssd1 vccd1 vccd1 _18679_/CLK sky130_fd_sc_hd__inv_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ _18227_/Q _11065_/X _11122_/S vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15930_ _15932_/B _15930_/B vssd1 vssd1 vccd1 vccd1 _15931_/B sky130_fd_sc_hd__nand2_1
X_11053_ _18665_/Q vssd1 vssd1 vccd1 vccd1 _11053_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _18762_/Q _09955_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16700__324 _16700__324/A vssd1 vssd1 vccd1 vccd1 _19099_/CLK sky130_fd_sc_hd__inv_2
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _15861_/A vssd1 vssd1 vccd1 vccd1 _15861_/X sky130_fd_sc_hd__buf_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14329__518 _14329__518/A vssd1 vssd1 vccd1 vccd1 _18153_/CLK sky130_fd_sc_hd__inv_2
X_17600_ _17609_/CLK _17600_/D vssd1 vssd1 vccd1 vccd1 _17600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18580_ _18580_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _18031_/CLK _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _19249_/Q vssd1 vssd1 vccd1 vccd1 _17225_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17462_ _17741_/Q _19335_/Q _17468_/S vssd1 vssd1 vccd1 vccd1 _17463_/B sky130_fd_sc_hd__mux2_1
X_10906_ _10906_/A vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _19152_/Q _18417_/Q _18311_/Q _18295_/Q _14563_/X _14564_/X vssd1 vssd1 vccd1
+ vccd1 _14675_/B sky130_fd_sc_hd__mux4_1
XFILLER_189_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19201_ _19201_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
X_16413_ _16413_/A _16413_/B vssd1 vssd1 vccd1 vccd1 _16416_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ _13635_/B vssd1 vssd1 vccd1 vccd1 _13626_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10837_ _18353_/Q _10794_/X _10843_/S vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ _19132_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13556_ _13441_/X _13549_/X _13553_/Y _13555_/X vssd1 vssd1 vccd1 vccd1 _17829_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10768_ _18379_/Q _10713_/X _10768_/S vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12507_ _12408_/X _12770_/A _12580_/A vssd1 vssd1 vccd1 vccd1 _12507_/Y sky130_fd_sc_hd__a21oi_1
X_19063_ _19063_/CLK _19063_/D vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16275_ _18531_/Q _18539_/Q _18547_/Q _18555_/Q _10420_/A _16117_/X vssd1 vssd1 vccd1
+ vccd1 _16276_/B sky130_fd_sc_hd__mux4_2
X_13487_ _13540_/A vssd1 vssd1 vccd1 vccd1 _14186_/D sky130_fd_sc_hd__clkbuf_4
X_10699_ _18408_/Q _10698_/X _10705_/S vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18014_ _18014_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15226_ _18828_/Q _18820_/Q _18812_/Q _18679_/Q _15214_/X _15225_/X vssd1 vssd1 vccd1
+ vccd1 _15226_/X sky130_fd_sc_hd__mux4_1
X_12438_ _12436_/X _12437_/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12438_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12369_ _12706_/A _12717_/C _12717_/B _12717_/A _12366_/X _12368_/X vssd1 vssd1 vccd1
+ vccd1 _12369_/X sky130_fd_sc_hd__mux4_2
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ _16570_/A vssd1 vssd1 vccd1 vccd1 _14108_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _14039_/A vssd1 vssd1 vccd1 vccd1 _14039_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18916_ _18919_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ _18847_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03396_ clkbuf_0__03396_/X vssd1 vssd1 vccd1 vccd1 _14759_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09580_ _10219_/A _09639_/A _10219_/C vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__nand3_2
X_18778_ _18778_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17729_ _17737_/CLK _17729_/D vssd1 vssd1 vccd1 vccd1 _17729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17061__49 _17061__49/A vssd1 vssd1 vccd1 vccd1 _19198_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15797__118 _15798__119/A vssd1 vssd1 vccd1 vccd1 _18790_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16090__203 _16090__203/A vssd1 vssd1 vccd1 vccd1 _18908_/CLK sky130_fd_sc_hd__inv_2
XFILLER_163_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ _09856_/B _09857_/C _09857_/A vssd1 vssd1 vccd1 vccd1 _09016_/C sky130_fd_sc_hd__a21o_1
X_14434__602 _14434__602/A vssd1 vssd1 vccd1 vccd1 _18237_/CLK sky130_fd_sc_hd__inv_2
XFILLER_151_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09916_ _10094_/A _10274_/A vssd1 vssd1 vccd1 vccd1 _09932_/S sky130_fd_sc_hd__nor2_2
XFILLER_113_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09847_ _16902_/A vssd1 vssd1 vccd1 vccd1 _16875_/S sky130_fd_sc_hd__buf_2
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09778_/A vssd1 vssd1 vccd1 vccd1 _18841_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08729_ _13128_/A _11779_/A vssd1 vssd1 vccd1 vccd1 _08855_/C sky130_fd_sc_hd__nor2_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11740_ _17915_/Q _18558_/Q _17826_/Q vssd1 vssd1 vccd1 vccd1 _11741_/A sky130_fd_sc_hd__mux2_4
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _17507_/Q _09697_/A _11671_/S vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _17787_/Q _13393_/X _13409_/Y vssd1 vssd1 vccd1 vccd1 _17787_/D sky130_fd_sc_hd__o21a_1
X_10622_ _18444_/Q _10112_/A _10630_/S vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13341_ _17773_/Q vssd1 vssd1 vccd1 vccd1 _17101_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ _10553_/A vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _16060_/A _16061_/B vssd1 vssd1 vccd1 vccd1 _18886_/D sky130_fd_sc_hd__nor2_1
X_13272_ _13271_/X _13259_/X _13260_/X vssd1 vssd1 vccd1 vccd1 _13272_/Y sky130_fd_sc_hd__a21oi_1
X_10484_ _18535_/Q _10342_/X _10484_/S vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15011_ _18461_/Q _14991_/X _15010_/X _14993_/X vssd1 vssd1 vccd1 vccd1 _15012_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12223_ _12229_/A vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__buf_1
XFILLER_154_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12154_ _12149_/X _12154_/B vssd1 vssd1 vccd1 vccd1 _12155_/A sky130_fd_sc_hd__and2b_1
XFILLER_123_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11105_ _11105_/A vssd1 vssd1 vccd1 vccd1 _18235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12085_ _17264_/A _19260_/Q _19261_/Q _17276_/A _11980_/X _11977_/S vssd1 vssd1 vccd1
+ vccd1 _12085_/X sky130_fd_sc_hd__mux4_1
X_16962_ _18249_/Q _18241_/Q _18233_/Q _18225_/Q _16799_/X _16801_/X vssd1 vssd1 vccd1
+ vccd1 _16963_/B sky130_fd_sc_hd__mux4_1
X_18701_ _18701_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15913_ _18870_/Q _15913_/B vssd1 vssd1 vccd1 vccd1 _15936_/C sky130_fd_sc_hd__xnor2_1
X_11036_ _18261_/Q _09139_/X _11040_/S vssd1 vssd1 vccd1 vccd1 _11037_/A sky130_fd_sc_hd__mux2_1
X_16893_ _16893_/A vssd1 vssd1 vccd1 vccd1 _16893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18632_ _18632_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03181_ clkbuf_0__03181_/X vssd1 vssd1 vccd1 vccd1 _14447__613/A sky130_fd_sc_hd__clkbuf_16
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18563_ _18563_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_1
X_12987_ _12975_/X _12987_/B vssd1 vssd1 vccd1 vccd1 _12988_/A sky130_fd_sc_hd__and2b_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14724_/X _14725_/X _14726_/S vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__mux2_1
X_17514_ _17514_/CLK _17514_/D vssd1 vssd1 vccd1 vccd1 _17514_/Q sky130_fd_sc_hd__dfxtp_1
X_11938_ _11938_/A vssd1 vssd1 vccd1 vccd1 _12017_/S sky130_fd_sc_hd__buf_2
X_18494_ _18494_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17445_ _17746_/Q _19330_/Q _17451_/S vssd1 vssd1 vccd1 vccd1 _17446_/B sky130_fd_sc_hd__mux2_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _19175_/Q _19167_/Q _19199_/Q _18334_/Q _14580_/A _14546_/X vssd1 vssd1 vccd1
+ vccd1 _14657_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11869_ _17930_/Q _11869_/B vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__or2_4
XFILLER_232_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13608_ _17847_/Q _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17376_ _19277_/Q _17490_/B vssd1 vssd1 vccd1 vccd1 _17377_/D sky130_fd_sc_hd__xnor2_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14588_ _16536_/C vssd1 vssd1 vccd1 vccd1 _14623_/A sky130_fd_sc_hd__clkbuf_2
X_12342__402 _12342__402/A vssd1 vssd1 vccd1 vccd1 _17583_/CLK sky130_fd_sc_hd__inv_2
XFILLER_220_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19115_ _19115_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_1
X_16327_ _16333_/A vssd1 vssd1 vccd1 vccd1 _16327_/X sky130_fd_sc_hd__buf_1
XFILLER_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ _16520_/A _13523_/X _13526_/X _15927_/A _15083_/B vssd1 vssd1 vccd1 vccd1
+ _17825_/D sky130_fd_sc_hd__a221o_1
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19046_ _19046_/CLK _19046_/D vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _18599_/Q _18615_/Q _18741_/Q _18522_/Q _16195_/X _16112_/X vssd1 vssd1 vccd1
+ vccd1 _16259_/B sky130_fd_sc_hd__mux4_1
X_15209_ _15273_/A vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16189_ _18916_/Q _16098_/X _16188_/Y _14247_/X vssd1 vssd1 vccd1 vccd1 _18916_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_9 _09726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15418__915 _15419__916/A vssd1 vssd1 vccd1 vccd1 _18602_/CLK sky130_fd_sc_hd__inv_2
X_09701_ _09716_/S vssd1 vssd1 vccd1 vccd1 _09710_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _18922_/Q _16294_/C _09631_/X vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09563_ _09578_/S vssd1 vssd1 vccd1 vccd1 _09572_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17034__27 _17036__29/A vssd1 vssd1 vccd1 vccd1 _19176_/CLK sky130_fd_sc_hd__inv_2
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ _09494_/A vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12910_ _12910_/A vssd1 vssd1 vccd1 vccd1 _17666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _13783_/X _13885_/X _13880_/X vssd1 vssd1 vccd1 vccd1 _13890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12841_ _17645_/Q _13093_/B vssd1 vssd1 vccd1 vccd1 _12841_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15558_/X _15559_/Y _15553_/X vssd1 vssd1 vccd1 vccd1 _18646_/D sky130_fd_sc_hd__a21oi_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12772_ _12524_/X _13081_/B _12772_/C _12850_/A vssd1 vssd1 vccd1 vccd1 _12773_/D
+ sky130_fd_sc_hd__and4bb_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04586_ clkbuf_0__04586_/X vssd1 vssd1 vccd1 vccd1 _16706__329/A sky130_fd_sc_hd__clkbuf_16
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A vssd1 vssd1 vccd1 vccd1 _14511_/X sky130_fd_sc_hd__buf_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11717_/X _17911_/Q vssd1 vssd1 vccd1 vccd1 _11724_/A sky130_fd_sc_hd__and2b_4
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15491_ _17832_/Q _15494_/B vssd1 vssd1 vccd1 vccd1 _15492_/B sky130_fd_sc_hd__xor2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _19251_/Q vssd1 vssd1 vccd1 vccd1 _17237_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11654_ _11654_/A vssd1 vssd1 vccd1 vccd1 _17532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ _17161_/A vssd1 vssd1 vccd1 vccd1 _19231_/D sky130_fd_sc_hd__clkbuf_1
X_10605_ _10605_/A vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11585_ _17580_/Q _10690_/A _11593_/S vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03399_ clkbuf_0__03399_/X vssd1 vssd1 vccd1 vccd1 _14764__704/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16112_ _16198_/A vssd1 vssd1 vccd1 vccd1 _16112_/X sky130_fd_sc_hd__buf_2
X_13324_ _17768_/Q _13304_/X _13323_/Y vssd1 vssd1 vccd1 vccd1 _17768_/D sky130_fd_sc_hd__o21a_1
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665__300 _16666__301/A vssd1 vssd1 vccd1 vccd1 _19074_/CLK sky130_fd_sc_hd__inv_2
X_17092_ _17776_/Q _17774_/Q _12214_/A vssd1 vssd1 vccd1 vccd1 _17092_/X sky130_fd_sc_hd__a21bo_1
XFILLER_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10536_ _18512_/Q _10339_/X _10538_/S vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16043_ _16044_/B _16050_/A _16042_/Y _16010_/X vssd1 vssd1 vccd1 vccd1 _18877_/D
+ sky130_fd_sc_hd__a211oi_1
X_13255_ _17745_/Q _13252_/X _13254_/Y vssd1 vssd1 vccd1 vccd1 _17745_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10467_ _10467_/A vssd1 vssd1 vccd1 vccd1 _18543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _12206_/A vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17969_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13186_ _17731_/Q _13208_/B vssd1 vssd1 vccd1 vccd1 _13186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _16172_/A vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12137_ _12132_/X _12137_/B vssd1 vssd1 vccd1 vccd1 _12138_/A sky130_fd_sc_hd__and2b_1
X_17994_ _18021_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03402_ _14777_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03402_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__07170_ _11876_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07170_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12068_ _12035_/X _12036_/X _12066_/X _12067_/X _12109_/S _12116_/A vssd1 vssd1 vccd1
+ vccd1 _12069_/B sky130_fd_sc_hd__mux4_1
X_16945_ _18208_/Q _18128_/Q _19185_/Q _18256_/Q _16822_/X _16823_/X vssd1 vssd1 vccd1
+ vccd1 _16946_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11019_ _11019_/A vssd1 vssd1 vccd1 vccd1 _18269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16876_ _16900_/A vssd1 vssd1 vccd1 vccd1 _16963_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_226_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18615_ _18615_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13101__408 _13102__409/A vssd1 vssd1 vccd1 vccd1 _17704_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03164_ clkbuf_0__03164_/X vssd1 vssd1 vccd1 vccd1 _14358__541/A sky130_fd_sc_hd__clkbuf_16
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18546_ _18546_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03195_ _14512_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03195_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_244_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03095_ clkbuf_0__03095_/X vssd1 vssd1 vccd1 vccd1 _14162__441/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14709_ _18859_/Q _18353_/Q _19194_/Q _18361_/Q _14553_/X _14600_/X vssd1 vssd1 vccd1
+ vccd1 _14709_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18477_ _18477_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17428_ _17751_/Q _19325_/Q _17497_/B vssd1 vssd1 vccd1 vccd1 _17429_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _17359_/A vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19029_ _19040_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08994_ _09880_/B vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _09615_/A _09628_/A vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__and2_1
XFILLER_244_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09546_ _08910_/X _18958_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09477_ _09467_/B _09477_/B _09477_/C vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__and3b_1
XFILLER_169_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04371_ clkbuf_0__04371_/X vssd1 vssd1 vccd1 vccd1 _16332__229/A sky130_fd_sc_hd__clkbuf_16
XFILLER_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _11370_/A vssd1 vssd1 vccd1 vccd1 _18129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03184_ clkbuf_0__03184_/X vssd1 vssd1 vccd1 vccd1 _14461__624/A sky130_fd_sc_hd__clkbuf_16
XFILLER_192_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _10321_/A vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _17947_/Q _17691_/Q _13053_/S vssd1 vssd1 vccd1 vccd1 _13041_/B sky130_fd_sc_hd__mux2_1
X_14371__552 _14373__554/A vssd1 vssd1 vccd1 vccd1 _18187_/CLK sky130_fd_sc_hd__inv_2
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ _18634_/Q _10195_/X _10254_/S vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10183_ _18478_/Q vssd1 vssd1 vccd1 vccd1 _10183_/X sky130_fd_sc_hd__buf_4
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14991_ _14991_/A vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16660__296 _16663__299/A vssd1 vssd1 vccd1 vccd1 _19070_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _13161_/X _13929_/B _13941_/Y _13937_/X vssd1 vssd1 vccd1 vccd1 _17958_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _13873_/A _13873_/B _13873_/C _13873_/D vssd1 vssd1 vccd1 vccd1 _16516_/D
+ sky130_fd_sc_hd__nor4_4
XFILLER_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15612_ _18656_/Q _15612_/B vssd1 vssd1 vccd1 vccd1 _15612_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18400_ _18400_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
X_12824_ _12824_/A vssd1 vssd1 vccd1 vccd1 _17649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16592_ _19025_/Q _16593_/C _16591_/Y vssd1 vssd1 vccd1 vccd1 _19025_/D sky130_fd_sc_hd__o21a_1
XFILLER_216_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _18644_/Q _18643_/Q _15543_/C vssd1 vssd1 vccd1 vccd1 _15557_/C sky130_fd_sc_hd__and3_1
XFILLER_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18331_ _18331_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
X_12755_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__and3_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04569_ clkbuf_0__04569_/X vssd1 vssd1 vccd1 vccd1 _16638__279/A sky130_fd_sc_hd__clkbuf_16
XFILLER_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ _13845_/A _11707_/S vssd1 vssd1 vccd1 vccd1 _11706_/Y sky130_fd_sc_hd__nor2_8
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18262_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
X_15474_ _17838_/Q _17837_/Q _17836_/Q _15517_/B vssd1 vssd1 vccd1 vccd1 _15505_/B
+ sky130_fd_sc_hd__or4_2
X_12686_ _17614_/Q _12686_/B vssd1 vssd1 vccd1 vccd1 _12694_/D sky130_fd_sc_hd__and2_1
XFILLER_124_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17213_ _17213_/A vssd1 vssd1 vccd1 vccd1 _19245_/D sky130_fd_sc_hd__clkbuf_1
X_14425_ _14425_/A vssd1 vssd1 vccd1 vccd1 _14425_/X sky130_fd_sc_hd__buf_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11637_ _11637_/A hold2/X vssd1 vssd1 vccd1 vccd1 _11653_/S sky130_fd_sc_hd__or2_2
X_18193_ _18193_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17144_ _17142_/X _17289_/A _17144_/C vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__and3b_1
XFILLER_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14356_ _14380_/A vssd1 vssd1 vccd1 vccd1 _14356_/X sky130_fd_sc_hd__buf_1
XFILLER_156_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ _11568_/A vssd1 vssd1 vccd1 vccd1 _17588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12226__372 _12226__372/A vssd1 vssd1 vccd1 vccd1 _17536_/CLK sky130_fd_sc_hd__inv_2
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13307_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__buf_2
XFILLER_7_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17075_ _17081_/A vssd1 vssd1 vccd1 vccd1 _17075_/X sky130_fd_sc_hd__buf_1
X_10519_ _10519_/A vssd1 vssd1 vccd1 vccd1 _18520_/D sky130_fd_sc_hd__clkbuf_1
X_14287_ _14287_/A vssd1 vssd1 vccd1 vccd1 _14287_/X sky130_fd_sc_hd__buf_1
X_11499_ _18045_/Q _11329_/A _11503_/S vssd1 vssd1 vccd1 vccd1 _11500_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16026_ _16024_/X _16025_/Y _16010_/X vssd1 vssd1 vccd1 vccd1 _18873_/D sky130_fd_sc_hd__a21oi_1
X_13238_ _13237_/X _13232_/X _13224_/X vssd1 vssd1 vccd1 vccd1 _13238_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14272__472 _14274__474/A vssd1 vssd1 vccd1 vccd1 _18107_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13169_ _14113_/A _13169_/B vssd1 vssd1 vccd1 vccd1 _13212_/B sky130_fd_sc_hd__and2_1
XFILLER_111_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17977_ _18001_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16928_ _18183_/Q _18175_/Q _18167_/Q _18159_/Q _16881_/X _16882_/X vssd1 vssd1 vccd1
+ vccd1 _16929_/B sky130_fd_sc_hd__mux4_1
XFILLER_226_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16859_ _16819_/X _16852_/Y _16854_/Y _16856_/Y _16858_/Y vssd1 vssd1 vccd1 vccd1
+ _16859_/X sky130_fd_sc_hd__o32a_1
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09400_ _08917_/X _19065_/Q _09406_/S vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03147_ clkbuf_0__03147_/X vssd1 vssd1 vccd1 vccd1 _14274__474/A sky130_fd_sc_hd__clkbuf_16
XFILLER_241_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _09331_/A vssd1 vssd1 vccd1 vccd1 _19095_/D sky130_fd_sc_hd__clkbuf_1
X_18529_ _18529_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03178_ _14425_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03178_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_240_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _18479_/Q vssd1 vssd1 vccd1 vccd1 _09262_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_179_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09193_ _09193_/A vssd1 vssd1 vccd1 vccd1 _19161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17079__63 _17080__64/A vssd1 vssd1 vccd1 vccd1 _19212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08977_ _08977_/A vssd1 vssd1 vccd1 vccd1 _19218_/D sky130_fd_sc_hd__clkbuf_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15652__957 _15654__959/A vssd1 vssd1 vccd1 vccd1 _18674_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18870_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _10885_/S vssd1 vssd1 vccd1 vccd1 _10879_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09529_/A vssd1 vssd1 vccd1 vccd1 _18966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _12408_/A _12392_/A _12580_/A vssd1 vssd1 vccd1 vccd1 _12540_/Y sky130_fd_sc_hd__a21oi_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14854__776 _14857__779/A vssd1 vssd1 vccd1 vccd1 _18421_/CLK sky130_fd_sc_hd__inv_2
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _17624_/Q vssd1 vssd1 vccd1 vccd1 _12727_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ _13488_/A input34/X _14218_/S vssd1 vssd1 vccd1 vccd1 _14211_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11422_ _18106_/Q _11259_/X _11430_/S vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__mux2_1
X_15190_ _15535_/A _15190_/B vssd1 vssd1 vccd1 vccd1 _15630_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11353_ _18136_/Q _11267_/X _11357_/S vssd1 vssd1 vccd1 vccd1 _11354_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03167_ clkbuf_0__03167_/X vssd1 vssd1 vccd1 vccd1 _14378__558/A sky130_fd_sc_hd__clkbuf_16
XFILLER_180_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10304_ _18611_/Q _10192_/X _10308_/S vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__mux2_1
X_14072_ _14072_/A _14083_/B vssd1 vssd1 vccd1 vccd1 _14072_/Y sky130_fd_sc_hd__nor2_2
X_11284_ _11284_/A vssd1 vssd1 vccd1 vccd1 _18163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03098_ clkbuf_0__03098_/X vssd1 vssd1 vccd1 vccd1 _14252__456/A sky130_fd_sc_hd__clkbuf_16
X_13023_ _13023_/A vssd1 vssd1 vccd1 vccd1 _17686_/D sky130_fd_sc_hd__clkbuf_1
X_17900_ _17923_/CLK _17900_/D vssd1 vssd1 vccd1 vccd1 _17900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10235_ _10235_/A vssd1 vssd1 vccd1 vccd1 _18672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18880_ _18886_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17831_ _17935_/CLK _17831_/D vssd1 vssd1 vccd1 vccd1 _17831_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10166_ _10166_/A vssd1 vssd1 vccd1 vccd1 _18699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17762_ _19288_/CLK _17762_/D vssd1 vssd1 vccd1 vccd1 _17762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14974_ _14991_/A vssd1 vssd1 vccd1 vccd1 _15080_/C sky130_fd_sc_hd__inv_2
X_10097_ _10097_/A vssd1 vssd1 vccd1 vccd1 _18726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ _16713_/A vssd1 vssd1 vccd1 vccd1 _19109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _13943_/B vssd1 vssd1 vccd1 vccd1 _13925_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17693_ _18007_/CLK _17693_/D vssd1 vssd1 vccd1 vccd1 _17693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13856_ input70/X _13867_/B vssd1 vssd1 vccd1 vccd1 _13856_/X sky130_fd_sc_hd__and2_1
XFILLER_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _12807_/A vssd1 vssd1 vccd1 vccd1 _17644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16575_ _19019_/Q _16576_/C _16574_/Y vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__o21a_1
X_13787_ _13786_/X _13778_/X _13774_/X vssd1 vssd1 vccd1 vccd1 _13787_/Y sky130_fd_sc_hd__a21oi_1
X_10999_ _10999_/A vssd1 vssd1 vccd1 vccd1 _18278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18314_ _18314_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_1
X_12738_ _12737_/A _12736_/A _12734_/X vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__o21ai_1
X_15526_ _15498_/Y _15499_/X _15525_/X vssd1 vssd1 vccd1 vccd1 _15526_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _19294_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18245_ _18245_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
X_12669_ _12673_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _17608_/D sky130_fd_sc_hd__nor2_1
XFILLER_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14378__558 _14378__558/A vssd1 vssd1 vccd1 vccd1 _18193_/CLK sky130_fd_sc_hd__inv_2
XFILLER_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14755__696 _14757__698/A vssd1 vssd1 vccd1 vccd1 _18339_/CLK sky130_fd_sc_hd__inv_2
XFILLER_175_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_72_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19037_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18176_ _18176_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17127_ _17129_/B _17129_/C _17126_/X vssd1 vssd1 vccd1 vccd1 _17127_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03796_ _15398_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03796_/X sky130_fd_sc_hd__clkbuf_16
X_08900_ _08900_/A vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16009_ _18870_/Q _16020_/B vssd1 vssd1 vccd1 vccd1 _16009_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _10583_/B _09880_/B _09894_/B vssd1 vssd1 vccd1 vccd1 _10985_/B sky130_fd_sc_hd__and3_2
XFILLER_112_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ hold12/X vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16678__310 _16680__312/A vssd1 vssd1 vccd1 vccd1 _19084_/CLK sky130_fd_sc_hd__inv_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08762_ hold4/A hold14/A _18925_/Q vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__and3_1
XFILLER_245_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14322__513 _14323__514/A vssd1 vssd1 vccd1 vccd1 _18148_/CLK sky130_fd_sc_hd__inv_2
X_09314_ _08933_/X _19102_/Q _09318_/S vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _18564_/Q _18559_/Q vssd1 vssd1 vccd1 vccd1 _10403_/D sky130_fd_sc_hd__xnor2_2
XFILLER_107_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13114__418 _13115__419/A vssd1 vssd1 vccd1 vccd1 _17714_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14279__478 _14280__479/A vssd1 vssd1 vccd1 vccd1 _18113_/CLK sky130_fd_sc_hd__inv_2
X_09176_ _19168_/Q _09100_/X _09178_/S vssd1 vssd1 vccd1 vccd1 _09177_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10020_ _18755_/Q _09951_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15887__177 _15889__179/A vssd1 vssd1 vccd1 vccd1 _18853_/CLK sky130_fd_sc_hd__inv_2
XFILLER_245_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11971_ _17777_/Q vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13710_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ _10922_/A vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _18858_/Q _18352_/Q _19193_/Q _18360_/Q _14553_/X _14600_/X vssd1 vssd1 vccd1
+ vccd1 _14690_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ _17859_/Q vssd1 vssd1 vccd1 vccd1 _14940_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10853_ _18346_/Q _10789_/X _10861_/S vssd1 vssd1 vccd1 vccd1 _10854_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13572_ _13589_/S vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__buf_2
X_10784_ _10784_/A vssd1 vssd1 vccd1 vccd1 _18373_/D sky130_fd_sc_hd__clkbuf_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15311_ _15311_/A vssd1 vssd1 vccd1 vccd1 _15311_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12523_/A vssd1 vssd1 vccd1 vccd1 _13095_/B sky130_fd_sc_hd__buf_4
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16291_ _16291_/A _16291_/B vssd1 vssd1 vccd1 vccd1 _16291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18030_ _18031_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
X_15242_ _16064_/A vssd1 vssd1 vccd1 vccd1 _15242_/X sky130_fd_sc_hd__clkbuf_2
X_12454_ _17626_/Q vssd1 vssd1 vccd1 vccd1 _12727_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11405_ _11405_/A vssd1 vssd1 vccd1 vccd1 _18114_/D sky130_fd_sc_hd__clkbuf_1
X_12385_ _17603_/Q vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14124_ _13748_/A _14120_/X _14123_/X vssd1 vssd1 vccd1 vccd1 _14124_/Y sky130_fd_sc_hd__a21oi_1
X_11336_ _11335_/X _18142_/Q _11336_/S vssd1 vssd1 vccd1 vccd1 _11337_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14055_ _14055_/A vssd1 vssd1 vccd1 vccd1 _14055_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18932_ _18932_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_2
X_11267_ _18666_/Q vssd1 vssd1 vccd1 vccd1 _11267_/X sky130_fd_sc_hd__clkbuf_4
X_13006_ _17682_/Q _12845_/A _12838_/A _17685_/Q _13005_/Y vssd1 vssd1 vccd1 vccd1
+ _13006_/X sky130_fd_sc_hd__o221a_1
X_10218_ _10218_/A vssd1 vssd1 vccd1 vccd1 _18679_/D sky130_fd_sc_hd__clkbuf_1
X_18863_ _18876_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11198_ _18197_/Q _11059_/X _11202_/S vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17814_ _19108_/CLK _17814_/D vssd1 vssd1 vccd1 vccd1 _17814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_239_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10149_ _18706_/Q _10063_/X _10149_/S vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18794_ _18794_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ _19336_/CLK _17745_/D vssd1 vssd1 vccd1 vccd1 _17745_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__05082_ clkbuf_0__05082_/X vssd1 vssd1 vccd1 vccd1 _17420__109/A sky130_fd_sc_hd__clkbuf_16
XFILLER_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14957_ _14960_/B _14963_/B _14957_/C vssd1 vssd1 vccd1 vccd1 _15076_/B sky130_fd_sc_hd__nor3_1
XFILLER_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13908_/A vssd1 vssd1 vccd1 vccd1 _13908_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17676_ _19037_/CLK _17676_/D vssd1 vssd1 vccd1 vccd1 _17676_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_200 _17454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_211 _11833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_222 _10175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16627_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16627_/X sky130_fd_sc_hd__buf_1
X_13839_ _17923_/Q _13829_/X _13838_/X _13826_/X vssd1 vssd1 vccd1 vccd1 _17923_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19346_ _19346_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15509_ _18647_/Q _15509_/B vssd1 vssd1 vccd1 vccd1 _15524_/A sky130_fd_sc_hd__xnor2_1
X_19277_ _19290_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16489_ _18980_/Q _16499_/B vssd1 vssd1 vccd1 vccd1 _16489_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ _18667_/Q vssd1 vssd1 vccd1 vccd1 _11326_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_248_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18228_ _18228_/CLK _18228_/D vssd1 vssd1 vccd1 vccd1 _18228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18159_ _18159_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09932_ _18783_/Q _09280_/X _09932_/S vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _09845_/X _09860_/X _09895_/C vssd1 vssd1 vccd1 vccd1 _09863_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _19323_/Q _08724_/X _08822_/S vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__mux2_1
X_14805__737 _14807__739/A vssd1 vssd1 vccd1 vccd1 _18380_/CLK sky130_fd_sc_hd__inv_2
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _18834_/Q _09749_/X _09800_/S vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__mux2_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08745_ _11787_/B vssd1 vssd1 vccd1 vccd1 _08747_/B sky130_fd_sc_hd__inv_2
XFILLER_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09228_ _18560_/Q vssd1 vssd1 vccd1 vccd1 _09972_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09159_ _09159_/A vssd1 vssd1 vccd1 vccd1 _19176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12170_ _17528_/Q _17723_/Q _12170_/S vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15854__154 _15854__154/A vssd1 vssd1 vccd1 vccd1 _18829_/CLK sky130_fd_sc_hd__inv_2
X_11121_ _11121_/A vssd1 vssd1 vccd1 vccd1 _18228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11052_ _11052_/A vssd1 vssd1 vccd1 vccd1 _18256_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10003_ _10003_/A vssd1 vssd1 vccd1 vccd1 _18763_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_55_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _18031_/CLK _17530_/D vssd1 vssd1 vccd1 vccd1 _17530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ _19247_/Q _19248_/Q _11956_/S vssd1 vssd1 vccd1 vccd1 _11954_/X sky130_fd_sc_hd__mux2_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _18330_/Q _14543_/A _14623_/A _14741_/X vssd1 vssd1 vccd1 vccd1 _18330_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15411__910 _15413__912/A vssd1 vssd1 vccd1 vccd1 _18597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_229_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _18317_/Q _10904_/X _10911_/S vssd1 vssd1 vccd1 vccd1 _10906_/A sky130_fd_sc_hd__mux2_1
X_17461_ _17461_/A vssd1 vssd1 vccd1 vccd1 _19334_/D sky130_fd_sc_hd__clkbuf_1
X_14673_ _14669_/X _14672_/X _14673_/S vssd1 vssd1 vccd1 vccd1 _14673_/X sky130_fd_sc_hd__mux2_2
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19200_ _19200_/CLK _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
X_13624_ _13642_/S vssd1 vssd1 vccd1 vccd1 _13635_/B sky130_fd_sc_hd__clkbuf_2
X_16412_ _17804_/Q _16412_/B vssd1 vssd1 vccd1 vccd1 _16413_/B sky130_fd_sc_hd__and2_1
XFILLER_232_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10836_ _10836_/A vssd1 vssd1 vccd1 vccd1 _18354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15665__967 _15667__969/A vssd1 vssd1 vccd1 vccd1 _18684_/CLK sky130_fd_sc_hd__inv_2
XFILLER_232_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19131_ _19132_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13555_ _13636_/A vssd1 vssd1 vccd1 vccd1 _13555_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10767_ _10767_/A vssd1 vssd1 vccd1 vccd1 _18380_/D sky130_fd_sc_hd__clkbuf_1
X_12506_ _18008_/Q vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16274_ _18920_/Q _16164_/X _16273_/Y _16216_/X vssd1 vssd1 vccd1 vccd1 _18920_/D
+ sky130_fd_sc_hd__o211a_1
X_19062_ _19062_/CLK _19062_/D vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _13486_/A vssd1 vssd1 vccd1 vccd1 _17808_/D sky130_fd_sc_hd__clkbuf_1
X_10698_ _10698_/A vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18013_ _18013_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15225_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__buf_2
X_12437_ _12647_/A _17604_/Q _12440_/S vssd1 vssd1 vccd1 vccd1 _12437_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03602_ clkbuf_0__03602_/X vssd1 vssd1 vccd1 vccd1 _15172__878/A sky130_fd_sc_hd__clkbuf_16
X_15156_ _15168_/A vssd1 vssd1 vccd1 vccd1 _15156_/X sky130_fd_sc_hd__buf_1
X_12368_ _12487_/S vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__buf_2
XFILLER_236_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _18019_/Q _14092_/X _14106_/Y vssd1 vssd1 vccd1 vccd1 _18019_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11319_ _11165_/X _18147_/Q _11319_/S vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12299_ _17557_/Q _17487_/B vssd1 vssd1 vccd1 vccd1 _12299_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14038_ _17993_/Q _14032_/X _14037_/Y vssd1 vssd1 vccd1 vccd1 _17993_/D sky130_fd_sc_hd__o21a_1
X_18915_ _18919_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18846_ _18846_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03395_ clkbuf_0__03395_/X vssd1 vssd1 vccd1 vccd1 _14870_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_110_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18777_ _18777_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17046__36 _17048__38/A vssd1 vssd1 vccd1 vccd1 _19185_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15989_ _15989_/A vssd1 vssd1 vccd1 vccd1 _16024_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_208_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17728_ _17878_/CLK _17728_/D vssd1 vssd1 vccd1 vccd1 _17728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _17969_/CLK _17659_/D vssd1 vssd1 vccd1 vccd1 _17659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19329_ _19329_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09013_ _18807_/Q _09880_/B vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__and2b_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14811__741 _14813__743/A vssd1 vssd1 vccd1 vccd1 _18384_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__04849_ clkbuf_0__04849_/X vssd1 vssd1 vccd1 vccd1 _17071__57/A sky130_fd_sc_hd__clkbuf_16
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09915_ _10138_/C _10424_/A _09975_/C vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__nand3b_4
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09846_ _18810_/Q vssd1 vssd1 vccd1 vccd1 _16902_/A sky130_fd_sc_hd__buf_2
XFILLER_219_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _08871_/X _18841_/Q _09781_/S vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__mux2_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16322__220 _16323__221/A vssd1 vssd1 vccd1 vccd1 _18936_/CLK sky130_fd_sc_hd__inv_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ input67/X _19145_/Q _14243_/C vssd1 vssd1 vccd1 vccd1 _08728_/X sky130_fd_sc_hd__and3_4
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11670_ _11670_/A vssd1 vssd1 vccd1 vccd1 _17508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10621_ _10636_/S vssd1 vssd1 vccd1 vccd1 _10630_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_169_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ _13431_/B vssd1 vssd1 vccd1 vccd1 _16518_/B sky130_fd_sc_hd__buf_6
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _18505_/Q _10120_/A _10556_/S vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13755_/A vssd1 vssd1 vccd1 vccd1 _13271_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10483_ _10483_/A vssd1 vssd1 vccd1 vccd1 _18536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _18461_/Q _15014_/C vssd1 vssd1 vccd1 vccd1 _15010_/X sky130_fd_sc_hd__xor2_1
XFILLER_154_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14335__523 _14336__524/A vssd1 vssd1 vccd1 vccd1 _18158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144__855 _15147__858/A vssd1 vssd1 vccd1 vccd1 _18531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12153_ _17523_/Q _17728_/Q _12153_/S vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__mux2_1
XFILLER_194_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11104_ _09055_/X _18235_/Q _11104_/S vssd1 vssd1 vccd1 vccd1 _11105_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12084_ _12084_/A vssd1 vssd1 vccd1 vccd1 _12084_/Y sky130_fd_sc_hd__clkinv_2
X_16961_ _16957_/X _16960_/X _16980_/S vssd1 vssd1 vccd1 vccd1 _16961_/X sky130_fd_sc_hd__mux2_2
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16624__267 _16626__269/A vssd1 vssd1 vccd1 vccd1 _19041_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18700_ _18700_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15912_ _17816_/Q _15938_/A vssd1 vssd1 vccd1 vccd1 _15913_/B sky130_fd_sc_hd__xor2_1
X_11035_ _11035_/A vssd1 vssd1 vccd1 vccd1 _18262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16892_ _16892_/A vssd1 vssd1 vccd1 vccd1 _16892_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_231_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18631_ _18631_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15843_ _15843_/A vssd1 vssd1 vccd1 vccd1 _15843_/X sky130_fd_sc_hd__buf_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03180_ clkbuf_0__03180_/X vssd1 vssd1 vccd1 vccd1 _14440__607/A sky130_fd_sc_hd__clkbuf_16
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18562_ _18562_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _17956_/Q _17681_/Q _12993_/S vssd1 vssd1 vccd1 vccd1 _12987_/B sky130_fd_sc_hd__mux2_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17513_ _17513_/CLK _17513_/D vssd1 vssd1 vccd1 vccd1 _17513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14725_ _18410_/Q _18402_/Q _19315_/Q _17719_/Q _14641_/A _14546_/X vssd1 vssd1 vccd1
+ vccd1 _14725_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11937_ _17780_/Q vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _18493_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17444_ _17444_/A vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11868_ _11868_/A vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__clkbuf_1
X_14656_ _14673_/S _14649_/Y _14651_/Y _14653_/Y _14655_/Y vssd1 vssd1 vccd1 vccd1
+ _14656_/X sky130_fd_sc_hd__o32a_1
XFILLER_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13607_ _13441_/X _13601_/X _13606_/Y _13604_/X vssd1 vssd1 vccd1 vccd1 _17846_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _18361_/Q _10794_/X _10825_/S vssd1 vssd1 vccd1 vccd1 _10820_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17375_ _19288_/Q _17489_/B vssd1 vssd1 vccd1 vccd1 _17377_/C sky130_fd_sc_hd__xnor2_1
X_14496__652 _14496__652/A vssd1 vssd1 vccd1 vccd1 _18287_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11799_ _13168_/A vssd1 vssd1 vccd1 vccd1 _16689_/A sky130_fd_sc_hd__buf_4
X_14587_ _08857_/X _14244_/X _14095_/A vssd1 vssd1 vccd1 vccd1 _16536_/C sky130_fd_sc_hd__a21oi_2
XFILLER_229_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19114_ _19114_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13538_ _17825_/Q vssd1 vssd1 vccd1 vccd1 _15927_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19045_ _19045_/CLK _19045_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_16257_ _16257_/A _16257_/B vssd1 vssd1 vccd1 vccd1 _16257_/Y sky130_fd_sc_hd__nor2_1
X_13469_ _13469_/A vssd1 vssd1 vccd1 vccd1 _17803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15208_ _15208_/A vssd1 vssd1 vccd1 vccd1 _15273_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16188_ _10391_/X _16177_/X _16187_/Y _16164_/X vssd1 vssd1 vccd1 vccd1 _16188_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880__363 _11881__364/A vssd1 vssd1 vccd1 vccd1 _17510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_173_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _09826_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09716_/S sky130_fd_sc_hd__or2_2
XFILLER_96_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09631_ _09631_/A vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__buf_4
XFILLER_56_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18829_ _18829_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _10310_/A _10967_/A vssd1 vssd1 vccd1 vccd1 _09578_/S sky130_fd_sc_hd__nor2_2
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09493_ _19009_/Q _09492_/X _09496_/S vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__05079_ _17397_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05079_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14397__572 _14399__574/A vssd1 vssd1 vccd1 vccd1 _18207_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09829_ _09829_/A vssd1 vssd1 vccd1 vccd1 _18819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12840_ _12840_/A vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__buf_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12764_/Y _12766_/Y _12769_/Y _12770_/Y _12568_/A _12469_/S vssd1 vssd1 vccd1
+ vccd1 _12850_/A sky130_fd_sc_hd__mux4_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04585_ clkbuf_0__04585_/X vssd1 vssd1 vccd1 vccd1 _16700__324/A sky130_fd_sc_hd__clkbuf_16
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A vssd1 vssd1 vccd1 vccd1 _11722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_215_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _18654_/Q _15490_/B vssd1 vssd1 vccd1 vccd1 _15528_/C sky130_fd_sc_hd__xnor2_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14818__747 _14818__747/A vssd1 vssd1 vccd1 vccd1 _18390_/CLK sky130_fd_sc_hd__inv_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _08804_/X _17532_/Q _11653_/S vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__mux2_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ _10112_/X _18452_/Q _10612_/S vssd1 vssd1 vccd1 vccd1 _10605_/A sky130_fd_sc_hd__mux2_1
X_17160_ _17158_/X _17189_/B _17160_/C vssd1 vssd1 vccd1 vccd1 _17161_/A sky130_fd_sc_hd__and3b_1
X_11584_ _11599_/S vssd1 vssd1 vccd1 vccd1 _11593_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _13274_/X _13311_/A _13320_/X vssd1 vssd1 vccd1 vccd1 _13323_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03398_ clkbuf_0__03398_/X vssd1 vssd1 vccd1 vccd1 _14758__699/A sky130_fd_sc_hd__clkbuf_16
X_16111_ _16276_/A vssd1 vssd1 vccd1 vccd1 _16223_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ _10535_/A vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__clkbuf_1
X_17091_ _12206_/A _17089_/X _17090_/X _13346_/B vssd1 vssd1 vccd1 vccd1 _17091_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ _13173_/X _13253_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _13254_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16042_ _15812_/Y _15958_/B _16044_/B vssd1 vssd1 vccd1 vccd1 _16042_/Y sky130_fd_sc_hd__a21oi_1
X_10466_ _18543_/Q _10342_/X _10466_/S vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12205_ _12205_/A vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__buf_2
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13212_/B vssd1 vssd1 vccd1 vccd1 _13208_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__04019_ clkbuf_0__04019_/X vssd1 vssd1 vccd1 vccd1 _15893__182/A sky130_fd_sc_hd__clkbuf_16
X_10397_ _16195_/A vssd1 vssd1 vccd1 vccd1 _16172_/A sky130_fd_sc_hd__buf_2
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18455_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_16329__226 _16329__226/A vssd1 vssd1 vccd1 vccd1 _18942_/CLK sky130_fd_sc_hd__inv_2
XFILLER_233_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ _17518_/Q _17733_/Q _12136_/S vssd1 vssd1 vccd1 vccd1 _12137_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ _18021_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03401_ _14771_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03401_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ _11933_/X _11935_/X _12067_/S vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__mux2_1
X_16944_ _16963_/A _16944_/B vssd1 vssd1 vccd1 vccd1 _16944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_97_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18993_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_238_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ _09047_/X _18269_/Q _11022_/S vssd1 vssd1 vccd1 vccd1 _11019_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _17737_/CLK sky130_fd_sc_hd__clkbuf_16
X_16875_ _16866_/X _16874_/X _16875_/S vssd1 vssd1 vccd1 vccd1 _16875_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18614_ _18614_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03163_ clkbuf_0__03163_/X vssd1 vssd1 vccd1 vccd1 _14374_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15867__164 _15867__164/A vssd1 vssd1 vccd1 vccd1 _18839_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03194_ _14511_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03194_/X sky130_fd_sc_hd__clkbuf_16
X_18545_ _18545_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03094_ clkbuf_0__03094_/X vssd1 vssd1 vccd1 vccd1 _14256_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12969_ _12957_/X _12969_/B vssd1 vssd1 vccd1 vccd1 _12970_/A sky130_fd_sc_hd__and2b_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _18369_/Q _18321_/Q _18377_/Q _17710_/Q _14599_/X _14627_/X vssd1 vssd1 vccd1
+ vccd1 _14708_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18476_ _18477_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17427_ _17427_/A vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ _14679_/A _14639_/B vssd1 vssd1 vccd1 vccd1 _14639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17358_ _17356_/X _17358_/B vssd1 vssd1 vccd1 vccd1 _17359_/A sky130_fd_sc_hd__and2b_1
XFILLER_146_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16309_ _16315_/A vssd1 vssd1 vccd1 vccd1 _16309_/X sky130_fd_sc_hd__buf_1
XFILLER_158_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15424__920 _15425__921/A vssd1 vssd1 vccd1 vccd1 _18607_/CLK sky130_fd_sc_hd__inv_2
X_17289_ _17289_/A _17289_/B _17289_/C vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__and3_1
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19028_ _19037_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08993_ _18802_/Q vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04579_ _16683_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04579_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_60_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09614_ _09614_/A _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__and3_1
XFILLER_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09545_ _09560_/S vssd1 vssd1 vccd1 vccd1 _09554_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09476_ _09476_/A _09480_/A vssd1 vssd1 vccd1 vccd1 _09477_/B sky130_fd_sc_hd__or2_1
XFILLER_212_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04370_ clkbuf_0__04370_/X vssd1 vssd1 vccd1 vccd1 _16326__224/A sky130_fd_sc_hd__clkbuf_16
XFILLER_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03183_ clkbuf_0__03183_/X vssd1 vssd1 vccd1 vccd1 _14455__619/A sky130_fd_sc_hd__clkbuf_16
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ _09688_/X _18604_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10251_/A vssd1 vssd1 vccd1 vccd1 _18635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10182_ _10182_/A vssd1 vssd1 vccd1 vccd1 _18693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14990_ _14990_/A vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447__613 _14447__613/A vssd1 vssd1 vccd1 vccd1 _18248_/CLK sky130_fd_sc_hd__inv_2
X_13941_ _17958_/Q _13941_/B vssd1 vssd1 vccd1 vccd1 _13941_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13872_ _17935_/Q _13863_/B _13871_/Y _13868_/X vssd1 vssd1 vccd1 vccd1 _17935_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _15611_/A _15615_/C _15611_/C vssd1 vssd1 vccd1 vccd1 _15611_/X sky130_fd_sc_hd__or3_1
X_12823_ _12812_/X _12823_/B vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__and2b_1
XFILLER_216_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16591_ _19025_/Q _16593_/C _16564_/X vssd1 vssd1 vccd1 vccd1 _16591_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18330_ _18996_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15542_ _15624_/A _15542_/B vssd1 vssd1 vccd1 vccd1 _18643_/D sky130_fd_sc_hd__nor2_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12758_/B _12758_/C _12758_/D vssd1 vssd1 vccd1 vccd1 _12755_/C sky130_fd_sc_hd__nand3_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04568_ clkbuf_0__04568_/X vssd1 vssd1 vccd1 vccd1 _16632__274/A sky130_fd_sc_hd__clkbuf_16
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ _17926_/Q vssd1 vssd1 vccd1 vccd1 _13845_/A sky130_fd_sc_hd__inv_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18261_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 _18261_/Q sky130_fd_sc_hd__dfxtp_1
X_12685_ _12686_/B _12687_/A _12684_/Y vssd1 vssd1 vccd1 vccd1 _17613_/D sky130_fd_sc_hd__a21oi_1
XFILLER_163_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15473_ _17839_/Q _15516_/B vssd1 vssd1 vccd1 vccd1 _15517_/B sky130_fd_sc_hd__or2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17210_/X _17235_/B _17212_/C vssd1 vssd1 vccd1 vccd1 _17213_/A sky130_fd_sc_hd__and3b_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _11636_/A vssd1 vssd1 vccd1 vccd1 _17540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18192_ _18192_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
X_17143_ _17142_/B _17142_/C _17142_/A vssd1 vssd1 vccd1 vccd1 _17144_/C sky130_fd_sc_hd__a21o_1
X_11567_ _17588_/Q _10887_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__mux2_1
X_14355_ _14355_/A vssd1 vssd1 vccd1 vccd1 _14355_/X sky130_fd_sc_hd__buf_1
XFILLER_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13306_ _17761_/Q _13303_/X _13305_/Y vssd1 vssd1 vccd1 vccd1 _17761_/D sky130_fd_sc_hd__o21a_1
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ _18520_/Q _10339_/X _10520_/S vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17074_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17074_/X sky130_fd_sc_hd__buf_1
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ _11498_/A vssd1 vssd1 vccd1 vccd1 _18046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13237_ _13783_/A vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__buf_4
X_16025_ _18873_/Q _16025_/B vssd1 vssd1 vccd1 vccd1 _16025_/Y sky130_fd_sc_hd__nand2_1
X_10449_ _10449_/A vssd1 vssd1 vccd1 vccd1 _18551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13168_ _13168_/A vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__buf_2
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12119_ _12116_/X _12117_/X _12118_/X _17777_/Q vssd1 vssd1 vccd1 vccd1 _17487_/B
+ sky130_fd_sc_hd__a22o_4
X_17976_ _18001_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_1
X_13099_ _11888_/X _13099_/B _13099_/C vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__and3b_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16927_ _16927_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_226_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ _09868_/X _16857_/X _16836_/X vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15157__865 _15158__866/A vssd1 vssd1 vccd1 vccd1 _18541_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15809_ _15809_/A vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03146_ clkbuf_0__03146_/X vssd1 vssd1 vccd1 vccd1 _14265__466/A sky130_fd_sc_hd__clkbuf_16
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ _16765_/X _16786_/Y _16788_/Y _14074_/A _16762_/A vssd1 vssd1 vccd1 vccd1
+ _16790_/B sky130_fd_sc_hd__o32a_1
XFILLER_53_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09330_ _19095_/Q _08958_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18528_ _18528_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03177_ _14419_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03177_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ _09261_/A vssd1 vssd1 vccd1 vccd1 _19127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18459_ _19039_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09192_ _19161_/Q _09130_/X _09196_/S vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03979_ clkbuf_0__03979_/X vssd1 vssd1 vccd1 vccd1 _15737__1025/A sky130_fd_sc_hd__clkbuf_16
XFILLER_174_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_15101__820 _15103__822/A vssd1 vssd1 vccd1 vccd1 _18496_/CLK sky130_fd_sc_hd__inv_2
X_08976_ _19218_/Q _08949_/X _08982_/S vssd1 vssd1 vccd1 vccd1 _08977_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09528_ _18966_/Q _09481_/X _09536_/S vssd1 vssd1 vccd1 vccd1 _09529_/A sky130_fd_sc_hd__mux2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _14580_/A vssd1 vssd1 vccd1 vccd1 _09459_/X sky130_fd_sc_hd__buf_4
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ _12470_/A vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__buf_4
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11421_ _11436_/S vssd1 vssd1 vccd1 vccd1 _11430_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_177_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ _11352_/A vssd1 vssd1 vccd1 vccd1 _18137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03166_ clkbuf_0__03166_/X vssd1 vssd1 vccd1 vccd1 _14373__554/A sky130_fd_sc_hd__clkbuf_16
XFILLER_152_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10303_ _10303_/A vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__clkbuf_1
X_14071_ _14071_/A vssd1 vssd1 vccd1 vccd1 _14083_/B sky130_fd_sc_hd__clkbuf_2
X_11283_ _18163_/Q _11282_/X _11283_/S vssd1 vssd1 vccd1 vccd1 _11284_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _16620_/A _13022_/B _13022_/C vssd1 vssd1 vccd1 vccd1 _13023_/A sky130_fd_sc_hd__and3b_1
Xclkbuf_1_0__f__03097_ clkbuf_0__03097_/X vssd1 vssd1 vccd1 vccd1 _14177__454/A sky130_fd_sc_hd__clkbuf_16
X_10234_ _18672_/Q _09764_/X hold3/X vssd1 vssd1 vccd1 vccd1 _10235_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17830_ _18919_/CLK _17830_/D vssd1 vssd1 vccd1 vccd1 _17830_/Q sky130_fd_sc_hd__dfxtp_1
X_10165_ _18699_/Q _10060_/X _10167_/S vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17761_ _19288_/CLK _17761_/D vssd1 vssd1 vccd1 vccd1 _17761_/Q sky130_fd_sc_hd__dfxtp_1
X_14973_ _14979_/C _15057_/A vssd1 vssd1 vccd1 vccd1 _14973_/Y sky130_fd_sc_hd__nand2_1
X_10096_ _18726_/Q _10048_/X _10104_/S vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16712_ _13066_/X _19109_/Q vssd1 vssd1 vccd1 vccd1 _16713_/A sky130_fd_sc_hd__and2b_1
X_13924_ _14053_/A _13945_/B vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__and2_2
X_17692_ _18007_/CLK _17692_/D vssd1 vssd1 vccd1 vccd1 _17692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13855_ _14243_/A _13855_/B _14076_/B vssd1 vssd1 vccd1 vccd1 _13867_/B sky130_fd_sc_hd__and3_1
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12806_ _12795_/X _12806_/B vssd1 vssd1 vccd1 vccd1 _12807_/A sky130_fd_sc_hd__and2b_1
X_16574_ _19019_/Q _16576_/C _16564_/X vssd1 vssd1 vccd1 vccd1 _16574_/Y sky130_fd_sc_hd__a21oi_1
X_13786_ _13786_/A vssd1 vssd1 vccd1 vccd1 _13786_/X sky130_fd_sc_hd__clkbuf_4
X_10998_ _18278_/Q _09136_/X _10998_/S vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18313_ _18313_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15525_ _15525_/A _15525_/B _15525_/C _15525_/D vssd1 vssd1 vccd1 vccd1 _15525_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12737_/A _12737_/B _12737_/C _12737_/D vssd1 vssd1 vccd1 vccd1 _12746_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19293_ _19293_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18244_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12668_ _17608_/Q _12665_/A _12663_/X vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__o21ai_1
XFILLER_176_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11619_ _11655_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11635_/S sky130_fd_sc_hd__nor2_2
X_18175_ _18175_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
X_12599_ _12603_/B _12759_/A _12599_/C vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__and3b_1
XFILLER_237_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ _17191_/A vssd1 vssd1 vccd1 vccd1 _17126_/X sky130_fd_sc_hd__buf_2
XFILLER_184_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14269_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14269_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__03795_ _15392_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03795_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_98_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16008_ _16024_/A _16008_/B _16018_/C vssd1 vssd1 vccd1 vccd1 _16008_/X sky130_fd_sc_hd__or3_1
XFILLER_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_41_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _18994_/Q vssd1 vssd1 vccd1 vccd1 _08830_/X sky130_fd_sc_hd__buf_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08757_/X _08761_/B vssd1 vssd1 vccd1 vccd1 _08761_/X sky130_fd_sc_hd__and2b_1
XFILLER_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17959_ _17959_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _09313_/A vssd1 vssd1 vccd1 vccd1 _19103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09244_ _09244_/A vssd1 vssd1 vccd1 vccd1 _09244_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09175_ _09175_/A vssd1 vssd1 vccd1 vccd1 _19169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ _19270_/Q _08958_/X _08959_/S vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860__781 _14862__783/A vssd1 vssd1 vccd1 vccd1 _18426_/CLK sky130_fd_sc_hd__inv_2
XFILLER_217_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11970_ _12083_/A _12084_/A _12034_/A vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__mux2_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10921_ _18311_/Q _10898_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10922_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13640_ _13640_/A vssd1 vssd1 vccd1 vccd1 _17858_/D sky130_fd_sc_hd__clkbuf_1
X_10852_ _10867_/S vssd1 vssd1 vccd1 vccd1 _10861_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13571_ _13623_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _13589_/S sky130_fd_sc_hd__nor2_1
X_10783_ _18373_/Q _10707_/X _10787_/S vssd1 vssd1 vccd1 vccd1 _10784_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15310_ _19070_/Q _19062_/Q _19054_/Q _19008_/Q _15232_/X _15233_/X vssd1 vssd1 vccd1
+ vccd1 _15311_/A sky130_fd_sc_hd__mux4_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12520_/X _12521_/X _18008_/Q vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16286_/X _16289_/X _16290_/S vssd1 vssd1 vccd1 vccd1 _16291_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _16036_/B vssd1 vssd1 vccd1 vccd1 _16064_/A sky130_fd_sc_hd__clkbuf_2
X_12453_ _17622_/Q _17623_/Q _17624_/Q _17625_/Q _12436_/S _12464_/S vssd1 vssd1 vccd1
+ vccd1 _12453_/X sky130_fd_sc_hd__mux4_2
XFILLER_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11404_ _11321_/X _18114_/Q _11412_/S vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__mux2_1
X_12384_ _17602_/Q vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14490__647 _14490__647/A vssd1 vssd1 vccd1 vccd1 _18282_/CLK sky130_fd_sc_hd__inv_2
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ _16570_/A vssd1 vssd1 vccd1 vccd1 _14123_/X sky130_fd_sc_hd__clkbuf_2
X_11335_ _11335_/A vssd1 vssd1 vccd1 vccd1 _11335_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108__826 _15109__827/A vssd1 vssd1 vccd1 vccd1 _18502_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03149_ clkbuf_0__03149_/X vssd1 vssd1 vccd1 vccd1 _14286__484/A sky130_fd_sc_hd__clkbuf_16
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18931_ _18931_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_2
X_14054_ _14055_/A vssd1 vssd1 vccd1 vccd1 _14054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11266_ _11266_/A vssd1 vssd1 vccd1 vccd1 _18169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _17681_/Q _12835_/A _12834_/A _17671_/Q _13004_/X vssd1 vssd1 vccd1 vccd1
+ _13005_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _18679_/Q _09767_/X hold6/X vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18862_ _18889_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_1
X_11197_ _11197_/A vssd1 vssd1 vccd1 vccd1 _18198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17813_ _19339_/CLK _17813_/D vssd1 vssd1 vccd1 vccd1 _17813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _10148_/A vssd1 vssd1 vccd1 vccd1 _18707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18793_ _18793_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _19336_/CLK _17744_/D vssd1 vssd1 vccd1 vccd1 _17744_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14956_ _14960_/A _14963_/A _14956_/C vssd1 vssd1 vccd1 vccd1 _14957_/C sky130_fd_sc_hd__or3_1
X_10079_ _10079_/A vssd1 vssd1 vccd1 vccd1 _18734_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__05081_ clkbuf_0__05081_/X vssd1 vssd1 vccd1 vccd1 _17414__104/A sky130_fd_sc_hd__clkbuf_16
XFILLER_48_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14384__563 _14385__564/A vssd1 vssd1 vccd1 vccd1 _18198_/CLK sky130_fd_sc_hd__inv_2
X_13907_ _17945_/Q _13902_/X _13906_/Y vssd1 vssd1 vccd1 vccd1 _17945_/D sky130_fd_sc_hd__o21a_1
XFILLER_223_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17675_ _19037_/CLK _17675_/D vssd1 vssd1 vccd1 vccd1 _17675_/Q sky130_fd_sc_hd__dfxtp_1
X_17073__59 _17073__59/A vssd1 vssd1 vccd1 vccd1 _19208_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_201 _16715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_212 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_223 _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13838_ input58/X _13847_/B vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__and2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19345_ _19345_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
X_13769_ _13769_/A _13795_/B vssd1 vssd1 vccd1 vccd1 _13778_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15508_ _17837_/Q _15511_/A vssd1 vssd1 vccd1 vccd1 _15509_/B sky130_fd_sc_hd__xnor2_1
X_19276_ _19340_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16488_ _16498_/A _16488_/B _16491_/B vssd1 vssd1 vccd1 vccd1 _16488_/X sky130_fd_sc_hd__or3_1
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18227_ _18227_/CLK _18227_/D vssd1 vssd1 vccd1 vccd1 _18227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18158_ _18158_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 _18158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17109_ _17109_/A _17109_/B vssd1 vssd1 vccd1 vccd1 _17114_/A sky130_fd_sc_hd__and2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14391__567 _14391__567/A vssd1 vssd1 vccd1 vccd1 _18202_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18089_ _18870_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _09931_/A vssd1 vssd1 vccd1 vccd1 _18784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348__240 _16349__241/A vssd1 vssd1 vccd1 vccd1 _18956_/CLK sky130_fd_sc_hd__inv_2
X_15709__1003 _15710__1004/A vssd1 vssd1 vccd1 vccd1 _18720_/CLK sky130_fd_sc_hd__inv_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _15808_/B vssd1 vssd1 vccd1 vccd1 _09895_/C sky130_fd_sc_hd__clkbuf_2
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08813_ _08828_/S vssd1 vssd1 vccd1 vccd1 _08822_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12239__383 _12239__383/A vssd1 vssd1 vccd1 vccd1 _17547_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09793_ _09793_/A vssd1 vssd1 vccd1 vccd1 _18835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _18068_/Q _18074_/Q _18075_/Q _13130_/B vssd1 vssd1 vccd1 vccd1 _11787_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_227_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120__423 _13120__423/A vssd1 vssd1 vccd1 vccd1 _17719_/CLK sky130_fd_sc_hd__inv_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14285__483 _14286__484/A vssd1 vssd1 vccd1 vccd1 _18118_/CLK sky130_fd_sc_hd__inv_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ _10049_/A _10075_/B _10437_/B vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__or3b_4
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09158_ _19176_/Q _09100_/X _09160_/S vssd1 vssd1 vccd1 vccd1 _09159_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09089_ _19195_/Q _09080_/X _09105_/S vssd1 vssd1 vccd1 vccd1 _09090_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15893__182 _15893__182/A vssd1 vssd1 vccd1 vccd1 _18858_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _18228_/Q _11062_/X _11122_/S vssd1 vssd1 vccd1 vccd1 _11121_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _18256_/Q _11050_/X _11057_/S vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ _18763_/Q _09951_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14741_ _14544_/X _14730_/X _14740_/Y vssd1 vssd1 vccd1 vccd1 _14741_/X sky130_fd_sc_hd__a21o_1
XFILLER_229_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11953_ _11949_/X _11950_/X _11977_/S vssd1 vssd1 vccd1 vccd1 _11953_/X sky130_fd_sc_hd__mux2_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17454_/X _17460_/B vssd1 vssd1 vccd1 vccd1 _17461_/A sky130_fd_sc_hd__and2b_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _18989_/Q vssd1 vssd1 vccd1 vccd1 _10904_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14670_/X _14671_/X _14726_/S vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__mux2_1
X_16411_ _16411_/A _16411_/B _16411_/C _16410_/X vssd1 vssd1 vccd1 vccd1 _16417_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_233_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13623_ _13623_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13642_/S sky130_fd_sc_hd__nor2_1
X_10835_ _18354_/Q _10789_/X _10843_/S vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__mux2_1
X_17391_ _17415_/A vssd1 vssd1 vccd1 vccd1 _17391_/X sky130_fd_sc_hd__buf_1
XFILLER_220_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19130_ _19132_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13554_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13636_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10766_ _18380_/Q _10710_/X _10768_/S vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _12447_/X _12438_/X _12765_/S vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__mux2_1
X_19061_ _19061_/CLK _19061_/D vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16273_ _16190_/X _16264_/X _16272_/Y _16214_/X vssd1 vssd1 vccd1 vccd1 _16273_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10697_ _10697_/A vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__clkbuf_1
X_13485_ _13560_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__or2_1
XFILLER_201_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18012_ _18012_/CLK _18012_/D vssd1 vssd1 vccd1 vccd1 _18012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _16294_/C _15955_/A vssd1 vssd1 vccd1 vccd1 _15267_/A sky130_fd_sc_hd__nand2_2
X_12436_ _12383_/X _17602_/Q _12436_/S vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03601_ clkbuf_0__03601_/X vssd1 vssd1 vccd1 vccd1 _15165__872/A sky130_fd_sc_hd__clkbuf_16
X_15155_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__buf_1
X_12367_ _18011_/Q vssd1 vssd1 vccd1 vccd1 _12487_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106_ _13786_/A _14099_/X _14096_/X vssd1 vssd1 vccd1 vccd1 _14106_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _11318_/A vssd1 vssd1 vccd1 vccd1 _18148_/D sky130_fd_sc_hd__clkbuf_1
X_12298_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12298_/X sky130_fd_sc_hd__clkbuf_2
X_15086_ _15086_/A vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__buf_1
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14867__787 _14869__789/A vssd1 vssd1 vccd1 vccd1 _18432_/CLK sky130_fd_sc_hd__inv_2
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14037_ _13400_/A _14033_/X _14034_/X vssd1 vssd1 vccd1 vccd1 _14037_/Y sky130_fd_sc_hd__a21oi_1
X_18914_ _18919_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
X_11249_ _11153_/X _18175_/Q _11251_/S vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18845_ _18845_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18776_ _18776_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15988_ _15986_/X _15987_/Y _15982_/X vssd1 vssd1 vccd1 vccd1 _18866_/D sky130_fd_sc_hd__a21oi_1
XFILLER_83_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17727_ _17878_/CLK _17727_/D vssd1 vssd1 vccd1 vccd1 _17727_/Q sky130_fd_sc_hd__dfxtp_1
X_14939_ _18461_/Q _14939_/B vssd1 vssd1 vccd1 vccd1 _14961_/A sky130_fd_sc_hd__xor2_1
XFILLER_247_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__04015_ clkbuf_0__04015_/X vssd1 vssd1 vccd1 vccd1 _15882__176/A sky130_fd_sc_hd__clkbuf_16
X_17658_ _17969_/CLK _17658_/D vssd1 vssd1 vccd1 vccd1 _17658_/Q sky130_fd_sc_hd__dfxtp_1
X_16716__333 _16717__334/A vssd1 vssd1 vccd1 vccd1 _19112_/CLK sky130_fd_sc_hd__inv_2
XFILLER_247_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16609_ _19033_/Q _16607_/B _16608_/Y vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17589_ _18010_/CLK _17589_/D vssd1 vssd1 vccd1 vccd1 _17589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19328_ _19329_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19259_ _19261_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _18802_/Q _18807_/Q vssd1 vssd1 vccd1 vccd1 _09857_/C sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__04848_ clkbuf_0__04848_/X vssd1 vssd1 vccd1 vccd1 _17067__54/A sky130_fd_sc_hd__clkbuf_16
XFILLER_145_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _09914_/A vssd1 vssd1 vccd1 vccd1 _18791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09845_ _16892_/A vssd1 vssd1 vccd1 vccd1 _09845_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09776_ _09776_/A vssd1 vssd1 vccd1 vccd1 _18842_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _13128_/A _11779_/A vssd1 vssd1 vccd1 vccd1 _14243_/C sky130_fd_sc_hd__and2b_1
XFILLER_233_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441__608 _14442__609/A vssd1 vssd1 vccd1 vccd1 _18243_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ _10620_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10636_/S sky130_fd_sc_hd__nor2_2
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10551_/A vssd1 vssd1 vccd1 vccd1 _18506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13270_ _17750_/Q _13253_/X _13269_/Y vssd1 vssd1 vccd1 vccd1 _17750_/D sky130_fd_sc_hd__o21a_1
X_10482_ _18536_/Q _10339_/X _10484_/S vssd1 vssd1 vccd1 vccd1 _10483_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ _12152_/A vssd1 vssd1 vccd1 vccd1 _17522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11103_ _11103_/A vssd1 vssd1 vccd1 vccd1 _18236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12083_ _12083_/A vssd1 vssd1 vccd1 vccd1 _12083_/Y sky130_fd_sc_hd__clkinv_2
X_16960_ _16958_/X _16959_/X _16979_/S vssd1 vssd1 vccd1 vccd1 _16960_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15911_ _17817_/Q _15937_/B vssd1 vssd1 vccd1 vccd1 _15938_/A sky130_fd_sc_hd__or2_1
X_11034_ _18262_/Q _09136_/X _11034_/S vssd1 vssd1 vccd1 vccd1 _11035_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16891_ _19139_/Q _16797_/X _16890_/X _15628_/X vssd1 vssd1 vccd1 vccd1 _19139_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_238_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15671__972 _15671__972/A vssd1 vssd1 vccd1 vccd1 _18689_/CLK sky130_fd_sc_hd__inv_2
XFILLER_209_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18630_ _18630_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _18561_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15773_ _15779_/A vssd1 vssd1 vccd1 vccd1 _15773_/X sky130_fd_sc_hd__buf_1
X_12985_ _12985_/A vssd1 vssd1 vccd1 vccd1 _17680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17512_ _17512_/CLK _17512_/D vssd1 vssd1 vccd1 vccd1 _17512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _19179_/Q _19171_/Q _19203_/Q _18338_/Q _14594_/X _14595_/X vssd1 vssd1 vccd1
+ vccd1 _14724_/X sky130_fd_sc_hd__mux4_1
X_11936_ _19228_/Q _19229_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__mux2_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _18492_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17443_ _17437_/X _17443_/B vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__and2b_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14655_ _14651_/A _14654_/X _14673_/S vssd1 vssd1 vccd1 vccd1 _14655_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11867_ _17928_/Q _17843_/Q vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__or2_4
X_17051__40 _17053__42/A vssd1 vssd1 vccd1 vccd1 _19189_/CLK sky130_fd_sc_hd__inv_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13606_ _17846_/Q _13608_/B vssd1 vssd1 vccd1 vccd1 _13606_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17374_ _19287_/Q _17492_/B vssd1 vssd1 vccd1 vccd1 _17377_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10818_ _10818_/A vssd1 vssd1 vccd1 vccd1 _18362_/D sky130_fd_sc_hd__clkbuf_1
X_14586_ _14544_/X _14560_/X _14585_/Y vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__a21o_1
X_15708__1002 _15710__1004/A vssd1 vssd1 vccd1 vccd1 _18719_/CLK sky130_fd_sc_hd__inv_2
X_11798_ _19145_/Q _11826_/A vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__and2_1
XFILLER_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14873__791 _14873__791/A vssd1 vssd1 vccd1 vccd1 _18436_/CLK sky130_fd_sc_hd__inv_2
X_19113_ _19113_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13537_ _16522_/A _13523_/X _13526_/X _17824_/Q _15083_/B vssd1 vssd1 vccd1 vccd1
+ _17824_/D sky130_fd_sc_hd__a221o_1
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10749_ _10749_/A vssd1 vssd1 vccd1 vccd1 _18388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19044_ _19044_/CLK _19044_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
X_16256_ _18530_/Q _18538_/Q _18546_/Q _18554_/Q _10420_/A _16117_/X vssd1 vssd1 vccd1
+ vccd1 _16257_/B sky130_fd_sc_hd__mux4_2
X_13468_ _13560_/A _13468_/B vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__or2_1
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12419_ _12432_/S vssd1 vssd1 vccd1 vccd1 _12555_/A sky130_fd_sc_hd__buf_2
X_16187_ _16234_/A _16187_/B vssd1 vssd1 vccd1 vccd1 _16187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13399_ _13414_/B vssd1 vssd1 vccd1 vccd1 _13405_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15069_ _16057_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _18476_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _18931_/D sky130_fd_sc_hd__nor2_1
X_18828_ _18828_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _09561_/A vssd1 vssd1 vccd1 vccd1 _18951_/D sky130_fd_sc_hd__clkbuf_1
X_18759_ _18759_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ _18884_/Q vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__05078_ _17391_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05078_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_3_0_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09828_ _09674_/X _18819_/Q _09836_/S vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09759_ _18847_/Q _09758_/X _09759_/S vssd1 vssd1 vccd1 vccd1 _09760_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ _12770_/A vssd1 vssd1 vccd1 vccd1 _12770_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11721_ _17910_/Q _11720_/X _11869_/B vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__mux2_8
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A vssd1 vssd1 vccd1 vccd1 _17533_/D sky130_fd_sc_hd__clkbuf_1
X_15150__860 _15154__864/A vssd1 vssd1 vccd1 vccd1 _18536_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10603_ _10618_/S vssd1 vssd1 vccd1 vccd1 _10612_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11583_ _11601_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11599_/S sky130_fd_sc_hd__nor2_2
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03397_ clkbuf_0__03397_/X vssd1 vssd1 vccd1 vccd1 _14752__694/A sky130_fd_sc_hd__clkbuf_16
X_16110_ _16171_/A _16110_/B vssd1 vssd1 vccd1 vccd1 _16110_/Y sky130_fd_sc_hd__nor2_1
X_13322_ _17767_/Q _13304_/X _13321_/Y vssd1 vssd1 vccd1 vccd1 _17767_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16630__272 _16631__273/A vssd1 vssd1 vccd1 vccd1 _19046_/CLK sky130_fd_sc_hd__inv_2
X_17090_ _17775_/Q _11947_/A vssd1 vssd1 vccd1 vccd1 _17090_/X sky130_fd_sc_hd__or2b_1
X_14298__493 _14299__494/A vssd1 vssd1 vccd1 vccd1 _18128_/CLK sky130_fd_sc_hd__inv_2
X_10534_ _18513_/Q _10336_/X _10538_/S vssd1 vssd1 vccd1 vccd1 _10535_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16041_ _16063_/B _16040_/Y _15955_/A vssd1 vssd1 vccd1 vccd1 _16050_/A sky130_fd_sc_hd__a21o_1
X_13253_ _13259_/A vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__clkbuf_2
X_10465_ _10465_/A vssd1 vssd1 vccd1 vccd1 _18544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _12204_/A vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13184_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13184_/X sky130_fd_sc_hd__buf_6
X_10396_ _18565_/Q vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__buf_4
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12135_ _12135_/A vssd1 vssd1 vccd1 vccd1 _17517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17992_ _18021_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03400_ _14765_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03400_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16943_ _18248_/Q _18240_/Q _18232_/Q _18224_/Q _16849_/X _16850_/X vssd1 vssd1 vccd1
+ vccd1 _16944_/B sky130_fd_sc_hd__mux4_2
X_12066_ _17117_/C _17117_/B _19222_/Q _19223_/Q _11961_/X _11957_/S vssd1 vssd1 vccd1
+ vccd1 _12066_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14760__700 _14764__704/A vssd1 vssd1 vccd1 vccd1 _18343_/CLK sky130_fd_sc_hd__inv_2
X_11017_ _11017_/A vssd1 vssd1 vccd1 vccd1 _18270_/D sky130_fd_sc_hd__clkbuf_1
X_16874_ _16869_/X _16872_/X _16976_/S vssd1 vssd1 vccd1 vccd1 _16874_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18613_ _18613_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03162_ clkbuf_0__03162_/X vssd1 vssd1 vccd1 vccd1 _14354__539/A sky130_fd_sc_hd__clkbuf_16
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16672__306 _16674__308/A vssd1 vssd1 vccd1 vccd1 _19080_/CLK sky130_fd_sc_hd__inv_2
XFILLER_218_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03193_ _14505_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03193_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _18544_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_1
X_12968_ _17961_/Q _17676_/Q _12976_/S vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03093_ clkbuf_0__03093_/X vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_66_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17959_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14707_ _14705_/X _14706_/X _14726_/S vssd1 vssd1 vccd1 vccd1 _14707_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11919_ _19231_/Q vssd1 vssd1 vccd1 vccd1 _17159_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18475_ _18477_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _17973_/Q _17663_/Q _12908_/S vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17356_/X _17426_/B vssd1 vssd1 vccd1 vccd1 _17427_/A sky130_fd_sc_hd__and2b_1
X_14638_ _17583_/Q _18381_/Q _18389_/Q _18423_/Q _14554_/X _14637_/X vssd1 vssd1 vccd1
+ vccd1 _14639_/B sky130_fd_sc_hd__mux4_1
XFILLER_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _17753_/Q _19290_/Q _17357_/S vssd1 vssd1 vccd1 vccd1 _17358_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14569_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14569_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16308_ _16308_/A vssd1 vssd1 vccd1 vccd1 _16308_/X sky130_fd_sc_hd__buf_1
X_17288_ _19265_/Q _17288_/B _17288_/C _17288_/D vssd1 vssd1 vccd1 vccd1 _17289_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_173_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19027_ _19027_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17422__5 _17502__9/A vssd1 vssd1 vccd1 vccd1 _19323_/CLK sky130_fd_sc_hd__inv_2
X_16239_ _18598_/Q _18614_/Q _18740_/Q _18521_/Q _16195_/X _16138_/X vssd1 vssd1 vccd1
+ vccd1 _16240_/B sky130_fd_sc_hd__mux4_1
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15678__978 _15679__979/A vssd1 vssd1 vccd1 vccd1 _18695_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ hold26/X vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_248_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04578_ _16677_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04578_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09613_ _09613_/A _18922_/Q _16294_/C vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__and3_1
XFILLER_244_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09544_ _09826_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _09560_/S sky130_fd_sc_hd__or2_2
XFILLER_225_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09475_ _10770_/C _09467_/B _09464_/Y vssd1 vssd1 vccd1 vccd1 _19043_/D sky130_fd_sc_hd__o21a_1
XFILLER_211_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03182_ clkbuf_0__03182_/X vssd1 vssd1 vccd1 vccd1 _14474_/A sky130_fd_sc_hd__clkbuf_16
X_16729__343 _16730__344/A vssd1 vssd1 vccd1 vccd1 _19122_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10250_ _18635_/Q _10192_/X _10254_/S vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _18693_/Q _10180_/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15707__1001 _15707__1001/A vssd1 vssd1 vccd1 vccd1 _18718_/CLK sky130_fd_sc_hd__inv_2
X_13940_ _13155_/X _13929_/B _13939_/Y _13937_/X vssd1 vssd1 vccd1 vccd1 _17957_/D
+ sky130_fd_sc_hd__a211oi_1
X_14824__752 _14824__752/A vssd1 vssd1 vccd1 vccd1 _18395_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13871_ _13871_/A _13871_/B vssd1 vssd1 vccd1 vccd1 _13871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15610_ _18656_/Q _15610_/B vssd1 vssd1 vccd1 vccd1 _15611_/C sky130_fd_sc_hd__nor2_1
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12822_ _17649_/Q _17986_/Q _12822_/S vssd1 vssd1 vccd1 vccd1 _12823_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16590_ _19024_/Q _16587_/B _16589_/Y vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15541_ _18643_/Q _15612_/B _15540_/Y _15551_/A vssd1 vssd1 vccd1 vccd1 _15542_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12753_ _12758_/C _12747_/A _12758_/B vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__a21o_1
XFILLER_199_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11704_ _11704_/A vssd1 vssd1 vccd1 vccd1 _11704_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18260_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ _17842_/Q _17841_/Q _17840_/Q vssd1 vssd1 vccd1 vccd1 _15516_/B sky130_fd_sc_hd__or3_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12684_ _12686_/B _12687_/A _12607_/X vssd1 vssd1 vccd1 vccd1 _12684_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17209_/B _17210_/A _19245_/Q vssd1 vssd1 vccd1 vccd1 _17212_/C sky130_fd_sc_hd__a21o_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _17540_/Q _09697_/A _11635_/S vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__mux2_1
X_18191_ _18191_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
X_16335__231 _16337__233/A vssd1 vssd1 vccd1 vccd1 _18947_/CLK sky130_fd_sc_hd__inv_2
XFILLER_168_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17142_ _17142_/A _17142_/B _17142_/C vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__and3_1
XFILLER_128_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11566_ _11581_/S vssd1 vssd1 vccd1 vccd1 _11575_/S sky130_fd_sc_hd__clkbuf_2
X_14454__618 _14455__619/A vssd1 vssd1 vccd1 vccd1 _18253_/CLK sky130_fd_sc_hd__inv_2
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _13173_/X _13304_/X _13293_/X vssd1 vssd1 vccd1 vccd1 _13305_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_155_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10517_ _10517_/A vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ _18046_/Q _11326_/A _11503_/S vssd1 vssd1 vccd1 vccd1 _11498_/A sky130_fd_sc_hd__mux2_1
X_16024_ _16024_/A _16024_/B _16024_/C vssd1 vssd1 vccd1 vccd1 _16024_/X sky130_fd_sc_hd__or3_1
X_13236_ _17740_/Q _13218_/X _13235_/Y vssd1 vssd1 vccd1 vccd1 _17740_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ _10126_/X _18551_/Q _10448_/S vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13167_ _13147_/B _13165_/X _13166_/Y _13158_/X vssd1 vssd1 vccd1 vccd1 _17728_/D
+ sky130_fd_sc_hd__a211oi_1
X_10379_ _10379_/A vssd1 vssd1 vccd1 vccd1 _18582_/D sky130_fd_sc_hd__clkbuf_1
X_12118_ _11994_/X _11997_/X _12005_/X _11996_/X _17778_/Q _12111_/S vssd1 vssd1 vccd1
+ vccd1 _12118_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17975_ _18001_/CLK _17975_/D vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_1
X_13098_ _13087_/X _13088_/X _13097_/X _17703_/Q vssd1 vssd1 vccd1 vccd1 _13099_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_46_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ _12045_/X _12047_/X _12069_/A vssd1 vssd1 vccd1 vccd1 _17098_/A sky130_fd_sc_hd__mux2_1
X_16926_ _18207_/Q _18127_/Q _19184_/Q _18255_/Q _16822_/X _16823_/X vssd1 vssd1 vccd1
+ vccd1 _16927_/B sky130_fd_sc_hd__mux4_1
X_16342__235 _16344__237/A vssd1 vssd1 vccd1 vccd1 _18951_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14348__534 _14348__534/A vssd1 vssd1 vccd1 vccd1 _18169_/CLK sky130_fd_sc_hd__inv_2
X_15196__882 _15198__884/A vssd1 vssd1 vccd1 vccd1 _18561_/CLK sky130_fd_sc_hd__inv_2
XFILLER_238_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16857_ _18212_/Q _18196_/Q _18485_/Q _18188_/Q _16834_/X _09875_/X vssd1 vssd1 vccd1
+ vccd1 _16857_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _18641_/Q _15808_/B _15808_/C _17826_/Q vssd1 vssd1 vccd1 vccd1 _15809_/A
+ sky130_fd_sc_hd__and4b_1
Xclkbuf_1_1__f__03145_ clkbuf_0__03145_/X vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__clkbuf_16
X_12233__378 _12234__379/A vssd1 vssd1 vccd1 vccd1 _17542_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16788_ _16788_/A _16788_/B vssd1 vssd1 vccd1 vccd1 _16788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18527_ _18527_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03176_ _14418_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03176_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16637__278 _16638__279/A vssd1 vssd1 vccd1 vccd1 _19052_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _19127_/Q _09223_/X _09272_/S vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18458_ _19039_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17409_ _17409_/A vssd1 vssd1 vccd1 vccd1 _17409_/X sky130_fd_sc_hd__buf_1
X_09191_ _09191_/A vssd1 vssd1 vccd1 vccd1 _19162_/D sky130_fd_sc_hd__clkbuf_1
X_18389_ _18389_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_1
X_15387__890 _15389__892/A vssd1 vssd1 vccd1 vccd1 _18577_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03978_ clkbuf_0__03978_/X vssd1 vssd1 vccd1 vccd1 _15731__1020/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14767__706 _14768__707/A vssd1 vssd1 vccd1 vccd1 _18349_/CLK sky130_fd_sc_hd__inv_2
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ _08975_/A vssd1 vssd1 vccd1 vccd1 _19219_/D sky130_fd_sc_hd__clkbuf_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ _09542_/S vssd1 vssd1 vccd1 vccd1 _09536_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09458_ _14594_/A vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _09389_/A vssd1 vssd1 vccd1 vccd1 _19070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _11493_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11436_/S sky130_fd_sc_hd__nor2_2
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11351_ _18137_/Q _11264_/X _11357_/S vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03165_ clkbuf_0__03165_/X vssd1 vssd1 vccd1 vccd1 _14364__546/A sky130_fd_sc_hd__clkbuf_16
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ _18612_/Q _10189_/X _10302_/S vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__mux2_1
X_14070_ _14071_/A vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__buf_2
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _18661_/Q vssd1 vssd1 vccd1 vccd1 _11282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03096_ clkbuf_0__03096_/X vssd1 vssd1 vccd1 vccd1 _14168__446/A sky130_fd_sc_hd__clkbuf_16
X_13021_ _13010_/X _13011_/X _13020_/X _17686_/Q vssd1 vssd1 vccd1 vccd1 _13022_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ _10233_/A vssd1 vssd1 vccd1 vccd1 _18673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10164_ _10164_/A vssd1 vssd1 vccd1 vccd1 _18700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17760_ _19327_/CLK _17760_/D vssd1 vssd1 vccd1 vccd1 _17760_/Q sky130_fd_sc_hd__dfxtp_1
X_14972_ _15026_/A vssd1 vssd1 vccd1 vccd1 _15057_/A sky130_fd_sc_hd__clkbuf_2
X_10095_ _10110_/S vssd1 vssd1 vccd1 vccd1 _10104_/S sky130_fd_sc_hd__buf_2
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13923_ _13133_/B _13923_/B vssd1 vssd1 vccd1 vccd1 _13945_/B sky130_fd_sc_hd__and2b_1
X_16711_ _19108_/Q _16689_/X _13359_/X vssd1 vssd1 vccd1 vccd1 _19108_/D sky130_fd_sc_hd__o21ba_1
X_17085__68 _17086__69/A vssd1 vssd1 vccd1 vccd1 _19217_/CLK sky130_fd_sc_hd__inv_2
XFILLER_247_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17691_ _18007_/CLK _17691_/D vssd1 vssd1 vccd1 vccd1 _17691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _17928_/Q _13850_/X _13853_/Y _13841_/X vssd1 vssd1 vccd1 vccd1 _17928_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _17644_/Q _17991_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12806_/B sky130_fd_sc_hd__mux2_1
XFILLER_222_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16573_ _19018_/Q _16569_/B _16572_/Y vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__o21a_1
XFILLER_90_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13785_ _17905_/Q _13770_/X _13784_/Y vssd1 vssd1 vccd1 vccd1 _17905_/D sky130_fd_sc_hd__o21a_1
XFILLER_76_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ _10997_/A vssd1 vssd1 vccd1 vccd1 _18279_/D sky130_fd_sc_hd__clkbuf_1
X_15524_ _15524_/A _15524_/B _15524_/C _15524_/D vssd1 vssd1 vccd1 vccd1 _15525_/D
+ sky130_fd_sc_hd__nand4_1
X_18312_ _18312_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _12736_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _17628_/D sky130_fd_sc_hd__nor2_1
XFILLER_187_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19292_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18243_/CLK _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15455_ _15455_/A vssd1 vssd1 vccd1 vccd1 _15455_/X sky130_fd_sc_hd__buf_1
X_12667_ _12680_/C vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14406_ _14412_/A vssd1 vssd1 vccd1 vccd1 _14406_/X sky130_fd_sc_hd__buf_1
XFILLER_198_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11618_ _11618_/A vssd1 vssd1 vccd1 vccd1 _17565_/D sky130_fd_sc_hd__clkbuf_1
X_18174_ _18174_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15386_ _15410_/A vssd1 vssd1 vccd1 vccd1 _15386_/X sky130_fd_sc_hd__buf_1
X_12598_ _18013_/Q _17589_/Q _17590_/Q vssd1 vssd1 vccd1 vccd1 _12599_/C sky130_fd_sc_hd__a21o_1
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17125_ _17125_/A vssd1 vssd1 vccd1 vccd1 _19222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14337_ _14349_/A vssd1 vssd1 vccd1 vccd1 _14337_/X sky130_fd_sc_hd__buf_1
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11549_ _17711_/Q _10887_/X _11557_/S vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17056_ _17062_/A vssd1 vssd1 vccd1 vccd1 _17056_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__03794_ _15386_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03794_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163__870 _15165__872/A vssd1 vssd1 vccd1 vccd1 _18546_/CLK sky130_fd_sc_hd__inv_2
X_16007_ _18870_/Q _16007_/B vssd1 vssd1 vccd1 vccd1 _16018_/C sky130_fd_sc_hd__and2_1
X_13219_ _13232_/A vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _18071_/Q input51/X _14207_/S vssd1 vssd1 vccd1 vccd1 _14200_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _15244_/A _10219_/B vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17958_ _17959_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_81_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18655_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16909_ _16929_/A _16909_/B vssd1 vssd1 vccd1 vccd1 _16909_/Y sky130_fd_sc_hd__nor2_1
X_17889_ _18024_/CLK _17889_/D vssd1 vssd1 vccd1 vccd1 _17889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18572_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ _08929_/X _19103_/Q _09312_/S vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03159_ _14331_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03159_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09243_ _18564_/Q _09256_/B _10402_/A vssd1 vssd1 vccd1 vccd1 _09247_/C sky130_fd_sc_hd__a21oi_1
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706__1000 _15707__1001/A vssd1 vssd1 vccd1 vccd1 _18717_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _19169_/Q _09096_/X _09178_/S vssd1 vssd1 vccd1 vccd1 _09175_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16685__316 _16685__316/A vssd1 vssd1 vccd1 vccd1 _19090_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15437__931 _15439__933/A vssd1 vssd1 vccd1 vccd1 _18618_/CLK sky130_fd_sc_hd__inv_2
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08958_ _09688_/A vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__buf_4
XFILLER_248_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _08911_/B _08889_/B _08769_/B vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__or3b_4
XFILLER_99_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10920_ _10920_/A vssd1 vssd1 vccd1 vccd1 _18312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _10851_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _10867_/S sky130_fd_sc_hd__nor2_2
XFILLER_204_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ _13165_/X _13557_/B _13568_/Y _13569_/X vssd1 vssd1 vccd1 vccd1 _17835_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10782_ _10782_/A vssd1 vssd1 vccd1 vccd1 _18374_/D sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12459_/X _12453_/X _12464_/X _12458_/X _12474_/A _12407_/A vssd1 vssd1 vccd1
+ vccd1 _12521_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _08749_/X _14244_/A _17303_/A vssd1 vssd1 vccd1 vccd1 _16036_/B sky130_fd_sc_hd__a21oi_2
X_12452_ _12351_/X _12932_/A _13094_/B vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__o21ba_1
XFILLER_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11403_ _11418_/S vssd1 vssd1 vccd1 vccd1 _11412_/S sky130_fd_sc_hd__clkbuf_2
X_12383_ _17601_/Q vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14122_ _18024_/Q _14114_/X _14121_/Y vssd1 vssd1 vccd1 vccd1 _18024_/D sky130_fd_sc_hd__o21a_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11334_ _11334_/A vssd1 vssd1 vccd1 vccd1 _18143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03148_ clkbuf_0__03148_/X vssd1 vssd1 vccd1 vccd1 _14280__479/A sky130_fd_sc_hd__clkbuf_16
XFILLER_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14053_ _14053_/A _14053_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _14055_/A sky130_fd_sc_hd__and3_2
X_18930_ _18930_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_2
X_11265_ _18169_/Q _11264_/X _11274_/S vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13004_ _17672_/Q _13081_/B vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__xor2_1
XFILLER_140_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10216_ _10216_/A vssd1 vssd1 vccd1 vccd1 _18680_/D sky130_fd_sc_hd__clkbuf_1
X_18861_ _18876_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_1
X_11196_ _18198_/Q _11056_/X _11196_/S vssd1 vssd1 vccd1 vccd1 _11197_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17812_ _19339_/CLK _17812_/D vssd1 vssd1 vccd1 vccd1 _17812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _18707_/Q _10060_/X _10149_/S vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__mux2_1
X_18792_ _18792_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17058__46 _17058__46/A vssd1 vssd1 vccd1 vccd1 _19195_/CLK sky130_fd_sc_hd__inv_2
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ _14963_/C _14960_/C _14955_/C _14955_/D vssd1 vssd1 vccd1 vccd1 _14956_/C
+ sky130_fd_sc_hd__or4_1
X_17743_ _19336_/CLK _17743_/D vssd1 vssd1 vccd1 vccd1 _17743_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__05080_ clkbuf_0__05080_/X vssd1 vssd1 vccd1 vccd1 _17405__96/A sky130_fd_sc_hd__clkbuf_16
X_10078_ _18734_/Q _10048_/X _10086_/S vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__mux2_1
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _13256_/X _13903_/X _13894_/X vssd1 vssd1 vccd1 vccd1 _13906_/Y sky130_fd_sc_hd__a21oi_1
X_17674_ _19037_/CLK _17674_/D vssd1 vssd1 vccd1 vccd1 _17674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_202 _13192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_213 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ _17922_/Q _13829_/X _13836_/X _13826_/X vssd1 vssd1 vccd1 vccd1 _17922_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_224 _16715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081__195 _16081__195/A vssd1 vssd1 vccd1 vccd1 _18900_/CLK sky130_fd_sc_hd__inv_2
XFILLER_223_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16556_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16556_/X sky130_fd_sc_hd__buf_1
X_19344_ _19344_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
X_13768_ _17900_/Q _13762_/X _13767_/Y vssd1 vssd1 vccd1 vccd1 _17900_/D sky130_fd_sc_hd__o21a_1
XFILLER_149_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12719_ _12717_/A _12716_/A _12718_/X vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__o21ai_1
XFILLER_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15507_ _15505_/B _15505_/C _15572_/B vssd1 vssd1 vccd1 vccd1 _15525_/C sky130_fd_sc_hd__a21oi_1
X_19275_ _19340_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
X_16487_ _18980_/Q _16492_/C vssd1 vssd1 vccd1 vccd1 _16491_/B sky130_fd_sc_hd__and2_1
X_13699_ _17877_/Q _13683_/X _13698_/Y vssd1 vssd1 vccd1 vccd1 _17877_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18226_ _18226_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _19323_/Q _19307_/Q _19299_/Q _19274_/Q _15293_/X _15215_/X vssd1 vssd1 vccd1
+ vccd1 _15369_/X sky130_fd_sc_hd__mux4_2
X_18157_ _18157_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17108_ _17102_/Y _17103_/Y _17108_/C _17117_/A vssd1 vssd1 vccd1 vccd1 _17109_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_85_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18088_ _18482_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09930_ _18784_/Q _09277_/X _09932_/S vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09861_/A vssd1 vssd1 vccd1 vccd1 _15808_/B sky130_fd_sc_hd__buf_8
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _09508_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08828_/S sky130_fd_sc_hd__nor2_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _18835_/Q _09744_/X _09800_/S vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__mux2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08743_ _18069_/Q _08743_/B vssd1 vssd1 vccd1 vccd1 _13130_/B sky130_fd_sc_hd__or2_2
XFILLER_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09226_ _18562_/Q vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09157_ _09157_/A vssd1 vssd1 vccd1 vccd1 _19177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09088_ _09117_/S vssd1 vssd1 vccd1 vccd1 _09105_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17414__104 _17414__104/A vssd1 vssd1 vccd1 vccd1 _19317_/CLK sky130_fd_sc_hd__inv_2
X_11050_ _18666_/Q vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10001_ _10001_/A vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14740_ _14544_/A _14739_/X _14619_/A vssd1 vssd1 vccd1 vccd1 _14740_/Y sky130_fd_sc_hd__o21ai_1
X_11952_ _12005_/S vssd1 vssd1 vccd1 vccd1 _11977_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _10903_/A vssd1 vssd1 vccd1 vccd1 _18318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _18857_/Q _18351_/Q _19192_/Q _18359_/Q _14553_/X _14600_/X vssd1 vssd1 vccd1
+ vccd1 _14671_/X sky130_fd_sc_hd__mux4_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _12229_/A vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__buf_1
XFILLER_60_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _18968_/Q _17808_/Q _16410_/S vssd1 vssd1 vccd1 vccd1 _16410_/X sky130_fd_sc_hd__mux2_1
X_13622_ _13165_/X _13608_/B _13621_/Y _13619_/X vssd1 vssd1 vccd1 vccd1 _17852_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17390_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17390_/X sky130_fd_sc_hd__buf_1
X_10834_ _10849_/S vssd1 vssd1 vccd1 vccd1 _10843_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15114__831 _15114__831/A vssd1 vssd1 vccd1 vccd1 _18507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16341_ _16543_/A vssd1 vssd1 vccd1 vccd1 _16341_/X sky130_fd_sc_hd__buf_1
XFILLER_201_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _17829_/Q _13557_/B vssd1 vssd1 vccd1 vccd1 _13553_/Y sky130_fd_sc_hd__nor2_1
X_10765_ _10765_/A vssd1 vssd1 vccd1 vccd1 _18381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12504_ _12504_/A _12764_/A vssd1 vssd1 vccd1 vccd1 _12504_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19060_ _19060_/CLK _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16272_ _16291_/A _16272_/B vssd1 vssd1 vccd1 vccd1 _16272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _17808_/Q _16520_/A _13484_/S vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10696_ _18409_/Q _10695_/X _10705_/S vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _18012_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15223_ _15213_/X _15216_/X _15217_/X _15219_/X _15220_/X _15222_/X vssd1 vssd1 vccd1
+ vccd1 _15223_/X sky130_fd_sc_hd__mux4_1
X_12435_ _12435_/A vssd1 vssd1 vccd1 vccd1 _12436_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03600_ clkbuf_0__03600_/X vssd1 vssd1 vccd1 vccd1 _15161__869/A sky130_fd_sc_hd__clkbuf_16
X_12366_ _12432_/S vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_165_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14105_ _18018_/Q _14091_/X _14104_/Y vssd1 vssd1 vccd1 vccd1 _18018_/D sky130_fd_sc_hd__o21a_1
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11317_ _11162_/X _18148_/Q _11319_/S vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__mux2_1
X_12297_ _17549_/Q _12187_/X _12185_/X _17563_/Q vssd1 vssd1 vccd1 vccd1 _12301_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14036_ _17992_/Q _14032_/X _14035_/Y vssd1 vssd1 vccd1 vccd1 _17992_/D sky130_fd_sc_hd__o21a_1
X_18913_ _18913_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11248_ _11248_/A vssd1 vssd1 vccd1 vccd1 _18176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18844_ _18844_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_1
X_11179_ _11179_/A vssd1 vssd1 vccd1 vccd1 _18206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18775_ _18775_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _18866_/Q _15993_/B vssd1 vssd1 vccd1 vccd1 _15987_/Y sky130_fd_sc_hd__nand2_1
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17726_ _17878_/CLK _17726_/D vssd1 vssd1 vccd1 vccd1 _17726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14938_ _14938_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _14939_/B sky130_fd_sc_hd__nand2_1
XFILLER_224_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04014_ clkbuf_0__04014_/X vssd1 vssd1 vccd1 vccd1 _15879__174/A sky130_fd_sc_hd__clkbuf_16
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17657_ _17969_/CLK _17657_/D vssd1 vssd1 vccd1 vccd1 _17657_/Q sky130_fd_sc_hd__dfxtp_1
X_14165__444 _14165__444/A vssd1 vssd1 vccd1 vccd1 _18052_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16608_ _16620_/A _16608_/B vssd1 vssd1 vccd1 vccd1 _16608_/Y sky130_fd_sc_hd__nor2_1
X_17588_ _17588_/CLK _17588_/D vssd1 vssd1 vccd1 vccd1 _17588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19327_ _19327_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_32_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19258_ _19261_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09011_ _09011_/A _09010_/X vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__or2b_1
XFILLER_192_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18209_ _18209_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19189_ _19189_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__04847_ clkbuf_0__04847_/X vssd1 vssd1 vccd1 vccd1 _17061__49/A sky130_fd_sc_hd__clkbuf_16
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16723__338 _16723__338/A vssd1 vssd1 vccd1 vccd1 _19117_/CLK sky130_fd_sc_hd__inv_2
X_09913_ _18791_/Q _09741_/X _09913_/S vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09844_ _18811_/Q vssd1 vssd1 vccd1 vccd1 _16892_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09775_ _08868_/X _18842_/Q _09781_/S vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08726_ _18089_/Q vssd1 vssd1 vccd1 vccd1 _11779_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03620_ clkbuf_0__03620_/X vssd1 vssd1 vccd1 vccd1 _15203__888/A sky130_fd_sc_hd__clkbuf_16
XFILLER_227_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10550_ _18506_/Q _10117_/A _10556_/S vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _19154_/Q _09092_/X _09215_/S vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10481_ _10481_/A vssd1 vssd1 vccd1 vccd1 _18537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__05083_ clkbuf_0__05083_/X vssd1 vssd1 vccd1 vccd1 _17502__9/A sky130_fd_sc_hd__clkbuf_16
XFILLER_182_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ _12179_/Y _12218_/X _12136_/S _16619_/A vssd1 vssd1 vccd1 vccd1 _17531_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _12149_/X _12151_/B vssd1 vssd1 vccd1 vccd1 _12152_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11102_ _09051_/X _18236_/Q _11104_/S vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12082_ _12082_/A vssd1 vssd1 vccd1 vccd1 _12082_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15910_ _15937_/B _15909_/C _18868_/Q vssd1 vssd1 vccd1 vccd1 _15936_/B sky130_fd_sc_hd__a21oi_1
X_11033_ _11033_/A vssd1 vssd1 vccd1 vccd1 _18263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16890_ _09845_/X _16875_/X _16889_/Y vssd1 vssd1 vccd1 vccd1 _16890_/X sky130_fd_sc_hd__a21o_1
XFILLER_209_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18560_ _18560_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _12975_/X _12984_/B vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__and2b_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17511_ _17511_/CLK _17511_/D vssd1 vssd1 vccd1 vccd1 _17511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11935_ _19226_/Q _17142_/A _12025_/S vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__mux2_1
X_14723_ _18329_/Q _14543_/A _14623_/X _14722_/X vssd1 vssd1 vccd1 vccd1 _18329_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18491_ _18491_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14342__529 _14342__529/A vssd1 vssd1 vccd1 vccd1 _18164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _17747_/Q _19329_/Q _17451_/S vssd1 vssd1 vccd1 vccd1 _17443_/B sky130_fd_sc_hd__mux2_1
X_14654_ _18588_/Q _18302_/Q _17568_/Q _18839_/Q _14575_/X _09459_/X vssd1 vssd1 vccd1
+ vccd1 _14654_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ _11866_/A vssd1 vssd1 vccd1 vccd1 _11866_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _13434_/X _13601_/X _13603_/Y _13604_/X vssd1 vssd1 vccd1 vccd1 _17845_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_232_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10817_ _18362_/Q _10789_/X _10825_/S vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17373_ _19285_/Q _17491_/B vssd1 vssd1 vccd1 vccd1 _17377_/A sky130_fd_sc_hd__xnor2_1
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14585_ _14544_/A _14584_/X _14619_/A vssd1 vssd1 vccd1 vccd1 _14585_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ input9/X _11790_/Y _11793_/X _17916_/Q _11796_/X vssd1 vssd1 vccd1 vccd1
+ _11797_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19112_ _19112_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13536_ _17823_/Q _13522_/X _13535_/Y vssd1 vssd1 vccd1 vccd1 _17823_/D sky130_fd_sc_hd__o21a_1
X_10748_ _18388_/Q _10710_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10749_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16255_ _18919_/Q _16164_/X _16254_/Y _16216_/X vssd1 vssd1 vccd1 vccd1 _18919_/D
+ sky130_fd_sc_hd__o211a_1
X_19043_ _19043_/CLK _19043_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_13467_ _17803_/Q _16530_/A _13477_/B vssd1 vssd1 vccd1 vccd1 _13468_/B sky130_fd_sc_hd__mux2_1
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10679_ _10679_/A vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__clkbuf_1
X_15206_ _16294_/C _15955_/A vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__and2_1
X_12418_ _12415_/X _12416_/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12418_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16186_ _16180_/X _16184_/X _16271_/S vssd1 vssd1 vccd1 vccd1 _16187_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13398_ _14069_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13414_/B sky130_fd_sc_hd__or2_1
XFILLER_126_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15137_ _15149_/A vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__buf_1
XFILLER_245_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12349_ _18004_/Q vssd1 vssd1 vccd1 vccd1 _14065_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15068_ _16056_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _18475_/D sky130_fd_sc_hd__nor2_1
XFILLER_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14019_ _17986_/Q _14011_/X _14018_/Y vssd1 vssd1 vccd1 vccd1 _17986_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18827_ _18827_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09560_ _08941_/X _18951_/Q _09560_/S vssd1 vssd1 vccd1 vccd1 _09561_/A sky130_fd_sc_hd__mux2_1
X_18758_ _18758_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17709_ _17709_/CLK _17709_/D vssd1 vssd1 vccd1 vccd1 _17709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09491_ _09491_/A vssd1 vssd1 vccd1 vccd1 _19010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18689_ _18689_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__05077_ _17390_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05077_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_247_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _09842_/S vssd1 vssd1 vccd1 vccd1 _09836_/S sky130_fd_sc_hd__buf_2
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ _18883_/Q vssd1 vssd1 vccd1 vccd1 _09758_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09689_ _09688_/X _18901_/Q _09689_/S vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__mux2_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11720_ _17784_/Q _17785_/Q vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__and2b_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ _08801_/X _17533_/Q _11653_/S vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10602_ _10638_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10618_/S sky130_fd_sc_hd__or2_2
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11582_ _11582_/A vssd1 vssd1 vccd1 vccd1 _17581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13321_ _13271_/X _13311_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03396_ clkbuf_0__03396_/X vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__clkbuf_16
X_10533_ _10533_/A vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16040_ _18888_/Q _16049_/C vssd1 vssd1 vccd1 vccd1 _16040_/Y sky130_fd_sc_hd__nor2_1
X_13252_ _13259_/A vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10464_ _18544_/Q _10339_/X _10466_/S vssd1 vssd1 vccd1 vccd1 _10465_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12203_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__buf_2
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13183_ _13404_/A vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__buf_6
X_10395_ _16194_/A vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_237_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12134_ _12132_/X _12134_/B vssd1 vssd1 vccd1 vccd1 _12135_/A sky130_fd_sc_hd__and2b_1
XFILLER_150_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _17991_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12065_ _19220_/Q vssd1 vssd1 vccd1 vccd1 _17117_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_123_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16942_ _16938_/X _16941_/X _16980_/S vssd1 vssd1 vccd1 vccd1 _16942_/X sky130_fd_sc_hd__mux2_2
XFILLER_111_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _09043_/X _18270_/Q _11016_/S vssd1 vssd1 vccd1 vccd1 _11017_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16873_ _16900_/A vssd1 vssd1 vccd1 vccd1 _16976_/S sky130_fd_sc_hd__buf_2
XFILLER_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18612_ _18612_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03161_ clkbuf_0__03161_/X vssd1 vssd1 vccd1 vccd1 _14347__533/A sky130_fd_sc_hd__clkbuf_16
X_15824_ _15824_/A vssd1 vssd1 vccd1 vccd1 _15824_/X sky130_fd_sc_hd__buf_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03192_ _14499_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03192_/X sky130_fd_sc_hd__clkbuf_16
X_18543_ _18543_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_1
X_12967_ _12967_/A vssd1 vssd1 vccd1 vccd1 _17675_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03092_ clkbuf_0__03092_/X vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__clkbuf_16
X_15755_ _15779_/A vssd1 vssd1 vccd1 vccd1 _15755_/X sky130_fd_sc_hd__buf_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _11912_/X _11917_/X _12076_/S vssd1 vssd1 vccd1 vccd1 _11918_/X sky130_fd_sc_hd__mux2_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _18409_/Q _18401_/Q _19314_/Q _17718_/Q _14641_/A _14546_/X vssd1 vssd1 vccd1
+ vccd1 _14706_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18474_ _18477_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
X_12898_ _12898_/A vssd1 vssd1 vccd1 vccd1 _17662_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15686_ _15686_/A vssd1 vssd1 vccd1 vccd1 _15686_/X sky130_fd_sc_hd__buf_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17752_/Q _19324_/Q _17497_/B vssd1 vssd1 vccd1 vccd1 _17426_/B sky130_fd_sc_hd__mux2_1
XFILLER_178_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ _11849_/A vssd1 vssd1 vccd1 vccd1 _11849_/X sky130_fd_sc_hd__clkbuf_1
X_14637_ _14637_/A vssd1 vssd1 vccd1 vccd1 _14637_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17356_ _17437_/A vssd1 vssd1 vccd1 vccd1 _17356_/X sky130_fd_sc_hd__clkbuf_2
X_14568_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14568_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_158_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _17772_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13519_ _17818_/Q _13500_/X _13518_/Y vssd1 vssd1 vccd1 vccd1 _17818_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17287_ _17288_/B _17279_/A _17288_/D _19265_/Q vssd1 vssd1 vccd1 vccd1 _17289_/B
+ sky130_fd_sc_hd__a31o_1
X_14499_ _14505_/A vssd1 vssd1 vccd1 vccd1 _14499_/X sky130_fd_sc_hd__buf_1
XFILLER_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19026_ _19027_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16238_ _16257_/A _16238_/B vssd1 vssd1 vccd1 vccd1 _16238_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127__841 _15128__842/A vssd1 vssd1 vccd1 vccd1 _18517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_126_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _16257_/A _16169_/B vssd1 vssd1 vccd1 vccd1 _16169_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08991_ _11321_/A vssd1 vssd1 vccd1 vccd1 _08991_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04577_ _16676_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04577_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09612_ _09612_/A _09612_/B _09612_/C _08761_/X vssd1 vssd1 vccd1 vccd1 _16294_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_205_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431__926 _15433__928/A vssd1 vssd1 vccd1 vccd1 _18613_/CLK sky130_fd_sc_hd__inv_2
XFILLER_209_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09543_ _09543_/A vssd1 vssd1 vccd1 vccd1 _18959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09474_ _09474_/A vssd1 vssd1 vccd1 vccd1 _19044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03181_ clkbuf_0__03181_/X vssd1 vssd1 vccd1 vccd1 _14448__614/A sky130_fd_sc_hd__clkbuf_16
XFILLER_137_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ _18479_/Q vssd1 vssd1 vccd1 vccd1 _10180_/X sky130_fd_sc_hd__buf_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13870_ input55/X vssd1 vssd1 vccd1 vccd1 _13871_/A sky130_fd_sc_hd__inv_2
XFILLER_235_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ _12821_/A vssd1 vssd1 vccd1 vccd1 _17648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12752_ _12758_/C _12758_/D _12751_/Y vssd1 vssd1 vccd1 vccd1 _17633_/D sky130_fd_sc_hd__a21oi_1
XFILLER_199_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15540_ _18643_/Q _15543_/C vssd1 vssd1 vccd1 vccd1 _15540_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11703_ _17906_/Q _17721_/Q _11707_/S vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__mux2_8
XFILLER_70_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15471_ _18641_/Q _15624_/A _15616_/A vssd1 vssd1 vccd1 vccd1 _18641_/D sky130_fd_sc_hd__a21o_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12687_/A _12683_/B vssd1 vssd1 vccd1 vccd1 _17612_/D sky130_fd_sc_hd__nor2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17210_/A _17216_/D vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__and2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11634_ _11634_/A vssd1 vssd1 vccd1 vccd1 _17541_/D sky130_fd_sc_hd__clkbuf_1
X_18190_ _18190_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17141_ _17141_/A vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11565_ _11565_/A hold13/A vssd1 vssd1 vccd1 vccd1 _11581_/S sky130_fd_sc_hd__nor2_2
XFILLER_128_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13304_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13304_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10516_ _18521_/Q _10336_/X _10520_/S vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11496_ _11496_/A vssd1 vssd1 vccd1 vccd1 _18047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13235_ _13146_/X _13232_/X _13224_/X vssd1 vssd1 vccd1 vccd1 _13235_/Y sky130_fd_sc_hd__a21oi_1
X_16023_ _18873_/Q _16027_/C vssd1 vssd1 vccd1 vccd1 _16024_/C sky130_fd_sc_hd__and2_1
X_10447_ _10447_/A vssd1 vssd1 vccd1 vccd1 _18552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13166_ _17728_/Q _14134_/B vssd1 vssd1 vccd1 vccd1 _13166_/Y sky130_fd_sc_hd__nor2_1
XFILLER_237_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10378_ _08789_/X _18582_/Q _10382_/S vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__mux2_1
X_12117_ _17778_/Q _12057_/X _11944_/A vssd1 vssd1 vccd1 vccd1 _12117_/X sky130_fd_sc_hd__o21a_1
X_17974_ _18001_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_1
X_13097_ _13097_/A _13097_/B _13097_/C _13097_/D vssd1 vssd1 vccd1 vccd1 _13097_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _17777_/Q vssd1 vssd1 vccd1 vccd1 _12069_/A sky130_fd_sc_hd__clkbuf_2
X_16925_ _16963_/A _16925_/B vssd1 vssd1 vccd1 vccd1 _16925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16856_ _16929_/A _16856_/B vssd1 vssd1 vccd1 vccd1 _16856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_226_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03144_ clkbuf_0__03144_/X vssd1 vssd1 vccd1 vccd1 _14261__464/A sky130_fd_sc_hd__clkbuf_16
XFILLER_20_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16787_ _19136_/Q _19134_/Q _16787_/S vssd1 vssd1 vccd1 vccd1 _16788_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13999_ _17979_/Q _13988_/X _13998_/Y vssd1 vssd1 vccd1 vccd1 _17979_/D sky130_fd_sc_hd__o21a_1
XFILLER_209_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18526_ _18526_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03175_ _14412_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03175_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_248_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18457_ _19039_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15684__983 _15685__984/A vssd1 vssd1 vccd1 vccd1 _18700_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _19162_/Q _09127_/X _09196_/S vssd1 vssd1 vccd1 vccd1 _09191_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18388_ _18388_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _17339_/A vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03977_ clkbuf_0__03977_/X vssd1 vssd1 vccd1 vccd1 _15727__1017/A sky130_fd_sc_hd__clkbuf_16
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19009_ _19009_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04529_ clkbuf_0__04529_/X vssd1 vssd1 vccd1 vccd1 _16552__261/A sky130_fd_sc_hd__clkbuf_16
X_08974_ _19219_/Q _08944_/X _08982_/S vssd1 vssd1 vccd1 vccd1 _08975_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09526_ _10967_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _09542_/S sky130_fd_sc_hd__nor2_2
XFILLER_231_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _19046_/Q vssd1 vssd1 vccd1 vccd1 _14594_/A sky130_fd_sc_hd__buf_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ _19070_/Q _08958_/X _09388_/S vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11350_ _11350_/A vssd1 vssd1 vccd1 vccd1 _18138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03164_ clkbuf_0__03164_/X vssd1 vssd1 vccd1 vccd1 _14361__544/A sky130_fd_sc_hd__clkbuf_16
X_10301_ _10301_/A vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__clkbuf_1
X_11281_ _11281_/A vssd1 vssd1 vccd1 vccd1 _18164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _13020_/A _13020_/B _13020_/C _13020_/D vssd1 vssd1 vccd1 vccd1 _13020_/X
+ sky130_fd_sc_hd__and4_1
Xclkbuf_1_0__f__03095_ clkbuf_0__03095_/X vssd1 vssd1 vccd1 vccd1 _14165__444/A sky130_fd_sc_hd__clkbuf_16
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10232_ _18673_/Q _09761_/X hold3/X vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14152__435 _14155__438/A vssd1 vssd1 vccd1 vccd1 _18043_/CLK sky130_fd_sc_hd__inv_2
X_10163_ _18700_/Q _10057_/X _10167_/S vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _14971_/A vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__clkbuf_1
X_10094_ _10094_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10110_/S sky130_fd_sc_hd__nor2_2
XFILLER_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13922_ _17951_/Q _13903_/X _13921_/Y vssd1 vssd1 vccd1 vccd1 _17951_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17690_ _17959_/CLK _17690_/D vssd1 vssd1 vccd1 vccd1 _17690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13853_ _13853_/A _13863_/B vssd1 vssd1 vccd1 vccd1 _13853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14460__623 _14460__623/A vssd1 vssd1 vccd1 vccd1 _18258_/CLK sky130_fd_sc_hd__inv_2
X_12804_ _12804_/A vssd1 vssd1 vccd1 vccd1 _17643_/D sky130_fd_sc_hd__clkbuf_1
X_16572_ _16602_/A _16576_/C vssd1 vssd1 vccd1 vccd1 _16572_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13784_ _13783_/X _13778_/X _13774_/X vssd1 vssd1 vccd1 vccd1 _13784_/Y sky130_fd_sc_hd__a21oi_1
X_10996_ _18279_/Q _09133_/X _10998_/S vssd1 vssd1 vccd1 vccd1 _10997_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18311_ _18311_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15523_ _15523_/A _15523_/B _15523_/C _15523_/D vssd1 vssd1 vccd1 vccd1 _15524_/D
+ sky130_fd_sc_hd__nor4_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12737_/B _12732_/A _12734_/X vssd1 vssd1 vccd1 vccd1 _12736_/B sky130_fd_sc_hd__o21ai_1
X_19291_ _19340_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18242_ _18242_/CLK _18242_/D vssd1 vssd1 vccd1 vccd1 _18242_/Q sky130_fd_sc_hd__dfxtp_1
X_12666_ _17608_/Q _17607_/Q _12666_/C _12666_/D vssd1 vssd1 vccd1 vccd1 _12680_/C
+ sky130_fd_sc_hd__and4_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11617_ _17565_/Q _10713_/A _11617_/S vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__mux2_1
X_18173_ _18173_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
X_12597_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__clkbuf_4
X_15385_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15385_/X sky130_fd_sc_hd__buf_1
XFILLER_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17124_ _17129_/C _17124_/B _17277_/B vssd1 vssd1 vccd1 vccd1 _17125_/A sky130_fd_sc_hd__and3b_1
XFILLER_156_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11548_ _11563_/S vssd1 vssd1 vccd1 vccd1 _11557_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_237_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03793_ _15385_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03793_/X sky130_fd_sc_hd__clkbuf_16
X_11479_ _09127_/X _18054_/Q _11485_/S vssd1 vssd1 vccd1 vccd1 _11480_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _13232_/A vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__clkbuf_2
X_16006_ _18870_/Q _16007_/B vssd1 vssd1 vccd1 vccd1 _16008_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ _14231_/A vssd1 vssd1 vccd1 vccd1 _14207_/S sky130_fd_sc_hd__buf_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13149_ input57/X _13210_/B vssd1 vssd1 vccd1 vccd1 _13783_/A sky130_fd_sc_hd__nand2_4
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16643__283 _16643__283/A vssd1 vssd1 vccd1 vccd1 _19057_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _17963_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16908_ _18182_/Q _18174_/Q _18166_/Q _18158_/Q _16881_/X _16882_/X vssd1 vssd1 vccd1
+ vccd1 _16909_/B sky130_fd_sc_hd__mux4_1
X_17888_ _18024_/CLK _17888_/D vssd1 vssd1 vccd1 vccd1 _17888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16839_ _16818_/X _16838_/X _16797_/A vssd1 vssd1 vccd1 vccd1 _16839_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17991_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09311_ _09311_/A vssd1 vssd1 vccd1 vccd1 _19104_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03158_ _14325_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03158_/X sky130_fd_sc_hd__clkbuf_16
X_18509_ _18509_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14773__711 _14773__711/A vssd1 vssd1 vccd1 vccd1 _18354_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ _18565_/Q _09972_/A vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__xor2_2
Xclkbuf_0__03089_ _14139_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03089_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09173_ _09173_/A vssd1 vssd1 vccd1 vccd1 _19170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _08957_/A vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _08888_/A vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _10850_/A vssd1 vssd1 vccd1 vccd1 _18347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09524_/S vssd1 vssd1 vccd1 vccd1 _09518_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10781_ _18374_/Q _10704_/X _10781_/S vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__mux2_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12466_/X _12463_/X _12519_/X _12465_/X _12474_/A _12407_/A vssd1 vssd1 vccd1
+ vccd1 _12520_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A vssd1 vssd1 vccd1 vccd1 _13094_/B sky130_fd_sc_hd__buf_4
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _11475_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11418_/S sky130_fd_sc_hd__or2_2
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ _17600_/Q vssd1 vssd1 vccd1 vccd1 _12638_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14121_ _13746_/A _14120_/X _14108_/X vssd1 vssd1 vccd1 vccd1 _14121_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ _11332_/X _18143_/Q _11336_/S vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03147_ clkbuf_0__03147_/X vssd1 vssd1 vccd1 vccd1 _14271__471/A sky130_fd_sc_hd__clkbuf_16
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _17999_/Q _14033_/X _14051_/Y vssd1 vssd1 vccd1 vccd1 _17999_/D sky130_fd_sc_hd__o21a_1
XFILLER_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11264_ _18667_/Q vssd1 vssd1 vccd1 vccd1 _11264_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _17678_/Q _12920_/X _12921_/X _17677_/Q vssd1 vssd1 vccd1 vccd1 _13010_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10215_ _18680_/Q _09764_/X hold6/X vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_18860_ _18860_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_1
X_11195_ _11195_/A vssd1 vssd1 vccd1 vccd1 _18199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17811_ _19339_/CLK _17811_/D vssd1 vssd1 vccd1 vccd1 _17811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10146_ _10146_/A vssd1 vssd1 vccd1 vccd1 _18708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _18791_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _19336_/CLK _17742_/D vssd1 vssd1 vccd1 vccd1 _17742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14954_ _14962_/A _14964_/B _14954_/C vssd1 vssd1 vccd1 vccd1 _14955_/D sky130_fd_sc_hd__or3_1
X_10077_ _10092_/S vssd1 vssd1 vccd1 vccd1 _10086_/S sky130_fd_sc_hd__buf_2
XFILLER_43_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13905_ _17944_/Q _13902_/X _13904_/Y vssd1 vssd1 vccd1 vccd1 _17944_/D sky130_fd_sc_hd__o21a_1
X_17673_ _19037_/CLK _17673_/D vssd1 vssd1 vccd1 vccd1 _17673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_203 _16518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ input59/X _13845_/B vssd1 vssd1 vccd1 vccd1 _13836_/X sky130_fd_sc_hd__and2_1
XINSDIODE2_214 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_225 _16518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19343_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
X_13767_ _13712_/A _13762_/A _13701_/X vssd1 vssd1 vccd1 vccd1 _13767_/Y sky130_fd_sc_hd__a21oi_1
X_10979_ _18285_/Q _09761_/X hold11/X vssd1 vssd1 vccd1 vccd1 _10980_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ _18648_/Q vssd1 vssd1 vccd1 vccd1 _15572_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14837__763 _14838__764/A vssd1 vssd1 vccd1 vccd1 _18406_/CLK sky130_fd_sc_hd__inv_2
X_12718_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19274_ _19274_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ _18980_/Q _16492_/C vssd1 vssd1 vccd1 vccd1 _16488_/B sky130_fd_sc_hd__nor2_1
XFILLER_231_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13698_ _13271_/X _13688_/X _13689_/X vssd1 vssd1 vccd1 vccd1 _13698_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_176_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18225_ _18225_/CLK _18225_/D vssd1 vssd1 vccd1 vccd1 _18225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12649_ _12647_/X _12759_/A _12649_/C vssd1 vssd1 vccd1 vccd1 _12650_/A sky130_fd_sc_hd__and3b_1
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18156_ _18156_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15368_ _19119_/Q _18950_/Q _18608_/Q _19348_/Q _15251_/X _15291_/X vssd1 vssd1 vccd1
+ vccd1 _15368_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17107_ _13361_/X _17101_/A _13346_/B _17104_/X _17106_/Y vssd1 vssd1 vccd1 vccd1
+ _17108_/C sky130_fd_sc_hd__o41a_1
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18087_ _19339_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15299_ _15301_/A vssd1 vssd1 vccd1 vccd1 _15299_/X sky130_fd_sc_hd__buf_2
XFILLER_171_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09860_ _16875_/S _09872_/A vssd1 vssd1 vccd1 vccd1 _09860_/X sky130_fd_sc_hd__and2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _09377_/A _10219_/B _09789_/A vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__or3b_4
X_14467__629 _14467__629/A vssd1 vssd1 vccd1 vccd1 _18264_/CLK sky130_fd_sc_hd__inv_2
X_09791_ _09806_/S vssd1 vssd1 vccd1 vccd1 _09800_/S sky130_fd_sc_hd__buf_2
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18989_ _18993_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08742_ _18070_/Q _18071_/Q _18072_/Q _18073_/Q vssd1 vssd1 vccd1 vccd1 _08743_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16355__246 _16355__246/A vssd1 vssd1 vccd1 vccd1 _18962_/CLK sky130_fd_sc_hd__inv_2
XFILLER_224_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09225_ _18561_/Q vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _19177_/Q _09096_/X _09160_/S vssd1 vssd1 vccd1 vccd1 _09157_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _10833_/B _10752_/A vssd1 vssd1 vccd1 vccd1 _09117_/S sky130_fd_sc_hd__nor2_2
XFILLER_206_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15697__993 _15698__994/A vssd1 vssd1 vccd1 vccd1 _18710_/CLK sky130_fd_sc_hd__inv_2
XFILLER_190_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14292__489 _14292__489/A vssd1 vssd1 vccd1 vccd1 _18124_/CLK sky130_fd_sc_hd__inv_2
XFILLER_174_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10000_ _18764_/Q _09947_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _10001_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09989_ _09989_/A vssd1 vssd1 vccd1 vccd1 _18769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _17780_/Q vssd1 vssd1 vccd1 vccd1 _12005_/S sky130_fd_sc_hd__buf_2
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450__940 _15453__943/A vssd1 vssd1 vccd1 vccd1 _18627_/CLK sky130_fd_sc_hd__inv_2
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10902_ _18318_/Q _10901_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10903_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17063__50 _17067__54/A vssd1 vssd1 vccd1 vccd1 _19199_/CLK sky130_fd_sc_hd__inv_2
X_14670_ _18367_/Q _18319_/Q _18375_/Q _17708_/Q _14637_/A _14627_/X vssd1 vssd1 vccd1
+ vccd1 _14670_/X sky130_fd_sc_hd__mux4_1
X_11882_ _17421_/A vssd1 vssd1 vccd1 vccd1 _11882_/X sky130_fd_sc_hd__buf_1
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13621_ _17852_/Q _13621_/B vssd1 vssd1 vccd1 vccd1 _13621_/Y sky130_fd_sc_hd__nor2_1
X_10833_ _10851_/A _10833_/B vssd1 vssd1 vccd1 vccd1 _10849_/S sky130_fd_sc_hd__nor2_2
XFILLER_232_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16340_/X sky130_fd_sc_hd__buf_1
X_13552_ _13434_/X _13549_/X _13551_/Y _13472_/X vssd1 vssd1 vccd1 vccd1 _17828_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10764_ _18381_/Q _10707_/X _10768_/S vssd1 vssd1 vccd1 vccd1 _10765_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12503_ _12441_/X _12429_/X _12765_/S vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16271_ _16267_/X _16270_/X _16271_/S vssd1 vssd1 vccd1 vccd1 _16272_/B sky130_fd_sc_hd__mux2_1
X_13483_ input65/X _13483_/B vssd1 vssd1 vccd1 vccd1 _16520_/A sky130_fd_sc_hd__and2_4
XFILLER_41_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10695_ _10695_/A vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__buf_2
XFILLER_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18010_ _18010_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12434_ _12429_/X _12433_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12533_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15222_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15222_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12365_ _18012_/Q vssd1 vssd1 vccd1 vccd1 _12432_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16709__331 _16710__332/A vssd1 vssd1 vccd1 vccd1 _19106_/CLK sky130_fd_sc_hd__inv_2
XFILLER_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14104_ _13783_/A _14099_/X _14096_/X vssd1 vssd1 vccd1 vccd1 _14104_/Y sky130_fd_sc_hd__a21oi_1
X_11316_ _11316_/A vssd1 vssd1 vccd1 vccd1 _18149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12296_ _17551_/Q _12182_/X _12180_/X _17548_/Q vssd1 vssd1 vccd1 vccd1 _12301_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14035_ _13740_/A _14033_/X _14034_/X vssd1 vssd1 vccd1 vccd1 _14035_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18912_ _18912_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _11150_/X _18176_/Q _11251_/S vssd1 vssd1 vccd1 vccd1 _11248_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18843_ _18843_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11178_ _11156_/X _18206_/Q _11178_/S vssd1 vssd1 vccd1 vccd1 _11179_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10129_ _10129_/A vssd1 vssd1 vccd1 vccd1 _10129_/X sky130_fd_sc_hd__clkbuf_4
X_18774_ _18774_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15986_ _15986_/A _15986_/B _15991_/B vssd1 vssd1 vccd1 vccd1 _15986_/X sky130_fd_sc_hd__or3_1
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17725_ _18031_/CLK _17725_/D vssd1 vssd1 vccd1 vccd1 _17725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14937_ _17853_/Q _14930_/A _17852_/Q vssd1 vssd1 vccd1 vccd1 _14938_/B sky130_fd_sc_hd__o21ai_1
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04013_ clkbuf_0__04013_/X vssd1 vssd1 vccd1 vccd1 _15873__169/A sky130_fd_sc_hd__clkbuf_16
XFILLER_223_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17656_ _18006_/CLK _17656_/D vssd1 vssd1 vccd1 vccd1 _17656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16607_ _16613_/A _16607_/B _16607_/C vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__nor3_1
X_13819_ _13849_/B vssd1 vssd1 vccd1 vccd1 _13828_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17587_ _17587_/CLK _17587_/D vssd1 vssd1 vccd1 vccd1 _17587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19326_ _19327_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16538_ _16506_/A _16534_/X _16429_/Y _14589_/X vssd1 vssd1 vccd1 vccd1 _18996_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19257_ _19261_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16469_ _16469_/A vssd1 vssd1 vccd1 vccd1 _16469_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09010_ _18810_/Q hold25/A vssd1 vssd1 vccd1 vccd1 _09010_/X sky130_fd_sc_hd__xor2_1
X_18208_ _18208_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__04846_ clkbuf_0__04846_/X vssd1 vssd1 vccd1 vccd1 _17053__42/A sky130_fd_sc_hd__clkbuf_16
X_19188_ _19188_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _18139_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
X_14885__801 _14886__802/A vssd1 vssd1 vccd1 vccd1 _18446_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09912_ _09912_/A vssd1 vssd1 vccd1 vccd1 _18792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09843_ _09843_/A vssd1 vssd1 vccd1 vccd1 _18812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09774_ _09774_/A vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08725_ _18090_/Q vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16656__293 _16657__294/A vssd1 vssd1 vccd1 vccd1 _19067_/CLK sky130_fd_sc_hd__inv_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09208_ _09208_/A vssd1 vssd1 vccd1 vccd1 _19155_/D sky130_fd_sc_hd__clkbuf_1
X_10480_ _18537_/Q _10336_/X _10484_/S vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__05082_ clkbuf_0__05082_/X vssd1 vssd1 vccd1 vccd1 _17419__108/A sky130_fd_sc_hd__clkbuf_16
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09139_ _18663_/Q vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__buf_2
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12150_ _17522_/Q _17729_/Q _12153_/S vssd1 vssd1 vccd1 vccd1 _12151_/B sky130_fd_sc_hd__mux2_1
X_14786__721 _14786__721/A vssd1 vssd1 vccd1 vccd1 _18364_/CLK sky130_fd_sc_hd__inv_2
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17501__8 _17501__8/A vssd1 vssd1 vccd1 vccd1 _19343_/CLK sky130_fd_sc_hd__inv_2
X_11101_ _11101_/A vssd1 vssd1 vccd1 vccd1 _18237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _11974_/X _11977_/X _12087_/S vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11032_ _18263_/Q _09133_/X _11034_/S vssd1 vssd1 vccd1 vccd1 _11033_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _17957_/Q _17680_/Q _12993_/S vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__mux2_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _17510_/CLK _17510_/D vssd1 vssd1 vccd1 vccd1 _17510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _14544_/X _14711_/X _14721_/Y vssd1 vssd1 vccd1 vccd1 _14722_/X sky130_fd_sc_hd__a21o_1
X_11934_ _19227_/Q vssd1 vssd1 vccd1 vccd1 _17142_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _18490_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17441_/A vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _14679_/A _14653_/B vssd1 vssd1 vccd1 vccd1 _14653_/Y sky130_fd_sc_hd__nor2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _13820_/A _11865_/B _11865_/C vssd1 vssd1 vccd1 vccd1 _11866_/A sky130_fd_sc_hd__and3_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13636_/A vssd1 vssd1 vccd1 vccd1 _13604_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17372_ _19276_/Q _12187_/A _12185_/X _19290_/Q vssd1 vssd1 vccd1 vccd1 _17378_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_10816_ _10831_/S vssd1 vssd1 vccd1 vccd1 _10825_/S sky130_fd_sc_hd__buf_2
XFILLER_158_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11796_ _11802_/A vssd1 vssd1 vccd1 vccd1 _11796_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14584_ _14561_/X _14566_/Y _14571_/Y _14577_/Y _14583_/Y vssd1 vssd1 vccd1 vccd1
+ _14584_/X sky130_fd_sc_hd__o32a_1
XFILLER_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19111_ _19128_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13535_ _13411_/X _13523_/A _13532_/X vssd1 vssd1 vccd1 vccd1 _13535_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ _10747_/A vssd1 vssd1 vccd1 vccd1 _18389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19042_ _19042_/CLK _19042_/D vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
X_16254_ _16190_/X _16245_/X _16253_/Y _16214_/X vssd1 vssd1 vccd1 vccd1 _16254_/Y
+ sky130_fd_sc_hd__o211ai_1
X_13466_ input70/X _13483_/B vssd1 vssd1 vccd1 vccd1 _16530_/A sky130_fd_sc_hd__and2_4
X_10678_ _18418_/Q _09726_/X _10682_/S vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14537__685 _14539__687/A vssd1 vssd1 vccd1 vccd1 _18320_/CLK sky130_fd_sc_hd__inv_2
X_15205_ _18889_/Q _18888_/Q vssd1 vssd1 vccd1 vccd1 _15955_/A sky130_fd_sc_hd__nor2_2
X_12417_ _18011_/Q vssd1 vssd1 vccd1 vccd1 _12441_/S sky130_fd_sc_hd__buf_2
X_16185_ _16290_/S vssd1 vssd1 vccd1 vccd1 _16271_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13397_ _17784_/Q _13393_/X _13396_/Y vssd1 vssd1 vccd1 vccd1 _17784_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12279_ _12279_/A vssd1 vssd1 vccd1 vccd1 _17558_/D sky130_fd_sc_hd__clkbuf_1
X_15067_ _16055_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _18474_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _13777_/X _14017_/X _14005_/X vssd1 vssd1 vccd1 vccd1 _14018_/Y sky130_fd_sc_hd__a21oi_1
X_15457__946 _15457__946/A vssd1 vssd1 vccd1 vccd1 _18633_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18826_ _18826_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_1
X_14880__797 _14881__798/A vssd1 vssd1 vccd1 vccd1 _18442_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18757_ _18757_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_1
X_15969_ _15986_/A _15973_/B _15969_/C vssd1 vssd1 vccd1 vccd1 _15969_/X sky130_fd_sc_hd__or3_1
XFILLER_247_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17708_ _17708_/CLK _17708_/D vssd1 vssd1 vccd1 vccd1 _17708_/Q sky130_fd_sc_hd__dfxtp_1
X_09490_ _19010_/Q _09489_/X _09496_/S vssd1 vssd1 vccd1 vccd1 _09491_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18688_ _18688_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _19247_/CLK _17639_/D vssd1 vssd1 vccd1 vccd1 _17639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__05076_ _17384_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05076_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15648__954 _15648__954/A vssd1 vssd1 vccd1 vccd1 _18671_/CLK sky130_fd_sc_hd__inv_2
X_15844__145 _15846__147/A vssd1 vssd1 vccd1 vccd1 _18820_/CLK sky130_fd_sc_hd__inv_2
XFILLER_247_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _19309_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_54_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09826_ _09826_/A hold5/A vssd1 vssd1 vccd1 vccd1 _09842_/S sky130_fd_sc_hd__or2_2
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09757_ _09757_/A vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18888_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_227_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03602_ clkbuf_0__03602_/X vssd1 vssd1 vccd1 vccd1 _15173__879/A sky130_fd_sc_hd__clkbuf_16
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_243_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ _11650_/A vssd1 vssd1 vccd1 vccd1 _17534_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10601_ _10601_/A vssd1 vssd1 vccd1 vccd1 _18484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11581_ _17581_/Q _10910_/X _11581_/S vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03395_ clkbuf_0__03395_/X vssd1 vssd1 vccd1 vccd1 _14808_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_195_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13320_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10532_ _18514_/Q _10333_/X _10538_/S vssd1 vssd1 vccd1 vccd1 _10533_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13251_ _14031_/A _13365_/B _13987_/B vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__and3_2
X_10463_ _10463_/A vssd1 vssd1 vccd1 vccd1 _18545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12202_ _12202_/A vssd1 vssd1 vccd1 vccd1 _12202_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ input69/X _13650_/A vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10394_ _18566_/Q vssd1 vssd1 vccd1 vccd1 _16194_/A sky130_fd_sc_hd__clkbuf_2
X_12133_ _17517_/Q _17734_/Q _12136_/S vssd1 vssd1 vccd1 vccd1 _12134_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17990_ _17991_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12064_ _12023_/X _12024_/X _12031_/X _12032_/X _12037_/S _12098_/S vssd1 vssd1 vccd1
+ vccd1 _12064_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16941_ _16939_/X _16940_/X _16979_/S vssd1 vssd1 vccd1 vccd1 _16941_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11015_ _11015_/A vssd1 vssd1 vccd1 vccd1 _18271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16872_ _18058_/Q _18050_/Q _18042_/Q _18034_/Q _16870_/X _16871_/X vssd1 vssd1 vccd1
+ vccd1 _16872_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18611_ _18611_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03160_ clkbuf_0__03160_/X vssd1 vssd1 vccd1 vccd1 _14339__526/A sky130_fd_sc_hd__clkbuf_16
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04849_ clkbuf_0__04849_/X vssd1 vssd1 vccd1 vccd1 _17073__59/A sky130_fd_sc_hd__clkbuf_16
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03191_ _14493_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03191_/X sky130_fd_sc_hd__clkbuf_16
X_18542_ _18542_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15754_/A vssd1 vssd1 vccd1 vccd1 _15754_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_90 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ _12957_/X _12966_/B vssd1 vssd1 vccd1 vccd1 _12967_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__03091_ clkbuf_0__03091_/X vssd1 vssd1 vccd1 vccd1 _14156__439/A sky130_fd_sc_hd__clkbuf_16
XFILLER_45_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _19178_/Q _19170_/Q _19202_/Q _18337_/Q _14591_/X _14592_/X vssd1 vssd1 vccd1
+ vccd1 _14705_/X sky130_fd_sc_hd__mux4_2
X_11917_ _11913_/X _11916_/X _12032_/S vssd1 vssd1 vccd1 vccd1 _11917_/X sky130_fd_sc_hd__mux2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _18477_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12894_/X _12897_/B vssd1 vssd1 vccd1 vccd1 _12898_/A sky130_fd_sc_hd__and2b_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17424_ _17474_/S vssd1 vssd1 vccd1 vccd1 _17497_/B sky130_fd_sc_hd__buf_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14636_ _14696_/A _14636_/B vssd1 vssd1 vccd1 vccd1 _14636_/Y sky130_fd_sc_hd__nor2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__and2_2
XFILLER_92_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17355_ _17355_/A vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14567_ _19048_/Q vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__buf_2
XFILLER_159_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11779_ _11779_/A _11779_/B _13128_/A vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__or3b_1
Xclkbuf_1_1__f__03993_ clkbuf_0__03993_/X vssd1 vssd1 vccd1 vccd1 _15823__129/A sky130_fd_sc_hd__clkbuf_16
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16306_ _16506_/A _16298_/Y _14623_/A _16305_/X vssd1 vssd1 vccd1 vccd1 _18924_/D
+ sky130_fd_sc_hd__o211a_4
XFILLER_174_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13518_ _13247_/X _13499_/A _13513_/X vssd1 vssd1 vccd1 vccd1 _13518_/Y sky130_fd_sc_hd__a21oi_1
X_17286_ _17286_/A vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19025_ _19027_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16237_ _18529_/Q _18537_/Q _18545_/Q _18553_/Q _10420_/A _16117_/X vssd1 vssd1 vccd1
+ vccd1 _16238_/B sky130_fd_sc_hd__mux4_2
XFILLER_127_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13449_ _13449_/A vssd1 vssd1 vccd1 vccd1 _17797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19027_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16168_ _18526_/Q _18534_/Q _18542_/Q _18550_/Q _10404_/A _16102_/X vssd1 vssd1 vccd1
+ vccd1 _16169_/B sky130_fd_sc_hd__mux4_2
XFILLER_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08990_ _18668_/Q vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__buf_2
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16099_ _18566_/Q vssd1 vssd1 vccd1 vccd1 _16152_/A sky130_fd_sc_hd__inv_2
Xclkbuf_0__04576_ _16670_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04576_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09612_/C sky130_fd_sc_hd__nand2_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18809_ _18809_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09542_ _18959_/Q _09504_/X _09542_/S vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ _09473_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__and2_1
XFILLER_240_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03180_ clkbuf_0__03180_/X vssd1 vssd1 vccd1 vccd1 _14442__609/A sky130_fd_sc_hd__clkbuf_16
XFILLER_149_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15399__900 _15400__901/A vssd1 vssd1 vccd1 vccd1 _18587_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _09824_/S vssd1 vssd1 vccd1 vccd1 _09818_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12820_ _12812_/X _12820_/B vssd1 vssd1 vccd1 vccd1 _12821_/A sky130_fd_sc_hd__and2b_1
XFILLER_41_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12758_/C _12758_/D _12755_/A vssd1 vssd1 vccd1 vccd1 _12751_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11702_ _11702_/A vssd1 vssd1 vccd1 vccd1 _11702_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15470_ _15470_/A _15643_/B vssd1 vssd1 vccd1 vccd1 _15616_/A sky130_fd_sc_hd__nor2_2
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12682_ _17612_/Q _12679_/A _12663_/X vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__o21ai_1
XFILLER_230_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _17541_/Q _09694_/A _11635_/S vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__mux2_1
X_17140_ _17289_/A _17140_/B _17140_/C vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__and3_1
XFILLER_196_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11564_ _11564_/A vssd1 vssd1 vccd1 vccd1 _17704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13303_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14831__758 _14832__759/A vssd1 vssd1 vccd1 vccd1 _18401_/CLK sky130_fd_sc_hd__inv_2
X_10515_ _10515_/A vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__clkbuf_1
X_11495_ _18047_/Q _11321_/A _11503_/S vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ _18873_/Q _16027_/C vssd1 vssd1 vccd1 vccd1 _16024_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ _17739_/Q _13218_/X _13233_/Y vssd1 vssd1 vccd1 vccd1 _17739_/D sky130_fd_sc_hd__o21a_1
X_10446_ _10123_/X _18552_/Q _10448_/S vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13165_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__buf_6
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _10377_/A vssd1 vssd1 vccd1 vccd1 _18583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12116_/A _12116_/B vssd1 vssd1 vccd1 vccd1 _12116_/X sky130_fd_sc_hd__or2_1
X_17973_ _18001_/CLK _17973_/D vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_1
X_13096_ _13096_/A _13096_/B _13096_/C _13096_/D vssd1 vssd1 vccd1 vccd1 _13097_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_46_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12047_ _12024_/X _12026_/X _12028_/X _12046_/X _12087_/S _12029_/A vssd1 vssd1 vccd1
+ vccd1 _12047_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16924_ _18247_/Q _18239_/Q _18231_/Q _18223_/Q _16849_/X _16850_/X vssd1 vssd1 vccd1
+ vccd1 _16925_/B sky130_fd_sc_hd__mux4_2
XFILLER_242_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16855_ _18180_/Q _18172_/Q _18164_/Q _18156_/Q _16813_/X _09869_/A vssd1 vssd1 vccd1
+ vccd1 _16856_/B sky130_fd_sc_hd__mux4_1
XFILLER_225_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16786_ _19135_/Q _16786_/B vssd1 vssd1 vccd1 vccd1 _16786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13998_ _13748_/A _13995_/X _13992_/X vssd1 vssd1 vccd1 vccd1 _13998_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _18525_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03174_ _14406_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03174_/X sky130_fd_sc_hd__clkbuf_16
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _12911_/X _12949_/B vssd1 vssd1 vccd1 vccd1 _12950_/A sky130_fd_sc_hd__and2b_1
XFILLER_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18456_ _18462_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _15668_/A vssd1 vssd1 vccd1 vccd1 _15668_/X sky130_fd_sc_hd__buf_1
XFILLER_233_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _14619_/A vssd1 vssd1 vccd1 vccd1 _14619_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18387_ _18387_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
X_17402__94 _17402__94/A vssd1 vssd1 vccd1 vccd1 _19307_/CLK sky130_fd_sc_hd__inv_2
X_15599_ _18654_/Q _15605_/C vssd1 vssd1 vccd1 vccd1 _15601_/B sky130_fd_sc_hd__nor2_1
X_17338_ _17323_/X _17338_/B vssd1 vssd1 vccd1 vccd1 _17339_/A sky130_fd_sc_hd__and2b_1
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03976_ clkbuf_0__03976_/X vssd1 vssd1 vccd1 vccd1 _15730_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17269_ _17274_/C _17270_/C _17268_/Y vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__a21oi_1
XFILLER_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19008_ _19008_/CLK _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04528_ clkbuf_0__04528_/X vssd1 vssd1 vccd1 vccd1 _16633_/A sky130_fd_sc_hd__clkbuf_16
X_08973_ _08988_/S vssd1 vssd1 vccd1 vccd1 _08982_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_229_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15394__896 _15395__897/A vssd1 vssd1 vccd1 vccd1 _18583_/CLK sky130_fd_sc_hd__inv_2
XFILLER_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09525_ _09525_/A vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09456_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _19047_/D sky130_fd_sc_hd__nor2_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09387_ _09387_/A vssd1 vssd1 vccd1 vccd1 _19071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03163_ clkbuf_0__03163_/X vssd1 vssd1 vccd1 vccd1 _14380_/A sky130_fd_sc_hd__clkbuf_16
X_10300_ _18613_/Q _10186_/X _10302_/S vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11280_ _18164_/Q _11279_/X _11283_/S vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03094_ clkbuf_0__03094_/X vssd1 vssd1 vccd1 vccd1 _14166_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10231_ _10231_/A vssd1 vssd1 vccd1 vccd1 _18674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _10162_/A vssd1 vssd1 vccd1 vccd1 _18701_/D sky130_fd_sc_hd__clkbuf_1
X_16703__326 _16704__327/A vssd1 vssd1 vccd1 vccd1 _19101_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14970_ _15001_/A _14970_/B vssd1 vssd1 vccd1 vccd1 _14971_/A sky130_fd_sc_hd__and2_1
X_10093_ _10093_/A vssd1 vssd1 vccd1 vccd1 _18727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13921_ _13815_/X _13908_/A _13920_/X vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_247_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13852_ _13871_/B vssd1 vssd1 vccd1 vccd1 _13863_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12803_ _12795_/X _12803_/B vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__and2b_1
X_16571_ _16571_/A vssd1 vssd1 vccd1 vccd1 _16576_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13783_ _13783_/A vssd1 vssd1 vccd1 vccd1 _13783_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _10995_/A vssd1 vssd1 vccd1 vccd1 _18280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18310_ _18310_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15522_ _18644_/Q _15516_/B _15520_/Y _18642_/Q _17842_/Q vssd1 vssd1 vccd1 vccd1
+ _15523_/D sky130_fd_sc_hd__a32o_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19290_ _19290_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18241_/CLK _18241_/D vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _17607_/D sky130_fd_sc_hd__nor2_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ _11616_/A vssd1 vssd1 vccd1 vccd1 _17566_/D sky130_fd_sc_hd__clkbuf_1
X_18172_ _18172_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_1
X_15384_ _18576_/Q _15207_/A _16064_/A _15383_/X vssd1 vssd1 vccd1 vccd1 _18576_/D
+ sky130_fd_sc_hd__o211a_1
X_12596_ _18013_/Q _17590_/Q _17589_/Q vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__and3_1
X_15801__121 _15801__121/A vssd1 vssd1 vccd1 vccd1 _18793_/CLK sky130_fd_sc_hd__inv_2
X_17123_ _17239_/A vssd1 vssd1 vccd1 vccd1 _17277_/B sky130_fd_sc_hd__clkbuf_2
X_11547_ _11547_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11563_/S sky130_fd_sc_hd__nor2_2
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11478_ _11478_/A vssd1 vssd1 vccd1 vccd1 _18055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16005_ _16003_/X _16004_/Y _15982_/X vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__a21oi_1
X_13217_ _13279_/A _13365_/B _13987_/B vssd1 vssd1 vccd1 vccd1 _13232_/A sky130_fd_sc_hd__and3_2
XFILLER_83_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10429_ _10429_/A vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__clkbuf_1
X_14197_ _14197_/A vssd1 vssd1 vccd1 vccd1 _18070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13148_ _13135_/X _13146_/X _13147_/Y _16619_/A vssd1 vssd1 vccd1 vccd1 _17724_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_151_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13079_ _17699_/Q _12846_/B _12835_/X _17698_/Q vssd1 vssd1 vccd1 vccd1 _13087_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_17956_ _18007_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16907_ _16927_/A _16907_/B vssd1 vssd1 vccd1 vccd1 _16907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17887_ _18024_/CLK _17887_/D vssd1 vssd1 vccd1 vccd1 _17887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16838_ _16819_/X _16825_/Y _16830_/Y _16833_/Y _16837_/Y vssd1 vssd1 vccd1 vccd1
+ _16838_/X sky130_fd_sc_hd__o32a_1
XFILLER_226_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16769_ _16765_/X _16766_/Y _16768_/Y _14083_/A _16762_/X vssd1 vssd1 vccd1 vccd1
+ _16770_/B sky130_fd_sc_hd__o32a_1
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ _08925_/X _19104_/Q _09312_/S vssd1 vssd1 vccd1 vccd1 _09311_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361__544 _14361__544/A vssd1 vssd1 vccd1 vccd1 _18179_/CLK sky130_fd_sc_hd__inv_2
XFILLER_206_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03157_ _14324_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03157_/X sky130_fd_sc_hd__clkbuf_16
X_18508_ _18508_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15170__876 _15172__878/A vssd1 vssd1 vccd1 vccd1 _18552_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09241_ _09972_/A _09971_/A _10403_/B vssd1 vssd1 vccd1 vccd1 _09247_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18439_ _18439_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17387__82 _17389__84/A vssd1 vssd1 vccd1 vccd1 _19295_/CLK sky130_fd_sc_hd__inv_2
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _17850_/CLK sky130_fd_sc_hd__clkbuf_16
X_16093__205 _16096__208/A vssd1 vssd1 vccd1 vccd1 _18910_/CLK sky130_fd_sc_hd__inv_2
X_09172_ _19170_/Q _09092_/X _09178_/S vssd1 vssd1 vccd1 vccd1 _09173_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16650__288 _16651__289/A vssd1 vssd1 vccd1 vccd1 _19062_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780__716 _14782__718/A vssd1 vssd1 vccd1 vccd1 _18359_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08956_ _19271_/Q _08955_/X _08959_/S vssd1 vssd1 vccd1 vccd1 _08957_/A sky130_fd_sc_hd__mux2_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _19308_/Q _08886_/X _08887_/S vssd1 vssd1 vccd1 vccd1 _08888_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09508_ _09508_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _09524_/S sky130_fd_sc_hd__nor2_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10780_/A vssd1 vssd1 vccd1 vccd1 _18375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _14627_/A vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__buf_4
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12528_/A _12533_/A _12529_/A _12449_/X _12408_/X _12560_/S vssd1 vssd1 vccd1
+ vccd1 _12451_/A sky130_fd_sc_hd__mux4_1
XFILLER_184_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15444__937 _15444__937/A vssd1 vssd1 vccd1 vccd1 _18624_/CLK sky130_fd_sc_hd__inv_2
X_11401_ _11401_/A vssd1 vssd1 vccd1 vccd1 _18115_/D sky130_fd_sc_hd__clkbuf_1
X_12381_ _12539_/B vssd1 vssd1 vccd1 vccd1 _12381_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11332_ _11332_/A vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__buf_2
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03146_ clkbuf_0__03146_/X vssd1 vssd1 vccd1 vccd1 _14268__469/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14051_ _13815_/X _14039_/A _14046_/X vssd1 vssd1 vccd1 vccd1 _14051_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_181_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11263_ _11263_/A vssd1 vssd1 vccd1 vccd1 _18170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13002_ _17682_/Q _12846_/B _12835_/X _17681_/Q vssd1 vssd1 vccd1 vccd1 _13010_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10214_ _10214_/A vssd1 vssd1 vccd1 vccd1 _18681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ _18199_/Q _11053_/X _11196_/S vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17810_ _19146_/CLK _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/Q sky130_fd_sc_hd__dfxtp_1
X_10145_ _18708_/Q _10057_/X _10149_/S vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__mux2_1
X_18790_ _18790_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _19337_/CLK _17741_/D vssd1 vssd1 vccd1 vccd1 _17741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _14961_/A _14961_/C _14962_/C vssd1 vssd1 vccd1 vccd1 _14954_/C sky130_fd_sc_hd__or3_1
X_10076_ _10157_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10092_/S sky130_fd_sc_hd__nor2_2
XFILLER_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _13394_/X _13903_/X _13894_/X vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_0__f__03979_ clkbuf_0__03979_/X vssd1 vssd1 vccd1 vccd1 _15741__1029/A sky130_fd_sc_hd__clkbuf_16
X_17672_ _19037_/CLK _17672_/D vssd1 vssd1 vccd1 vccd1 _17672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16623_ _19040_/Q _16620_/B _16622_/Y vssd1 vssd1 vccd1 vccd1 _19040_/D sky130_fd_sc_hd__o21a_1
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _17921_/Q _13829_/X _13834_/X _13826_/X vssd1 vssd1 vccd1 vccd1 _17921_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_204 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_215 _19148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_226 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ _19342_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
X_13766_ _17899_/Q _13762_/X _13765_/Y vssd1 vssd1 vccd1 vccd1 _17899_/D sky130_fd_sc_hd__o21a_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _10978_/A vssd1 vssd1 vccd1 vccd1 _18286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15505_ _18648_/Q _15505_/B _15505_/C vssd1 vssd1 vccd1 vccd1 _15525_/B sky130_fd_sc_hd__and3_1
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _12717_/A _12717_/B _12717_/C _12717_/D vssd1 vssd1 vccd1 vccd1 _12727_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_241_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19273_ _19273_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16485_ _16483_/X _16484_/Y _16469_/X vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__a21oi_1
XFILLER_231_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13697_ _17876_/Q _13683_/X _13696_/Y vssd1 vssd1 vccd1 vccd1 _17876_/D sky130_fd_sc_hd__o21a_1
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18224_ _18224_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _12647_/B _12647_/C _12647_/A vssd1 vssd1 vccd1 vccd1 _12649_/C sky130_fd_sc_hd__a21o_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18155_ _18155_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15367_ _18575_/Q _15207_/A _15270_/X _15366_/X vssd1 vssd1 vccd1 vccd1 _18575_/D
+ sky130_fd_sc_hd__o211a_1
X_12579_ _12494_/X _12485_/X _12486_/X _12487_/X _12768_/S _12538_/A vssd1 vssd1 vccd1
+ vccd1 _12580_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17106_ _17491_/B _17105_/Y _11675_/A vssd1 vssd1 vccd1 vccd1 _17106_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14318_ _14318_/A vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__buf_1
XFILLER_89_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18086_ _19337_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15298_ _15303_/A vssd1 vssd1 vccd1 vccd1 _15298_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17037_ _17037_/A vssd1 vssd1 vccd1 vccd1 _17037_/X sky130_fd_sc_hd__buf_1
XFILLER_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14249_ _14249_/A _14249_/B vssd1 vssd1 vccd1 vccd1 _14249_/Y sky130_fd_sc_hd__nor2_1
XFILLER_217_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ hold10/X vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _10220_/A hold5/A vssd1 vssd1 vccd1 vccd1 _09806_/S sky130_fd_sc_hd__nor2_2
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844__768 _14845__769/A vssd1 vssd1 vccd1 vccd1 _18413_/CLK sky130_fd_sc_hd__inv_2
X_18988_ _18993_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _13488_/A _09250_/A _11786_/A _08741_/D vssd1 vssd1 vccd1 vccd1 _13759_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_245_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17939_ _18024_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539__251 _16541__253/A vssd1 vssd1 vccd1 vccd1 _18997_/CLK sky130_fd_sc_hd__inv_2
XFILLER_224_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _18563_/Q vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09155_ _09155_/A vssd1 vssd1 vccd1 vccd1 _19178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09086_ _11601_/A vssd1 vssd1 vccd1 vccd1 _10752_/A sky130_fd_sc_hd__buf_4
XFILLER_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _18769_/Q _09959_/X _09992_/S vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__mux2_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08939_ _08939_/A vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11950_ _19245_/Q _19246_/Q _11956_/S vssd1 vssd1 vccd1 vccd1 _11950_/X sky130_fd_sc_hd__mux2_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _18990_/Q vssd1 vssd1 vccd1 vccd1 _10901_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ _13161_/X _13608_/B _13618_/Y _13619_/X vssd1 vssd1 vccd1 vccd1 _17851_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10832_ _10832_/A vssd1 vssd1 vccd1 vccd1 _18355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13551_ _17828_/Q _13557_/B vssd1 vssd1 vccd1 vccd1 _13551_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10763_ _10763_/A vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ _12502_/A vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__buf_2
XFILLER_164_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16270_ _16268_/X _16269_/X _16289_/S vssd1 vssd1 vccd1 vccd1 _16270_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13482_ _13482_/A vssd1 vssd1 vccd1 vccd1 _17807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10694_ _10694_/A vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _18934_/Q vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__clkbuf_4
X_12433_ _12431_/X _12432_/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12433_/X sky130_fd_sc_hd__mux2_1
XFILLER_240_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12364_ _17623_/Q vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14103_ _18017_/Q _14091_/X _14102_/Y vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__o21a_1
XFILLER_126_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11315_ _11159_/X _18149_/Q _11319_/S vssd1 vssd1 vccd1 vccd1 _11316_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15083_ _18483_/Q _15083_/B _16689_/B vssd1 vssd1 vccd1 vccd1 _18483_/D sky130_fd_sc_hd__nor3_1
X_12295_ _12295_/A vssd1 vssd1 vccd1 vccd1 _17563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14034_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14034_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18911_ _18911_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _11246_/A vssd1 vssd1 vccd1 vccd1 _18177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18842_ _18842_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_1
X_15121__837 _15123__839/A vssd1 vssd1 vccd1 vccd1 _18513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11177_ _11177_/A vssd1 vssd1 vccd1 vccd1 _18207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10128_ _10128_/A vssd1 vssd1 vccd1 vccd1 _18714_/D sky130_fd_sc_hd__clkbuf_1
X_18773_ _18773_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
X_15985_ _18866_/Q _15985_/B _15985_/C vssd1 vssd1 vccd1 vccd1 _15991_/B sky130_fd_sc_hd__and3_1
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17724_ _17878_/CLK _17724_/D vssd1 vssd1 vccd1 vccd1 _17724_/Q sky130_fd_sc_hd__dfxtp_1
X_14936_ _14936_/A _14936_/B _14936_/C vssd1 vssd1 vccd1 vccd1 _14964_/B sky130_fd_sc_hd__and3_1
XFILLER_76_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10059_ _10059_/A vssd1 vssd1 vccd1 vccd1 _18740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19336_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04012_ clkbuf_0__04012_/X vssd1 vssd1 vccd1 vccd1 _15863__160/A sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17655_ _18006_/CLK _17655_/D vssd1 vssd1 vccd1 vccd1 _17655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16606_ _19031_/Q _16602_/B _19032_/Q vssd1 vssd1 vccd1 vccd1 _16607_/C sky130_fd_sc_hd__a21oi_1
X_13818_ _13855_/B _14053_/B vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__and2_1
XFILLER_56_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17586_ _17586_/CLK _17586_/D vssd1 vssd1 vccd1 vccd1 _17586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19325_ _19327_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
X_16537_ _16537_/A vssd1 vssd1 vccd1 vccd1 _18995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13749_ _17893_/Q _13738_/X _13748_/Y _13741_/X vssd1 vssd1 vccd1 vccd1 _17893_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19256_ _19261_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_1
X_16468_ _18976_/Q _16468_/B vssd1 vssd1 vccd1 vccd1 _16468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18207_ _18207_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
X_19187_ _19187_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04845_ clkbuf_0__04845_/X vssd1 vssd1 vccd1 vccd1 _17048__38/A sky130_fd_sc_hd__clkbuf_16
X_16399_ _17804_/Q _16412_/B vssd1 vssd1 vccd1 vccd1 _16413_/A sky130_fd_sc_hd__nor2_1
XFILLER_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14473__634 _14473__634/A vssd1 vssd1 vccd1 vccd1 _18269_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18138_ _18138_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18069_ _18072_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ _18792_/Q _09738_/X _09913_/S vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09842_ _09697_/X _18812_/Q _09842_/S vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03589_ clkbuf_0__03589_/X vssd1 vssd1 vccd1 vccd1 _15103__822/A sky130_fd_sc_hd__clkbuf_16
XFILLER_219_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09773_ _08830_/X _18843_/Q _09781_/S vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _18887_/Q vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__buf_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09207_ _19155_/Q _09080_/X _09215_/S vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__05081_ clkbuf_0__05081_/X vssd1 vssd1 vccd1 vccd1 _17412__102/A sky130_fd_sc_hd__clkbuf_16
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09138_ _09138_/A vssd1 vssd1 vccd1 vccd1 _19183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _19200_/Q _08874_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _09070_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11100_ _09047_/X _18237_/Q _11104_/S vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ _17489_/B _12080_/B _17492_/B _12079_/X vssd1 vssd1 vccd1 vccd1 _12123_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _11031_/A vssd1 vssd1 vccd1 vccd1 _18264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12982_/A vssd1 vssd1 vccd1 vccd1 _17679_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14544_/A _14720_/X _14619_/X vssd1 vssd1 vccd1 vccd1 _14721_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11933_ _17129_/A _19225_/Q _11980_/A vssd1 vssd1 vccd1 vccd1 _11933_/X sky130_fd_sc_hd__mux2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17437_/X _17440_/B vssd1 vssd1 vccd1 vccd1 _17441_/A sky130_fd_sc_hd__and2b_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _17584_/Q _18382_/Q _18390_/Q _18424_/Q _09459_/X _09444_/A vssd1 vssd1 vccd1
+ vccd1 _14653_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _17917_/Q _11802_/A _11812_/A _17898_/Q vssd1 vssd1 vccd1 vccd1 _11865_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _17845_/Q _13608_/B vssd1 vssd1 vccd1 vccd1 _13603_/Y sky130_fd_sc_hd__nor2_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _19278_/Q _12182_/A _12180_/A _19275_/Q vssd1 vssd1 vccd1 vccd1 _17378_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_10815_ _10833_/B _11547_/A vssd1 vssd1 vccd1 vccd1 _10831_/S sky130_fd_sc_hd__nor2_2
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14583_ _14696_/A _14581_/X _14604_/A vssd1 vssd1 vccd1 vccd1 _14583_/Y sky130_fd_sc_hd__o21ai_1
X_11795_ _11839_/A vssd1 vssd1 vccd1 vccd1 _11802_/A sky130_fd_sc_hd__buf_2
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19110_ _19128_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _17822_/Q _13522_/X _13533_/Y vssd1 vssd1 vccd1 vccd1 _17822_/D sky130_fd_sc_hd__o21a_1
X_10746_ _18389_/Q _10707_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10747_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19041_ _19041_/CLK _19041_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16253_ _16291_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _17454_/A vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _10677_/A vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ _17619_/Q _17620_/Q _12426_/S vssd1 vssd1 vccd1 vccd1 _12416_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16184_ _16181_/X _16183_/X _16286_/S vssd1 vssd1 vccd1 vccd1 _16184_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _13394_/X _13395_/X _13337_/X vssd1 vssd1 vccd1 vccd1 _13396_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04592_ _16731_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04592_/X sky130_fd_sc_hd__clkbuf_16
X_15066_ _16054_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _18473_/D sky130_fd_sc_hd__nor2_1
X_12278_ _12263_/X _12278_/B vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__and2b_1
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14017_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11229_ _11150_/X _18184_/Q _11233_/S vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18825_ _18825_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18756_ _18756_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _18862_/Q _15967_/C _18863_/Q vssd1 vssd1 vccd1 vccd1 _15969_/C sky130_fd_sc_hd__a21oi_1
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17707_ _17707_/CLK _17707_/D vssd1 vssd1 vccd1 vccd1 _17707_/Q sky130_fd_sc_hd__dfxtp_1
X_14919_ _17850_/Q _14934_/A vssd1 vssd1 vccd1 vccd1 _14920_/B sky130_fd_sc_hd__xnor2_1
XFILLER_209_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15899_ _17819_/Q _17818_/Q _15917_/B vssd1 vssd1 vccd1 vccd1 _15937_/B sky130_fd_sc_hd__or3_1
X_18687_ _18687_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17638_ _18014_/CLK _17638_/D vssd1 vssd1 vccd1 vccd1 _17638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _17569_/CLK _17569_/D vssd1 vssd1 vccd1 vccd1 _17569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19308_ _19308_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19239_ _19240_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15401__902 _15403__904/A vssd1 vssd1 vccd1 vccd1 _18589_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09825_ _09825_/A vssd1 vssd1 vccd1 vccd1 _18820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09756_ _18848_/Q _09755_/X _09759_/S vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03601_ clkbuf_0__03601_/X vssd1 vssd1 vccd1 vccd1 _15167__874/A sky130_fd_sc_hd__clkbuf_16
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09687_/A vssd1 vssd1 vccd1 vccd1 _18902_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10600_ _09055_/X _18484_/Q hold19/X vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _11580_/A vssd1 vssd1 vccd1 vccd1 _17582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10531_ _10531_/A vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13250_ _14113_/A vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10462_ _18545_/Q _10336_/X _10466_/S vssd1 vssd1 vccd1 vccd1 _10463_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12201_ _12201_/A vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__buf_2
XFILLER_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _13170_/X _16060_/A _13180_/Y _13158_/X vssd1 vssd1 vccd1 vccd1 _17730_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_136_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04015_ clkbuf_0__04015_/X vssd1 vssd1 vccd1 vccd1 _15889__179/A sky130_fd_sc_hd__clkbuf_16
X_10393_ _16290_/S vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719__1011 _15720__1012/A vssd1 vssd1 vccd1 vccd1 _18728_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _12099_/S _12056_/X _12062_/X vssd1 vssd1 vccd1 vccd1 _12186_/A sky130_fd_sc_hd__o21ai_1
XFILLER_151_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16940_ _18061_/Q _18053_/Q _18045_/Q _18037_/Q _16870_/X _16871_/X vssd1 vssd1 vccd1
+ vccd1 _16940_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11014_ _09039_/X _18271_/Q _11016_/S vssd1 vssd1 vccd1 vccd1 _11015_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16871_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18610_ _18610_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04848_ clkbuf_0__04848_/X vssd1 vssd1 vccd1 vccd1 _17066__53/A sky130_fd_sc_hd__clkbuf_16
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03190_ _14487_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03190_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18541_ _18541_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12965_ _17962_/Q _17675_/Q _12976_/S vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__mux2_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03090_ clkbuf_0__03090_/X vssd1 vssd1 vccd1 vccd1 _14149__433/A sky130_fd_sc_hd__clkbuf_16
XINSDIODE2_80 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_91 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _17209_/B _19245_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14704_ _18328_/Q _14543_/A _14623_/X _14703_/X vssd1 vssd1 vccd1 vccd1 _18328_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_233_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18472_ _18921_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12896_ _17974_/Q _17662_/Q _12908_/S vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__mux2_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17771_/Q _17423_/B vssd1 vssd1 vccd1 vccd1 _17474_/S sky130_fd_sc_hd__and2_2
X_14635_ _19077_/Q _18341_/Q _17575_/Q _18793_/Q _14579_/X _14580_/X vssd1 vssd1 vccd1
+ vccd1 _14636_/B sky130_fd_sc_hd__mux4_2
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11847_ _17922_/Q _11839_/X _11840_/X _17903_/Q vssd1 vssd1 vccd1 vccd1 _11848_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17354_ _17340_/X _17354_/B vssd1 vssd1 vccd1 vccd1 _17355_/A sky130_fd_sc_hd__and2b_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14566_ _14688_/S _14566_/B vssd1 vssd1 vccd1 vccd1 _14566_/Y sky130_fd_sc_hd__nor2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _18080_/Q _13759_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__nand3_1
XFILLER_53_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03992_ clkbuf_0__03992_/X vssd1 vssd1 vccd1 vccd1 _15804__124/A sky130_fd_sc_hd__clkbuf_16
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13517_ _17817_/Q _13500_/X _13516_/Y vssd1 vssd1 vccd1 vccd1 _17817_/D sky130_fd_sc_hd__o21a_1
X_16305_ _16514_/A _16534_/A _16305_/C vssd1 vssd1 vccd1 vccd1 _16305_/X sky130_fd_sc_hd__or3_1
X_17285_ _17289_/A _17285_/B _17285_/C vssd1 vssd1 vccd1 vccd1 _17286_/A sky130_fd_sc_hd__and3_1
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _10729_/A vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15463__951 _15464__952/A vssd1 vssd1 vccd1 vccd1 _18638_/CLK sky130_fd_sc_hd__inv_2
XFILLER_173_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19024_ _19027_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_1
X_16236_ _18918_/Q _16098_/X _16235_/Y _16216_/X vssd1 vssd1 vccd1 vccd1 _18918_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13448_ _16736_/A _13448_/B vssd1 vssd1 vccd1 vccd1 _13449_/A sky130_fd_sc_hd__or2_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16312__212 _16313__213/A vssd1 vssd1 vccd1 vccd1 _18928_/CLK sky130_fd_sc_hd__inv_2
XFILLER_186_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _16276_/A vssd1 vssd1 vccd1 vccd1 _16257_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13379_ _11931_/S _13366_/S _13378_/Y vssd1 vssd1 vccd1 vccd1 _17781_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17004__353 _17005__354/A vssd1 vssd1 vccd1 vccd1 _19152_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15118_/X sky130_fd_sc_hd__buf_1
XFILLER_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16098_ _16214_/A vssd1 vssd1 vccd1 vccd1 _16098_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15049_ _18468_/Q _15049_/B vssd1 vssd1 vccd1 vccd1 _15049_/X sky130_fd_sc_hd__or2_1
Xclkbuf_0__04575_ _16664_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04575_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19251_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15850__150 _15851__151/A vssd1 vssd1 vccd1 vccd1 _18825_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _09631_/A vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__buf_4
XFILLER_205_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18808_ _18808_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09541_ _09541_/A vssd1 vssd1 vccd1 vccd1 _18960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18739_ _18739_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09472_ _19014_/Q _08844_/A _09084_/C _10770_/B vssd1 vssd1 vccd1 vccd1 _09473_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15134__847 _15134__847/A vssd1 vssd1 vccd1 vccd1 _18523_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__04009_ _15849_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04009_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030__24 _17030__24/A vssd1 vssd1 vccd1 vccd1 _19173_/CLK sky130_fd_sc_hd__inv_2
XFILLER_189_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14486__644 _14486__644/A vssd1 vssd1 vccd1 vccd1 _18279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09808_ _11637_/A hold5/A vssd1 vssd1 vccd1 vccd1 _09824_/S sky130_fd_sc_hd__or2_1
XFILLER_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09739_ _18854_/Q _09738_/X _09742_/S vssd1 vssd1 vccd1 vccd1 _09740_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _17633_/Q vssd1 vssd1 vccd1 vccd1 _12758_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11707_/S _17925_/Q vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__and2b_4
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12694_/C vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11632_ _11632_/A vssd1 vssd1 vccd1 vccd1 _17542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15408__908 _15409__909/A vssd1 vssd1 vccd1 vccd1 _18595_/CLK sky130_fd_sc_hd__inv_2
X_11563_ _17704_/Q _10910_/X _11563_/S vssd1 vssd1 vccd1 vccd1 _11564_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _14031_/A _13365_/B _14031_/B vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__and3_2
XFILLER_156_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10514_ _18522_/Q _10333_/X _10520_/S vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11494_ _11509_/S vssd1 vssd1 vccd1 vccd1 _11503_/S sky130_fd_sc_hd__buf_2
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16021_ _16019_/X _16020_/Y _16010_/X vssd1 vssd1 vccd1 vccd1 _18872_/D sky130_fd_sc_hd__a21oi_1
X_13233_ _13231_/X _13232_/X _13224_/X vssd1 vssd1 vccd1 vccd1 _13233_/Y sky130_fd_sc_hd__a21oi_1
X_10445_ _10445_/A vssd1 vssd1 vccd1 vccd1 _18553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13164_ input72/X _13431_/B vssd1 vssd1 vccd1 vccd1 _13792_/A sky130_fd_sc_hd__nand2_4
XFILLER_237_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _08786_/X _18583_/Q _10382_/S vssd1 vssd1 vccd1 vccd1 _10377_/A sky130_fd_sc_hd__mux2_1
X_12115_ _12004_/X _12008_/X _12115_/S vssd1 vssd1 vccd1 vccd1 _12116_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17972_ _18010_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_1
X_13095_ _17692_/Q _13095_/B vssd1 vssd1 vccd1 vccd1 _13096_/D sky130_fd_sc_hd__xnor2_1
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12046_ _19260_/Q _17274_/B _17276_/A _17279_/A _11931_/S _12017_/S vssd1 vssd1 vccd1
+ vccd1 _12046_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16923_ _16919_/X _16922_/X _16980_/S vssd1 vssd1 vccd1 vccd1 _16923_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16854_ _16927_/A _16854_/B vssd1 vssd1 vccd1 vccd1 _16854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14799__732 _14799__732/A vssd1 vssd1 vccd1 vccd1 _18375_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _15824_/A vssd1 vssd1 vccd1 vccd1 _15805_/X sky130_fd_sc_hd__buf_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13997_ _17978_/Q _13988_/X _13996_/Y vssd1 vssd1 vccd1 vccd1 _17978_/D sky130_fd_sc_hd__o21a_1
X_16785_ _16795_/A _16785_/B vssd1 vssd1 vccd1 vccd1 _19134_/D sky130_fd_sc_hd__nor2_1
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_2_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16339_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03173_ _14400_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03173_/X sky130_fd_sc_hd__clkbuf_16
X_18524_ _18524_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_1
X_12948_ _17967_/Q _17670_/Q _13022_/B vssd1 vssd1 vccd1 vccd1 _12949_/B sky130_fd_sc_hd__mux2_1
X_15736_ _15748_/A vssd1 vssd1 vccd1 vccd1 _15736_/X sky130_fd_sc_hd__buf_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18455_ _18455_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
X_17399__91 _17399__91/A vssd1 vssd1 vccd1 vccd1 _19304_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _17979_/Q _17657_/Q _12891_/S vssd1 vssd1 vccd1 vccd1 _12880_/B sky130_fd_sc_hd__mux2_1
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14618_ _14607_/X _14609_/Y _14611_/Y _14614_/Y _14617_/Y vssd1 vssd1 vccd1 vccd1
+ _14618_/X sky130_fd_sc_hd__o32a_1
X_15598_ _15596_/X _15597_/Y _15581_/X vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__a21oi_1
X_18386_ _18386_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17337_ _17759_/Q _19284_/Q _17350_/S vssd1 vssd1 vccd1 vccd1 _17338_/B sky130_fd_sc_hd__mux2_1
X_14549_ _19048_/Q vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03975_ clkbuf_0__03975_/X vssd1 vssd1 vccd1 vccd1 _15722__1014/A sky130_fd_sc_hd__clkbuf_16
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17268_ _17274_/C _17270_/C _17112_/B vssd1 vssd1 vccd1 vccd1 _17268_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19007_ _19007_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ _16257_/A _16219_/B vssd1 vssd1 vccd1 vccd1 _16219_/Y sky130_fd_sc_hd__nor2_1
X_17199_ _17199_/A vssd1 vssd1 vccd1 vccd1 _19241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08972_ _09508_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _08988_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_1_1__f__04527_ clkbuf_0__04527_/X vssd1 vssd1 vccd1 vccd1 _16547__258/A sky130_fd_sc_hd__clkbuf_16
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_15691__989 _15691__989/A vssd1 vssd1 vccd1 vccd1 _18706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03409_ clkbuf_0__03409_/X vssd1 vssd1 vccd1 vccd1 _14814__744/A sky130_fd_sc_hd__clkbuf_16
XFILLER_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09524_ _18997_/Q _09504_/X _09524_/S vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09444_/A _09444_/B _09477_/C vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__o21ai_1
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16319__218 _16320__219/A vssd1 vssd1 vccd1 vccd1 _18934_/CLK sky130_fd_sc_hd__inv_2
XFILLER_212_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15718__1010 _15720__1012/A vssd1 vssd1 vccd1 vccd1 _18727_/CLK sky130_fd_sc_hd__inv_2
X_09386_ _19071_/Q _08955_/X _09388_/S vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03162_ clkbuf_0__03162_/X vssd1 vssd1 vccd1 vccd1 _14352__537/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15857__156 _15859__158/A vssd1 vssd1 vccd1 vccd1 _18831_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03093_ clkbuf_0__03093_/X vssd1 vssd1 vccd1 vccd1 _14293_/A sky130_fd_sc_hd__clkbuf_16
X_10230_ _18674_/Q _09758_/X _10230_/S vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ _18701_/Q _10054_/X _10167_/S vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _18727_/Q _10072_/X _10092_/S vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13920_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13920_/X sky130_fd_sc_hd__buf_2
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13851_ input71/X vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__inv_2
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12802_ _17643_/Q _17992_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12803_/B sky130_fd_sc_hd__mux2_1
XFILLER_210_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16570_ _16570_/A vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__clkbuf_2
X_13782_ _17904_/Q _13770_/X _13781_/Y vssd1 vssd1 vccd1 vccd1 _17904_/D sky130_fd_sc_hd__o21a_1
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _18280_/Q _09130_/X _10998_/S vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12733_ _12737_/B _12737_/C _12737_/D vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__and3_1
XFILLER_231_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15521_ _15516_/B _15520_/Y _18644_/Q vssd1 vssd1 vccd1 vccd1 _15523_/C sky130_fd_sc_hd__a21oi_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ _18240_/CLK _18240_/D vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
X_12664_ _17607_/Q _12658_/X _12663_/X vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__o21ai_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _17566_/Q _10710_/A _11617_/S vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15383_ _15244_/A _15372_/X _15382_/X _15267_/A vssd1 vssd1 vccd1 vccd1 _15383_/X
+ sky130_fd_sc_hd__a211o_1
X_18171_ _18171_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
X_12595_ _12595_/A vssd1 vssd1 vccd1 vccd1 _17589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17122_ _17117_/A _17117_/B _17117_/C _19222_/Q vssd1 vssd1 vccd1 vccd1 _17124_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _11546_/A vssd1 vssd1 vccd1 vccd1 _17712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11477_ _09119_/X _18055_/Q _11485_/S vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16004_ _18869_/Q _16020_/B vssd1 vssd1 vccd1 vccd1 _16004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13216_ _18066_/Q _13216_/B _13216_/C vssd1 vssd1 vccd1 vccd1 _13987_/B sky130_fd_sc_hd__and3_2
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _10424_/X _10428_/B _10433_/C vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__and3b_1
X_14196_ _18070_/Q input50/X _14196_/S vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13147_ _17724_/Q _13147_/B vssd1 vssd1 vccd1 vccd1 _13147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10359_/A vssd1 vssd1 vccd1 vccd1 _18591_/D sky130_fd_sc_hd__clkbuf_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13078_/A vssd1 vssd1 vccd1 vccd1 _17702_/D sky130_fd_sc_hd__clkbuf_1
X_17955_ _18007_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12029_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16906_ _18206_/Q _18126_/Q _19183_/Q _18254_/Q _16827_/X _16828_/X vssd1 vssd1 vccd1
+ vccd1 _16907_/B sky130_fd_sc_hd__mux4_1
X_17886_ _18024_/CLK _17886_/D vssd1 vssd1 vccd1 vccd1 _17886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ _09868_/X _16835_/X _16836_/X vssd1 vssd1 vccd1 vccd1 _16837_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_226_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16768_ _16783_/A _16768_/B vssd1 vssd1 vccd1 vccd1 _16768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03156_ _14318_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03156_/X sky130_fd_sc_hd__clkbuf_16
X_18507_ _18507_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09240_ _18559_/Q vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18438_ _18438_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _09171_/A vssd1 vssd1 vccd1 vccd1 _19171_/D sky130_fd_sc_hd__clkbuf_1
X_18369_ _18369_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03989_ _15786_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03989_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ _09685_/A vssd1 vssd1 vccd1 vccd1 _08955_/X sky130_fd_sc_hd__buf_4
XFILLER_131_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08886_ _18987_/Q vssd1 vssd1 vccd1 vccd1 _08886_/X sky130_fd_sc_hd__buf_4
XFILLER_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _10219_/B _09789_/A _09377_/A vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__or3b_4
XFILLER_213_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15863__160 _15863__160/A vssd1 vssd1 vccd1 vccd1 _18835_/CLK sky130_fd_sc_hd__inv_2
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09438_ _19046_/Q vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _19078_/Q _09104_/X _09369_/S vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _11344_/X _18115_/Q _11400_/S vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _12376_/X _12379_/X _12448_/A vssd1 vssd1 vccd1 vccd1 _12539_/B sky130_fd_sc_hd__mux2_1
XFILLER_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17393__86 _17396__89/A vssd1 vssd1 vccd1 vccd1 _19299_/CLK sky130_fd_sc_hd__inv_2
X_14338__525 _14339__526/A vssd1 vssd1 vccd1 vccd1 _18160_/CLK sky130_fd_sc_hd__inv_2
XFILLER_138_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11331_ _11331_/A vssd1 vssd1 vccd1 vccd1 _18144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03145_ clkbuf_0__03145_/X vssd1 vssd1 vccd1 vccd1 _14287_/A sky130_fd_sc_hd__clkbuf_16
X_14050_ _17998_/Q _14033_/X _14049_/Y vssd1 vssd1 vccd1 vccd1 _17998_/D sky130_fd_sc_hd__o21a_1
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11262_ _18170_/Q _11259_/X _11274_/S vssd1 vssd1 vccd1 vccd1 _11263_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13001_ _13001_/A vssd1 vssd1 vccd1 vccd1 _17685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10213_ _18681_/Q _09761_/X hold6/X vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ _11193_/A vssd1 vssd1 vccd1 vccd1 _18200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10144_ _10144_/A vssd1 vssd1 vccd1 vccd1 _18709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15741__1029 _15741__1029/A vssd1 vssd1 vccd1 vccd1 _18746_/CLK sky130_fd_sc_hd__inv_2
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _19336_/CLK _17740_/D vssd1 vssd1 vccd1 vccd1 _17740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14952_ _15005_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14962_/C sky130_fd_sc_hd__nor2_1
X_10075_ _18562_/Q _10075_/B _10049_/A vssd1 vssd1 vccd1 vccd1 _10564_/B sky130_fd_sc_hd__or3b_2
XFILLER_248_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03978_ clkbuf_0__03978_/X vssd1 vssd1 vccd1 vccd1 _15735__1024/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _13908_/A vssd1 vssd1 vccd1 vccd1 _13903_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17671_ _19037_/CLK _17671_/D vssd1 vssd1 vccd1 vccd1 _17671_/Q sky130_fd_sc_hd__dfxtp_1
X_14883_ _14883_/A vssd1 vssd1 vccd1 vccd1 _14883_/X sky130_fd_sc_hd__buf_1
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16622_ _19040_/Q _16620_/B _14184_/A vssd1 vssd1 vccd1 vccd1 _16622_/Y sky130_fd_sc_hd__a21oi_1
X_13834_ input60/X _13845_/B vssd1 vssd1 vccd1 vccd1 _13834_/X sky130_fd_sc_hd__and2_1
XINSDIODE2_205 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_216 _18846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19341_ _19341_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
X_13765_ _13709_/A _13762_/X _13701_/X vssd1 vssd1 vccd1 vccd1 _13765_/Y sky130_fd_sc_hd__a21oi_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10977_ _18286_/Q _09758_/X _10977_/S vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ _17837_/Q _15511_/A _17836_/Q vssd1 vssd1 vccd1 vccd1 _15505_/C sky130_fd_sc_hd__o21ai_1
X_12716_ _12716_/A _12716_/B vssd1 vssd1 vccd1 vccd1 _17622_/D sky130_fd_sc_hd__nor2_1
XFILLER_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19272_ _19272_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13696_ _13268_/X _13688_/X _13689_/X vssd1 vssd1 vccd1 vccd1 _13696_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16484_ _18979_/Q _16499_/B vssd1 vssd1 vccd1 vccd1 _16484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ _18223_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
X_12647_ _12647_/A _12647_/B _12647_/C vssd1 vssd1 vccd1 vccd1 _12647_/X sky130_fd_sc_hd__and3_1
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15435_ _15441_/A vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__buf_1
XFILLER_15_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18154_ _18154_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
X_15366_ _15244_/A _15355_/X _15365_/X _15267_/A vssd1 vssd1 vccd1 vccd1 _15366_/X
+ sky130_fd_sc_hd__a211o_1
X_12578_ _12489_/X _12513_/X _12557_/X _12577_/X _12569_/S _12568_/A vssd1 vssd1 vccd1
+ vccd1 _12578_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _17775_/Q _17774_/Q _17773_/Q vssd1 vssd1 vccd1 vccd1 _17105_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11545_/S sky130_fd_sc_hd__or2_2
XFILLER_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18085_ _19337_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
X_15297_ _15292_/X _15294_/X _15295_/X _15296_/X _15281_/X _09600_/X vssd1 vssd1 vccd1
+ vccd1 _15297_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _16097_/B _14242_/X _14247_/X vssd1 vssd1 vccd1 vccd1 _18088_/D sky130_fd_sc_hd__o21a_1
XFILLER_217_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__08201_ clkbuf_0__08201_/X vssd1 vssd1 vccd1 vccd1 _14138__424/A sky130_fd_sc_hd__clkbuf_16
XFILLER_171_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _18987_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _18078_/Q _11786_/A _18079_/Q vssd1 vssd1 vccd1 vccd1 _08741_/D sky130_fd_sc_hd__a21oi_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _18024_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17869_ _18031_/CLK _17869_/D vssd1 vssd1 vccd1 vccd1 _17869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ _18480_/Q vssd1 vssd1 vccd1 vccd1 _09223_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09154_ _19178_/Q _09092_/X _09160_/S vssd1 vssd1 vccd1 vccd1 _09155_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _09476_/A _09449_/A _09480_/A vssd1 vssd1 vccd1 vccd1 _11601_/A sky130_fd_sc_hd__or3b_4
XFILLER_190_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _09987_/A vssd1 vssd1 vccd1 vccd1 _18770_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ _08937_/X _19293_/Q _08942_/S vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__mux2_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _19314_/Q _08868_/X _08878_/S vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__mux2_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ _10900_/A vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10831_ _18355_/Q _10812_/X _10831_/S vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13550_ _13559_/S vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ _18382_/Q _10704_/X _10762_/S vssd1 vssd1 vccd1 vccd1 _10763_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _12421_/X _12500_/X _12433_/X _12418_/X _12567_/S _12408_/A vssd1 vssd1 vccd1
+ vccd1 _12501_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _13560_/A _13481_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__or2_1
X_10693_ _18410_/Q _10690_/X _10705_/S vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668__303 _16669__304/A vssd1 vssd1 vccd1 vccd1 _19077_/CLK sky130_fd_sc_hd__inv_2
X_15220_ _15303_/A vssd1 vssd1 vccd1 vccd1 _15220_/X sky130_fd_sc_hd__clkbuf_4
X_12432_ _17615_/Q _17616_/Q _12432_/S vssd1 vssd1 vccd1 vccd1 _12432_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _17622_/Q vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _13724_/A _14099_/X _14096_/X vssd1 vssd1 vccd1 vccd1 _14102_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11314_ _11314_/A vssd1 vssd1 vccd1 vccd1 _18150_/D sky130_fd_sc_hd__clkbuf_1
X_15082_ _19109_/Q _19108_/Q vssd1 vssd1 vccd1 vccd1 _16689_/B sky130_fd_sc_hd__nor2_1
X_12294_ _12280_/X _12294_/B vssd1 vssd1 vccd1 vccd1 _12295_/A sky130_fd_sc_hd__and2b_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14033_ _14039_/A vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18910_ _18910_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11245_ _11147_/X _18177_/Q _11251_/S vssd1 vssd1 vccd1 vccd1 _11246_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18841_ _18841_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_1
X_11176_ _11153_/X _18207_/Q _11178_/S vssd1 vssd1 vccd1 vccd1 _11177_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10127_ _10126_/X _18714_/Q _10127_/S vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18772_ _18772_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _15985_/B _15985_/C _18866_/Q vssd1 vssd1 vccd1 vccd1 _15986_/B sky130_fd_sc_hd__a21oi_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ _18031_/CLK _17723_/D vssd1 vssd1 vccd1 vccd1 _17723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ _18462_/Q _14935_/B vssd1 vssd1 vccd1 vccd1 _14962_/A sky130_fd_sc_hd__xnor2_1
X_10058_ _18740_/Q _10057_/X _10064_/S vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04011_ clkbuf_0__04011_/X vssd1 vssd1 vccd1 vccd1 _15880_/A sky130_fd_sc_hd__clkbuf_16
X_17654_ _18006_/CLK _17654_/D vssd1 vssd1 vccd1 vccd1 _17654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14507__661 _14510__664/A vssd1 vssd1 vccd1 vccd1 _18296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_224_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16605_ _19031_/Q _16602_/B _16604_/Y vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13817_ _17916_/Q _13797_/X _13816_/Y vssd1 vssd1 vccd1 vccd1 _17916_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17585_ _17585_/CLK _17585_/D vssd1 vssd1 vccd1 vccd1 _17585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19324_ _19327_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_69_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17935_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16536_ _16534_/X _16536_/B _16536_/C vssd1 vssd1 vccd1 vccd1 _16537_/A sky130_fd_sc_hd__and3b_1
XFILLER_204_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13748_ _13748_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13748_/Y sky130_fd_sc_hd__nor2_1
XFILLER_232_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19255_ _19261_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16467_ _16467_/A _16467_/B _16473_/B vssd1 vssd1 vccd1 vccd1 _16467_/X sky130_fd_sc_hd__or3_1
X_13679_ _13247_/X _13666_/A _13674_/X vssd1 vssd1 vccd1 vccd1 _13679_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18206_ _18206_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__04844_ clkbuf_0__04844_/X vssd1 vssd1 vccd1 vccd1 _17068_/A sky130_fd_sc_hd__clkbuf_16
X_19186_ _19186_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _16397_/B _16397_/C _18974_/Q vssd1 vssd1 vccd1 vccd1 _16418_/B sky130_fd_sc_hd__a21oi_1
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18137_ _18137_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
X_14850__773 _14850__773/A vssd1 vssd1 vccd1 vccd1 _18418_/CLK sky130_fd_sc_hd__inv_2
X_15349_ _15244_/X _15338_/X _15348_/X _15267_/X vssd1 vssd1 vccd1 vccd1 _15349_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18068_ _18870_/CLK _18068_/D vssd1 vssd1 vccd1 vccd1 _18068_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17019_ _17037_/A vssd1 vssd1 vccd1 vccd1 _17019_/X sky130_fd_sc_hd__buf_1
X_09910_ _09910_/A vssd1 vssd1 vccd1 vccd1 _18793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09841_ _09841_/A vssd1 vssd1 vccd1 vccd1 _18813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03588_ clkbuf_0__03588_/X vssd1 vssd1 vccd1 vccd1 _15095__815/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ _09787_/S vssd1 vssd1 vccd1 vccd1 _09781_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14892__807 _14892__807/A vssd1 vssd1 vccd1 vccd1 _18452_/CLK sky130_fd_sc_hd__inv_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408__581 _14410__583/A vssd1 vssd1 vccd1 vccd1 _18216_/CLK sky130_fd_sc_hd__inv_2
XFILLER_242_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ _09221_/S vssd1 vssd1 vccd1 vccd1 _09215_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_210_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15740__1028 _15741__1029/A vssd1 vssd1 vccd1 vccd1 _18745_/CLK sky130_fd_sc_hd__inv_2
XFILLER_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__05080_ clkbuf_0__05080_/X vssd1 vssd1 vccd1 vccd1 _17408__99/A sky130_fd_sc_hd__clkbuf_16
XFILLER_182_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09137_ _19183_/Q _09136_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14751__693 _14752__694/A vssd1 vssd1 vccd1 vccd1 _18336_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _09068_/A vssd1 vssd1 vccd1 vccd1 _19201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11030_ _18264_/Q _09130_/X _11034_/S vssd1 vssd1 vccd1 vccd1 _11031_/A sky130_fd_sc_hd__mux2_1
X_16663__299 _16663__299/A vssd1 vssd1 vccd1 vccd1 _19073_/CLK sky130_fd_sc_hd__inv_2
XFILLER_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12975_/X _12981_/B vssd1 vssd1 vccd1 vccd1 _12982_/A sky130_fd_sc_hd__and2b_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14607_/X _14713_/Y _14715_/Y _14717_/Y _14719_/Y vssd1 vssd1 vccd1 vccd1
+ _14720_/X sky130_fd_sc_hd__o32a_1
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11932_ _19224_/Q vssd1 vssd1 vccd1 vccd1 _17129_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _11863_/A vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14651_ _14651_/A _14651_/B vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14793__727 _14793__727/A vssd1 vssd1 vccd1 vccd1 _18370_/CLK sky130_fd_sc_hd__inv_2
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13602_ _13611_/S vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__clkbuf_2
X_10814_ _10814_/A vssd1 vssd1 vccd1 vccd1 _18363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _19284_/Q _17487_/B vssd1 vssd1 vccd1 vccd1 _17378_/A sky130_fd_sc_hd__xnor2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11794_ _11837_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14582_ _19049_/Q vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16321_ _16333_/A vssd1 vssd1 vccd1 vccd1 _16321_/X sky130_fd_sc_hd__buf_1
XFILLER_242_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13533_ _13407_/X _13523_/X _13532_/X vssd1 vssd1 vccd1 vccd1 _13533_/Y sky130_fd_sc_hd__a21oi_1
X_10745_ _10745_/A vssd1 vssd1 vccd1 vccd1 _18390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19040_ _19040_/CLK _19040_/D vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16252_ _16248_/X _16251_/X _16271_/S vssd1 vssd1 vccd1 vccd1 _16253_/B sky130_fd_sc_hd__mux2_1
X_13464_ _16061_/A _13463_/B _13463_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _17802_/D
+ sky130_fd_sc_hd__a211oi_1
X_10676_ _18419_/Q _09723_/X _10682_/S vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12415_ _12707_/B _17618_/Q _12432_/S vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13395_ _13395_/A vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__clkbuf_2
X_16183_ _18777_/Q _18635_/Q _18785_/Q _18619_/Q _16158_/X _16182_/X vssd1 vssd1 vccd1
+ vccd1 _16183_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__04591_ _16725_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04591_/X sky130_fd_sc_hd__clkbuf_16
X_15065_ _15177_/A vssd1 vssd1 vccd1 vccd1 _15070_/B sky130_fd_sc_hd__clkbuf_2
X_12277_ _17558_/Q _18019_/Q _12287_/S vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__mux2_1
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14016_ _17985_/Q _14011_/X _14015_/Y vssd1 vssd1 vccd1 vccd1 _17985_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _11228_/A vssd1 vssd1 vccd1 vccd1 _18185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18824_ _18824_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ _11338_/A vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__buf_2
XFILLER_68_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18755_ _18755_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15967_ _18863_/Q _18862_/Q _15967_/C vssd1 vssd1 vccd1 vccd1 _15973_/B sky130_fd_sc_hd__and3_1
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17706_ _17706_/CLK _17706_/D vssd1 vssd1 vccd1 vccd1 _17706_/Q sky130_fd_sc_hd__dfxtp_1
X_14918_ _17851_/Q _14938_/A vssd1 vssd1 vccd1 vccd1 _14934_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18686_ _18686_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _17821_/Q _17820_/Q _15932_/B vssd1 vssd1 vccd1 vccd1 _15917_/B sky130_fd_sc_hd__or3_2
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17637_ _18014_/CLK _17637_/D vssd1 vssd1 vccd1 vccd1 _17637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ _17568_/CLK _17568_/D vssd1 vssd1 vccd1 vccd1 _17568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19307_ _19307_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ _16519_/A vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19238_ _19248_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19169_ _19169_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03809_ _15461_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03809_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_160_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09824_ _09697_/X _18820_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09755_ _18884_/Q vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03600_ clkbuf_0__03600_/X vssd1 vssd1 vccd1 vccd1 _15158__866/A sky130_fd_sc_hd__clkbuf_16
X_09686_ _09685_/X _18902_/Q _09689_/S vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__mux2_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14857__779 _14857__779/A vssd1 vssd1 vccd1 vccd1 _18424_/CLK sky130_fd_sc_hd__inv_2
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10530_ _18515_/Q _10328_/X _10538_/S vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A vssd1 vssd1 vccd1 vccd1 _18546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12200_ _17516_/Q _12187_/X _12199_/X _17526_/Q vssd1 vssd1 vccd1 vccd1 _12217_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ _17730_/Q _13180_/B vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__04014_ clkbuf_0__04014_/X vssd1 vssd1 vccd1 vccd1 _15878__173/A sky130_fd_sc_hd__clkbuf_16
X_10392_ _18567_/Q vssd1 vssd1 vccd1 vccd1 _16290_/S sky130_fd_sc_hd__buf_2
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ _12131_/A vssd1 vssd1 vccd1 vccd1 _17516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _12075_/A _12057_/X _12061_/X _12069_/A vssd1 vssd1 vccd1 vccd1 _12062_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ _11013_/A vssd1 vssd1 vccd1 vccd1 _18272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _16893_/A vssd1 vssd1 vccd1 vccd1 _16870_/X sky130_fd_sc_hd__buf_2
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04847_ clkbuf_0__04847_/X vssd1 vssd1 vccd1 vccd1 _17058__46/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _18540_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_70 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ _12964_/A vssd1 vssd1 vccd1 vccd1 _17674_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801__734 _14801__734/A vssd1 vssd1 vccd1 vccd1 _18377_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_81 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_92 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14544_/X _14692_/X _14702_/Y vssd1 vssd1 vccd1 vccd1 _14703_/X sky130_fd_sc_hd__a21o_1
X_11915_ _11975_/S vssd1 vssd1 vccd1 vccd1 _12025_/S sky130_fd_sc_hd__buf_2
X_18471_ _18921_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12915_/S vssd1 vssd1 vccd1 vccd1 _12908_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14634_ _14732_/A _14634_/B vssd1 vssd1 vccd1 vccd1 _14634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11846_ _11846_/A vssd1 vssd1 vccd1 vccd1 _11846_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17754_/Q _19289_/Q _17357_/S vssd1 vssd1 vccd1 vccd1 _17354_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11786_/A _13386_/B _13386_/C _11776_/Y vssd1 vssd1 vccd1 vccd1 _13874_/C
+ sky130_fd_sc_hd__a211oi_2
X_14758__699 _14758__699/A vssd1 vssd1 vccd1 vccd1 _18342_/CLK sky130_fd_sc_hd__inv_2
X_14565_ _19148_/Q _18413_/Q _18307_/Q _18291_/Q _14563_/X _14564_/X vssd1 vssd1 vccd1
+ vccd1 _14566_/B sky130_fd_sc_hd__mux4_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03991_ clkbuf_0__03991_/X vssd1 vssd1 vccd1 vccd1 _15796__117/A sky130_fd_sc_hd__clkbuf_16
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16304_ _16302_/X _16303_/X _18986_/Q vssd1 vssd1 vccd1 vccd1 _16305_/C sky130_fd_sc_hd__mux2_1
X_13516_ _13244_/X _13499_/A _13513_/X vssd1 vssd1 vccd1 vccd1 _13516_/Y sky130_fd_sc_hd__a21oi_1
X_10728_ _18397_/Q _10707_/X _10732_/S vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__mux2_1
X_17284_ _17288_/B _17288_/C _17284_/C vssd1 vssd1 vccd1 vccd1 _17285_/C sky130_fd_sc_hd__nand3_1
XFILLER_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19023_ _19027_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16235_ _16190_/X _16226_/X _16234_/Y _16214_/X vssd1 vssd1 vccd1 vccd1 _16235_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_220_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13447_ _17797_/Q _13446_/X _13447_/S vssd1 vssd1 vccd1 vccd1 _13448_/B sky130_fd_sc_hd__mux2_1
X_10659_ _10659_/A vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13378_ _13271_/X _13366_/S _13337_/X vssd1 vssd1 vccd1 vccd1 _13378_/Y sky130_fd_sc_hd__a21oi_2
X_16166_ _18915_/Q _16098_/X _16165_/Y _14247_/X vssd1 vssd1 vccd1 vccd1 _18915_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16097_ _16097_/A _16097_/B vssd1 vssd1 vccd1 vccd1 _16214_/A sky130_fd_sc_hd__and2_1
XFILLER_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15048_ _18468_/Q _15049_/B vssd1 vssd1 vccd1 vccd1 _15048_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04574_ _16658_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04574_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18807_ _18807_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_84_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _17840_/CLK sky130_fd_sc_hd__clkbuf_16
X_09540_ _18960_/Q _09501_/X _09542_/S vssd1 vssd1 vccd1 vccd1 _09541_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18738_ _18738_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19133_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09471_ _10770_/A _09473_/A _10662_/S vssd1 vssd1 vccd1 vccd1 _19045_/D sky130_fd_sc_hd__a21o_1
X_18669_ _18670_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17015__11 _17016__12/A vssd1 vssd1 vccd1 vccd1 _19160_/CLK sky130_fd_sc_hd__inv_2
XFILLER_224_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04008_ _15843_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04008_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_211_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09807_ _09807_/A vssd1 vssd1 vccd1 vccd1 _18828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09738_ _10710_/A vssd1 vssd1 vccd1 vccd1 _09738_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_228_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ _09669_/A vssd1 vssd1 vccd1 vccd1 _18908_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _17722_/Q vssd1 vssd1 vccd1 vccd1 _11707_/S sky130_fd_sc_hd__buf_4
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12680_ _17612_/Q _17611_/Q _12680_/C _12680_/D vssd1 vssd1 vccd1 vccd1 _12694_/C
+ sky130_fd_sc_hd__and4_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _17542_/Q _09691_/A _11635_/S vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11562_ _11562_/A vssd1 vssd1 vccd1 vccd1 _17705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13301_ _17760_/Q _13282_/X _13300_/Y vssd1 vssd1 vccd1 vccd1 _17760_/D sky130_fd_sc_hd__o21a_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10513_ _10513_/A vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__clkbuf_1
X_14281_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14281_/X sky130_fd_sc_hd__buf_1
XFILLER_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11493_ _11493_/A hold23/X vssd1 vssd1 vccd1 vccd1 _11509_/S sky130_fd_sc_hd__nor2_2
X_16077__192 _16077__192/A vssd1 vssd1 vccd1 vccd1 _18897_/CLK sky130_fd_sc_hd__inv_2
XFILLER_183_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13232_ _13232_/A vssd1 vssd1 vccd1 vccd1 _13232_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16020_ _18872_/Q _16020_/B vssd1 vssd1 vccd1 vccd1 _16020_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10444_ _10120_/X _18553_/Q _10448_/S vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _13135_/X _13161_/X _13162_/Y _13158_/X vssd1 vssd1 vccd1 vccd1 _17727_/D
+ sky130_fd_sc_hd__a211oi_1
X_10375_ _10375_/A vssd1 vssd1 vccd1 vccd1 _18584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12114_ _12108_/Y _12110_/Y _12112_/Y _12113_/Y _12075_/A _12022_/A vssd1 vssd1 vccd1
+ vccd1 _12205_/A sky130_fd_sc_hd__mux4_1
XFILLER_124_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17971_ _18010_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
X_13094_ _17691_/Q _13094_/B vssd1 vssd1 vccd1 vccd1 _13096_/C sky130_fd_sc_hd__xnor2_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12045_ _12108_/A _12113_/A _12045_/S vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__mux2_1
X_16922_ _16920_/X _16921_/X _16979_/S vssd1 vssd1 vccd1 vccd1 _16922_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16853_ _18204_/Q _18124_/Q _19181_/Q _18252_/Q _16827_/X _16828_/X vssd1 vssd1 vccd1
+ vccd1 _16854_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16784_ _16765_/X _16781_/Y _16783_/Y _13746_/A _16762_/X vssd1 vssd1 vccd1 vccd1
+ _16785_/B sky130_fd_sc_hd__o32a_1
XFILLER_207_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13996_ _13529_/X _13995_/X _13992_/X vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_168_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03172_ _14394_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03172_/X sky130_fd_sc_hd__clkbuf_16
X_18523_ _18523_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12947_ _12999_/S vssd1 vssd1 vccd1 vccd1 _13022_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18454_ _18462_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12878_ _12915_/S vssd1 vssd1 vccd1 vccd1 _12891_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14617_ _14651_/A _14616_/X _14561_/X vssd1 vssd1 vccd1 vccd1 _14617_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11829_ _13279_/A vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__clkbuf_2
X_18385_ _18385_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_15597_ _18653_/Q _15597_/B vssd1 vssd1 vccd1 vccd1 _15597_/Y sky130_fd_sc_hd__nand2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17336_ _17357_/S vssd1 vssd1 vccd1 vccd1 _17350_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14548_ _18403_/Q _18395_/Q _19308_/Q _17712_/Q _14641_/A _14546_/X vssd1 vssd1 vccd1
+ vccd1 _14548_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03974_ clkbuf_0__03974_/X vssd1 vssd1 vccd1 vccd1 _15714__1007/A sky130_fd_sc_hd__clkbuf_16
XFILLER_202_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17267_ _19260_/Q vssd1 vssd1 vccd1 vccd1 _17274_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_146_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19006_ _19006_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_1
X_16218_ _18528_/Q _18536_/Q _18544_/Q _18552_/Q _10420_/A _16117_/X vssd1 vssd1 vccd1
+ vccd1 _16219_/B sky130_fd_sc_hd__mux4_2
XFILLER_179_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17198_ _17195_/X _17235_/B _17198_/C vssd1 vssd1 vccd1 vccd1 _17199_/A sky130_fd_sc_hd__and3b_1
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16149_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _09377_/A _09639_/A _10219_/C vssd1 vssd1 vccd1 vccd1 _10967_/B sky130_fd_sc_hd__or3_4
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15140__852 _15142__854/A vssd1 vssd1 vccd1 vccd1 _18528_/CLK sky130_fd_sc_hd__inv_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_229_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03408_ clkbuf_0__03408_/X vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14288__485 _14290__487/A vssd1 vssd1 vccd1 vccd1 _18120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09523_ _09523_/A vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09454_ _09454_/A vssd1 vssd1 vccd1 vccd1 _19048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09385_ _09385_/A vssd1 vssd1 vccd1 vccd1 _19072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329__391 _12329__391/A vssd1 vssd1 vccd1 vccd1 _17572_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03161_ clkbuf_0__03161_/X vssd1 vssd1 vccd1 vccd1 _14348__534/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03092_ clkbuf_0__03092_/X vssd1 vssd1 vccd1 vccd1 _15447_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _10160_/A vssd1 vssd1 vccd1 vccd1 _18702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10091_ _10091_/A vssd1 vssd1 vccd1 vccd1 _18728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _13871_/B vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15414__913 _15415__914/A vssd1 vssd1 vccd1 vccd1 _18600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12801_ _12801_/A vssd1 vssd1 vccd1 vccd1 _17642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13781_ _13669_/X _13778_/X _13774_/X vssd1 vssd1 vccd1 vccd1 _13781_/Y sky130_fd_sc_hd__a21oi_1
X_10993_ _10993_/A vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15520_ _17842_/Q _17841_/Q _17840_/Q vssd1 vssd1 vccd1 vccd1 _15520_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12732_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _17627_/D sky130_fd_sc_hd__nor2_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12695_/A vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14501__656 _14503__658/A vssd1 vssd1 vccd1 vccd1 _18291_/CLK sky130_fd_sc_hd__inv_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18170_ _18170_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
X_11614_ _11614_/A vssd1 vssd1 vccd1 vccd1 _17567_/D sky130_fd_sc_hd__clkbuf_1
X_15382_ _15376_/X _15381_/X _09620_/A vssd1 vssd1 vccd1 vccd1 _15382_/X sky130_fd_sc_hd__o21a_1
X_12594_ _17589_/Q _12755_/A vssd1 vssd1 vccd1 vccd1 _12595_/A sky130_fd_sc_hd__and2b_1
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _17133_/D vssd1 vssd1 vccd1 vccd1 _17129_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ _08886_/X _17712_/Q _11545_/S vssd1 vssd1 vccd1 vccd1 _11546_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11476_ _11491_/S vssd1 vssd1 vccd1 vccd1 _11485_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16003_ _16024_/A _16003_/B _16007_/B vssd1 vssd1 vccd1 vccd1 _16003_/X sky130_fd_sc_hd__or3_1
X_13215_ _14113_/B vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10427_ _10424_/B _10432_/A _10436_/A _10424_/A vssd1 vssd1 vccd1 vccd1 _10428_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _14195_/A vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13146_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__buf_6
X_10358_ _18591_/Q _09723_/X _10364_/S vssd1 vssd1 vccd1 vccd1 _10359_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13066_/X _13077_/B vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__and2b_1
X_17954_ _18007_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _10289_/A vssd1 vssd1 vccd1 vccd1 _18618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12028_ _17252_/A _19257_/Q _17262_/B _17264_/A _11931_/S _11981_/X vssd1 vssd1 vccd1
+ vccd1 _12028_/X sky130_fd_sc_hd__mux4_1
X_16905_ _16963_/A _16905_/B vssd1 vssd1 vccd1 vccd1 _16905_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17885_ _18001_/CLK _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16836_ _18810_/Q vssd1 vssd1 vccd1 vccd1 _16836_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16767_ _19132_/Q _19130_/Q _16767_/S vssd1 vssd1 vccd1 vccd1 _16768_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13979_ _13783_/X _13973_/X _13978_/X vssd1 vssd1 vccd1 vccd1 _13979_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03155_ _14312_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03155_/X sky130_fd_sc_hd__clkbuf_16
X_18506_ _18506_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18437_ _18437_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _15655_/A vssd1 vssd1 vccd1 vccd1 _15649_/X sky130_fd_sc_hd__buf_1
XFILLER_210_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09170_ _19171_/Q _09080_/X _09178_/S vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__mux2_1
X_18368_ _18368_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402__576 _14405__579/A vssd1 vssd1 vccd1 vccd1 _18211_/CLK sky130_fd_sc_hd__inv_2
XFILLER_175_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ _17357_/S vssd1 vssd1 vccd1 vccd1 _17333_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_159_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14814__744 _14814__744/A vssd1 vssd1 vccd1 vccd1 _18387_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18299_ _18299_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPeripherals_190 vssd1 vssd1 vccd1 vccd1 Peripherals_190/HI wb_data_o[29] sky130_fd_sc_hd__conb_1
Xclkbuf_0__03988_ _15785_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03988_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08954_ _08954_/A vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16325__223 _16326__224/A vssd1 vssd1 vccd1 vccd1 _18939_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08885_ _08885_/A vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09506_ _09506_/A vssd1 vssd1 vccd1 vccd1 _19005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ _14637_/A vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__clkbuf_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09368_ _09368_/A vssd1 vssd1 vccd1 vccd1 _19079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09299_ _19112_/Q _08967_/X _09299_/S vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11330_ _11329_/X _18144_/Q _11336_/S vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03144_ clkbuf_0__03144_/X vssd1 vssd1 vccd1 vccd1 _14260__463/A sky130_fd_sc_hd__clkbuf_16
X_15147__858 _15147__858/A vssd1 vssd1 vccd1 vccd1 _18534_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11261_ _11283_/S vssd1 vssd1 vccd1 vccd1 _11274_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_238_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13000_ _12992_/X _13000_/B vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__and2b_1
X_10212_ _10212_/A vssd1 vssd1 vccd1 vccd1 _18682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11192_ _18200_/Q _11050_/X _11196_/S vssd1 vssd1 vccd1 vccd1 _11193_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10143_ _18709_/Q _10054_/X _10149_/S vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _18460_/Q vssd1 vssd1 vccd1 vccd1 _15005_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10074_ _10074_/A vssd1 vssd1 vccd1 vccd1 _18735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13902_ _13908_/A vssd1 vssd1 vccd1 vccd1 _13902_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03977_ clkbuf_0__03977_/X vssd1 vssd1 vccd1 vccd1 _15729__1019/A sky130_fd_sc_hd__clkbuf_16
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17670_ _19037_/CLK _17670_/D vssd1 vssd1 vccd1 vccd1 _17670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16621_ _19039_/Q _16619_/B _16620_/Y vssd1 vssd1 vccd1 vccd1 _19039_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13833_ _17920_/Q _13829_/X _13832_/X _13826_/X vssd1 vssd1 vccd1 vccd1 _17920_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_206 _11818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19340_ _19340_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_217 _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13764_ _17898_/Q _13762_/X _13763_/Y vssd1 vssd1 vccd1 vccd1 _17898_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10976_ _10976_/A vssd1 vssd1 vccd1 vccd1 _18287_/D sky130_fd_sc_hd__clkbuf_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15503_ _17838_/Q _15517_/B vssd1 vssd1 vccd1 vccd1 _15511_/A sky130_fd_sc_hd__or2_1
X_12715_ _12717_/B _12713_/A _12695_/X vssd1 vssd1 vccd1 vccd1 _12716_/B sky130_fd_sc_hd__o21ai_1
X_19271_ _19271_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16483_ _16498_/A _16483_/B _16492_/C vssd1 vssd1 vccd1 vccd1 _16483_/X sky130_fd_sc_hd__or3_1
XFILLER_241_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13695_ _17875_/Q _13682_/X _13694_/Y vssd1 vssd1 vccd1 vccd1 _17875_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04529_ clkbuf_0__04529_/X vssd1 vssd1 vccd1 vccd1 _16555__264/A sky130_fd_sc_hd__clkbuf_16
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18222_ _18222_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12646_ _12647_/B _12647_/C _12645_/Y vssd1 vssd1 vccd1 vccd1 _17602_/D sky130_fd_sc_hd__o21a_1
XFILLER_176_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18153_ _18153_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15365_ _15359_/X _15364_/X _09620_/A vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__o21a_1
X_12577_ _12746_/B _12746_/A _17633_/Q _12758_/B _12555_/X _12556_/X vssd1 vssd1 vccd1
+ vccd1 _12577_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17104_ _17773_/Q _12187_/A _12121_/D vssd1 vssd1 vccd1 vccd1 _17104_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18084_ _19337_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11528_ _11528_/A vssd1 vssd1 vccd1 vccd1 _18032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15296_ _18938_/Q _18901_/Q _18893_/Q _18847_/Q _15251_/X _15252_/X vssd1 vssd1 vccd1
+ vccd1 _15296_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14247_ _16216_/A vssd1 vssd1 vccd1 vccd1 _14247_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11459_ _11321_/X _18063_/Q _11467_/S vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__08200_ clkbuf_0__08200_/X vssd1 vssd1 vccd1 vccd1 _13111__415/A sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14178_ _14256_/A vssd1 vssd1 vccd1 vccd1 _14178_/X sky130_fd_sc_hd__buf_1
XFILLER_140_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _18074_/Q _18075_/Q _13645_/A vssd1 vssd1 vccd1 vccd1 _13873_/D sky130_fd_sc_hd__or3_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _19013_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17049__39 _17049__39/A vssd1 vssd1 vccd1 vccd1 _19188_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17937_ _18024_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17868_ _18031_/CLK _17868_/D vssd1 vssd1 vccd1 vccd1 _17868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16819_ _16902_/A vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17799_ _19135_/CLK _17799_/D vssd1 vssd1 vccd1 vccd1 _17799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _09222_/A vssd1 vssd1 vccd1 vccd1 _19148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09153_ _09153_/A vssd1 vssd1 vccd1 vccd1 _19179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _09148_/B _19014_/Q _09084_/C vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__and3_1
XFILLER_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16546__257 _16548__259/A vssd1 vssd1 vccd1 vccd1 _19003_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09986_ _18770_/Q _09955_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__mux2_1
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08937_ _09694_/A vssd1 vssd1 vccd1 vccd1 _08937_/X sky130_fd_sc_hd__buf_2
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__buf_6
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08799_ _19343_/Q _08798_/X _08805_/S vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344__530 _14348__534/A vssd1 vssd1 vccd1 vccd1 _18165_/CLK sky130_fd_sc_hd__inv_2
X_10830_ _10830_/A vssd1 vssd1 vccd1 vccd1 _18356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10761_ _10761_/A vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _12727_/B _12727_/A _17627_/Q _17628_/Q _12555_/A _12429_/S vssd1 vssd1 vccd1
+ vccd1 _12500_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10692_ _10714_/S vssd1 vssd1 vccd1 vccd1 _10705_/S sky130_fd_sc_hd__clkbuf_2
X_13480_ _17807_/Q _16522_/A _13484_/S vssd1 vssd1 vccd1 vccd1 _13481_/B sky130_fd_sc_hd__mux2_1
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _12686_/B _17614_/Q _12440_/S vssd1 vssd1 vccd1 vccd1 _12431_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12362_ _17621_/Q vssd1 vssd1 vccd1 vccd1 _12717_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_194_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14101_ _18016_/Q _14091_/X _14100_/Y vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _11156_/X _18150_/Q _11313_/S vssd1 vssd1 vccd1 vccd1 _11314_/A sky130_fd_sc_hd__mux2_1
X_12293_ _17563_/Q _18014_/Q _12293_/S vssd1 vssd1 vccd1 vccd1 _12294_/B sky130_fd_sc_hd__mux2_1
X_15081_ _15081_/A vssd1 vssd1 vccd1 vccd1 _18482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14032_ _14039_/A vssd1 vssd1 vccd1 vccd1 _14032_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11244_ _11244_/A vssd1 vssd1 vccd1 vccd1 _18178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18840_ _18840_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_1
X_11175_ _11175_/A vssd1 vssd1 vccd1 vccd1 _18208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _10126_/A vssd1 vssd1 vccd1 vccd1 _10126_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18771_ _18771_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _15980_/Y _15981_/Y _15982_/X vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__a21oi_1
XFILLER_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _17953_/CLK _17722_/D vssd1 vssd1 vccd1 vccd1 _17722_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ _14934_/A _14934_/B vssd1 vssd1 vccd1 vccd1 _14935_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10057_ _10120_/A vssd1 vssd1 vccd1 vccd1 _10057_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04010_ clkbuf_0__04010_/X vssd1 vssd1 vccd1 vccd1 _15859__158/A sky130_fd_sc_hd__clkbuf_16
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _18006_/CLK _17653_/D vssd1 vssd1 vccd1 vccd1 _17653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16604_ _19031_/Q _16602_/B _14184_/A vssd1 vssd1 vccd1 vccd1 _16604_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13816_ _13815_/X _13802_/A _13805_/X vssd1 vssd1 vccd1 vccd1 _13816_/Y sky130_fd_sc_hd__a21oi_1
X_17584_ _17584_/CLK _17584_/D vssd1 vssd1 vccd1 vccd1 _17584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14796_ _14802_/A vssd1 vssd1 vccd1 vccd1 _14796_/X sky130_fd_sc_hd__buf_1
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19323_ _19323_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
X_16535_ _16534_/B _16507_/A _16534_/A _14619_/A vssd1 vssd1 vccd1 vccd1 _16536_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13747_ _17892_/Q _13738_/X _13746_/Y _13741_/X vssd1 vssd1 vccd1 vccd1 _17892_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10959_ _08877_/X _18294_/Q _10959_/S vssd1 vssd1 vccd1 vccd1 _10960_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19254_ _19261_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
X_15089__812 _15089__812/A vssd1 vssd1 vccd1 vccd1 _18488_/CLK sky130_fd_sc_hd__inv_2
X_16466_ _18976_/Q _16466_/B _16466_/C vssd1 vssd1 vccd1 vccd1 _16473_/B sky130_fd_sc_hd__and3_1
X_13678_ _17869_/Q _13660_/X _13677_/Y vssd1 vssd1 vccd1 vccd1 _17869_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18205_ _18205_/CLK _18205_/D vssd1 vssd1 vccd1 vccd1 _18205_/Q sky130_fd_sc_hd__dfxtp_1
X_15427__923 _15428__924/A vssd1 vssd1 vccd1 vccd1 _18610_/CLK sky130_fd_sc_hd__inv_2
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15417_ _15441_/A vssd1 vssd1 vccd1 vccd1 _15417_/X sky130_fd_sc_hd__buf_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ _17598_/Q _17597_/Q vssd1 vssd1 vccd1 vccd1 _12630_/D sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__04843_ clkbuf_0__04843_/X vssd1 vssd1 vccd1 vccd1 _17042__34/A sky130_fd_sc_hd__clkbuf_16
X_19185_ _19185_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
X_16397_ _18974_/Q _16397_/B _16397_/C vssd1 vssd1 vccd1 vccd1 _16418_/A sky130_fd_sc_hd__and3_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_38_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19281_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18136_ _18136_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15348_ _15342_/X _15347_/X _09620_/A vssd1 vssd1 vccd1 vccd1 _15348_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18067_ _19146_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15279_ _15279_/A _15307_/A vssd1 vssd1 vccd1 vccd1 _15279_/X sky130_fd_sc_hd__or2b_1
XFILLER_208_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14514__666 _14514__666/A vssd1 vssd1 vccd1 vccd1 _18301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_171_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ _09694_/X _18813_/Q _09842_/S vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03587_ clkbuf_0__03587_/X vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _11529_/B _11601_/B vssd1 vssd1 vccd1 vccd1 _09787_/S sky130_fd_sc_hd__or2_2
X_15096__816 _15099__819/A vssd1 vssd1 vccd1 vccd1 _18492_/CLK sky130_fd_sc_hd__inv_2
X_18969_ _18971_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16552__261 _16552__261/A vssd1 vssd1 vccd1 vccd1 _19007_/CLK sky130_fd_sc_hd__inv_2
X_09205_ _10691_/B hold8/A vssd1 vssd1 vccd1 vccd1 _09221_/S sky130_fd_sc_hd__nor2_2
XFILLER_167_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _18664_/Q vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09067_ _19201_/Q _08871_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16071__187 _16071__187/A vssd1 vssd1 vccd1 vccd1 _18892_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09969_ _09969_/A vssd1 vssd1 vccd1 vccd1 _18775_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12980_ _17958_/Q _17679_/Q _12993_/S vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__mux2_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _19222_/Q _17129_/B _11931_/S vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__mux2_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _19078_/Q _18342_/Q _17576_/Q _18794_/Q _14575_/X _09459_/X vssd1 vssd1 vccd1
+ vccd1 _14651_/B sky130_fd_sc_hd__mux4_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _13820_/A _11865_/B _11862_/C vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__and3_1
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13601_ _13621_/B vssd1 vssd1 vccd1 vccd1 _13601_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10813_ _18363_/Q _10812_/X _10813_/S vssd1 vssd1 vccd1 vccd1 _10814_/A sky130_fd_sc_hd__mux2_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14581_ _18585_/Q _18299_/Q _17565_/Q _18836_/Q _14579_/X _14580_/X vssd1 vssd1 vccd1
+ vccd1 _14581_/X sky130_fd_sc_hd__mux4_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11793_ _11812_/A vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13532_ _13689_/A vssd1 vssd1 vccd1 vccd1 _13532_/X sky130_fd_sc_hd__buf_2
XFILLER_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _18390_/Q _10704_/X _10744_/S vssd1 vssd1 vccd1 vccd1 _10745_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16251_ _16249_/X _16250_/X _16289_/S vssd1 vssd1 vccd1 vccd1 _16251_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _17802_/Q _13463_/B vssd1 vssd1 vccd1 vccd1 _13463_/Y sky130_fd_sc_hd__nor2_1
X_10675_ _10675_/A vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12414_ _17617_/Q vssd1 vssd1 vccd1 vccd1 _12707_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16182_ _16182_/A vssd1 vssd1 vccd1 vccd1 _16182_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13394_ _14072_/A vssd1 vssd1 vccd1 vccd1 _13394_/X sky130_fd_sc_hd__buf_4
XFILLER_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12345_ _13103_/A vssd1 vssd1 vccd1 vccd1 _12345_/X sky130_fd_sc_hd__buf_1
X_15876__171 _15878__173/A vssd1 vssd1 vccd1 vccd1 _18846_/CLK sky130_fd_sc_hd__inv_2
XFILLER_154_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04590_ _16719_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04590_/X sky130_fd_sc_hd__clkbuf_16
X_15064_ _15064_/A _15174_/B _16052_/C vssd1 vssd1 vccd1 vccd1 _15177_/A sky130_fd_sc_hd__nand3_4
X_12276_ _12276_/A vssd1 vssd1 vccd1 vccd1 _17557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14015_ _13719_/A _14012_/X _14005_/X vssd1 vssd1 vccd1 vccd1 _14015_/Y sky130_fd_sc_hd__a21oi_1
X_11227_ _11147_/X _18185_/Q _11233_/S vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18823_ _18823_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11158_ _11158_/A vssd1 vssd1 vccd1 vccd1 _18214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10109_ _10109_/A vssd1 vssd1 vccd1 vccd1 _18720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18754_ _18754_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_1
X_11089_ _11104_/S vssd1 vssd1 vccd1 vccd1 _11098_/S sky130_fd_sc_hd__clkbuf_2
X_15966_ _16033_/A _15966_/B vssd1 vssd1 vccd1 vccd1 _18862_/D sky130_fd_sc_hd__nor2_1
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14917_ _18464_/Q _14917_/B vssd1 vssd1 vccd1 vccd1 _14963_/C sky130_fd_sc_hd__xor2_1
X_17705_ _17705_/CLK _17705_/D vssd1 vssd1 vccd1 vccd1 _17705_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ _17825_/Q _17824_/Q _17823_/Q _17822_/Q vssd1 vssd1 vccd1 vccd1 _15932_/B
+ sky130_fd_sc_hd__or4_2
X_18685_ _18685_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17636_ _19247_/CLK _17636_/D vssd1 vssd1 vccd1 vccd1 _17636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17042__34 _17042__34/A vssd1 vssd1 vccd1 vccd1 _19183_/CLK sky130_fd_sc_hd__inv_2
X_17567_ _17567_/CLK _17567_/D vssd1 vssd1 vccd1 vccd1 _17567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19306_ _19306_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
X_16518_ input55/X _16518_/B _16530_/B vssd1 vssd1 vccd1 vccd1 _16519_/A sky130_fd_sc_hd__and3_1
XFILLER_182_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17498_ _17498_/A vssd1 vssd1 vccd1 vccd1 _19340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19237_ _19248_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16449_ _16453_/B _16453_/C vssd1 vssd1 vccd1 vccd1 _16449_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19168_ _19168_/CLK _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18119_ _18119_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_1
X_19099_ _19099_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03808_ _15455_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03808_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104__823 _15105__824/A vssd1 vssd1 vccd1 vccd1 _18499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09823_ _09823_/A vssd1 vssd1 vccd1 vccd1 _18821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _09754_/A vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ _09685_/A vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14148__432 _14149__433/A vssd1 vssd1 vccd1 vccd1 _18040_/CLK sky130_fd_sc_hd__inv_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10460_ _18546_/Q _10333_/X _10466_/S vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ _18668_/Q vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__buf_2
XFILLER_182_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10391_ _16291_/A vssd1 vssd1 vccd1 vccd1 _10391_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__04013_ clkbuf_0__04013_/X vssd1 vssd1 vccd1 vccd1 _15872__168/A sky130_fd_sc_hd__clkbuf_16
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _11888_/X _12130_/B vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__and2b_1
XFILLER_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12061_ _12018_/X _12051_/X _12060_/X _12045_/S vssd1 vssd1 vccd1 vccd1 _12061_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11012_ _09035_/X _18272_/Q _11016_/S vssd1 vssd1 vccd1 vccd1 _11013_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15820_ _18889_/Q _15812_/Y _16064_/A _15819_/X vssd1 vssd1 vccd1 vccd1 _18801_/D
+ sky130_fd_sc_hd__o211a_4
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04846_ clkbuf_0__04846_/X vssd1 vssd1 vccd1 vccd1 _17055__44/A sky130_fd_sc_hd__clkbuf_16
XFILLER_218_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _12957_/X _12963_/B vssd1 vssd1 vccd1 vccd1 _12964_/A sky130_fd_sc_hd__and2b_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_60 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_71 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_82 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14702_ _14664_/A _14701_/X _14619_/X vssd1 vssd1 vccd1 vccd1 _14702_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_93 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ _19244_/Q vssd1 vssd1 vccd1 vccd1 _17209_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18470_ _18921_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12894_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12894_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__buf_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14633_ _19150_/Q _18415_/Q _18309_/Q _18293_/Q _09443_/A _14575_/X vssd1 vssd1 vccd1
+ vccd1 _14634_/B sky130_fd_sc_hd__mux4_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11848_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__and2_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17352_ _17352_/A vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14575_/A vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _18081_/Q vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__inv_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03990_ clkbuf_0__03990_/X vssd1 vssd1 vccd1 vccd1 _15788__110/A sky130_fd_sc_hd__clkbuf_16
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16303_ _18327_/Q _18328_/Q _18329_/Q _18330_/Q _18984_/Q _18985_/Q vssd1 vssd1 vccd1
+ vccd1 _16303_/X sky130_fd_sc_hd__mux4_1
X_13515_ _17816_/Q _13499_/X _13514_/Y vssd1 vssd1 vccd1 vccd1 _17816_/D sky130_fd_sc_hd__o21a_1
X_17283_ _17279_/A _17288_/D _17288_/B vssd1 vssd1 vccd1 vccd1 _17285_/B sky130_fd_sc_hd__a21o_1
X_10727_ _10727_/A vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__clkbuf_1
X_19022_ _19027_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _16234_/A _16234_/B vssd1 vssd1 vccd1 vccd1 _16234_/Y sky130_fd_sc_hd__nand2_1
X_13446_ input58/X _13446_/B vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__and2_4
XFILLER_174_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10658_ _18427_/Q _09723_/X _10662_/S vssd1 vssd1 vccd1 vccd1 _10659_/A sky130_fd_sc_hd__mux2_1
X_14357__540 _14358__541/A vssd1 vssd1 vccd1 vccd1 _18175_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16165_ _10391_/X _16147_/X _16163_/Y _16164_/X vssd1 vssd1 vccd1 vccd1 _16165_/Y
+ sky130_fd_sc_hd__o211ai_1
X_13377_ _12017_/S _13355_/X _13375_/Y _13376_/X vssd1 vssd1 vccd1 vccd1 _17780_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10589_ _10589_/A vssd1 vssd1 vccd1 vccd1 _18490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15047_ _15047_/A vssd1 vssd1 vccd1 vccd1 _18467_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__04573_ _16652_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04573_/X sky130_fd_sc_hd__clkbuf_16
X_12259_ _17553_/Q _18024_/Q _12270_/S vssd1 vssd1 vccd1 vccd1 _12260_/B sky130_fd_sc_hd__mux2_1
XFILLER_218_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03424_ clkbuf_0__03424_/X vssd1 vssd1 vccd1 vccd1 _15085__809/A sky130_fd_sc_hd__clkbuf_16
XFILLER_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17410__100 _17412__102/A vssd1 vssd1 vccd1 vccd1 _19313_/CLK sky130_fd_sc_hd__inv_2
XFILLER_228_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18806_ _18806_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16998_ _16998_/A vssd1 vssd1 vccd1 vccd1 _19147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18737_ _18737_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15949_ _18875_/Q vssd1 vssd1 vccd1 vccd1 _15949_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09470_ _10670_/S vssd1 vssd1 vccd1 vccd1 _10662_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18668_ _14157_/A _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17619_ _17621_/CLK _17619_/D vssd1 vssd1 vccd1 vccd1 _17619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17011__359 _17011__359/A vssd1 vssd1 vccd1 vccd1 _19158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18599_ _18599_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__04007_ _15837_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04007_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_225_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18012_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_196_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__07559_ _12339_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07559_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_160_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14863__784 _14863__784/A vssd1 vssd1 vccd1 vccd1 _18429_/CLK sky130_fd_sc_hd__inv_2
X_09806_ _18828_/Q _09767_/X _09806_/S vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ _09737_/A vssd1 vssd1 vccd1 vccd1 _18855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09668_ _18908_/Q _09274_/X _09672_/S vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827__132 _15829__134/A vssd1 vssd1 vccd1 vccd1 _18807_/CLK sky130_fd_sc_hd__inv_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09599_ _18934_/Q vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11630_/A vssd1 vssd1 vccd1 vccd1 _17543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14161__440 _14162__441/A vssd1 vssd1 vccd1 vccd1 _18048_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _17705_/Q _10907_/X _11563_/S vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13300_ _13247_/X _13288_/A _13293_/X vssd1 vssd1 vccd1 vccd1 _13300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_195_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10512_ _18523_/Q _10328_/X _10520_/S vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11492_ _11492_/A vssd1 vssd1 vccd1 vccd1 _18048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13231_ _13777_/A vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__buf_4
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10443_ _10443_/A vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13162_ _17727_/Q _14134_/B vssd1 vssd1 vccd1 vccd1 _13162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10374_ _08724_/X _18584_/Q _10382_/S vssd1 vssd1 vccd1 vccd1 _10375_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ _12113_/A vssd1 vssd1 vccd1 vccd1 _12113_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_151_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17970_ _19016_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
X_13093_ _17696_/Q _13093_/B vssd1 vssd1 vccd1 vccd1 _13096_/B sky130_fd_sc_hd__xnor2_1
XFILLER_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12045_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16921_ _18060_/Q _18052_/Q _18044_/Q _18036_/Q _16870_/X _16871_/X vssd1 vssd1 vccd1
+ vccd1 _16921_/X sky130_fd_sc_hd__mux4_2
XFILLER_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16852_ _16986_/A _16852_/B vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16783_ _16783_/A _16783_/B vssd1 vssd1 vccd1 vccd1 _16783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13995_ _13995_/A vssd1 vssd1 vccd1 vccd1 _13995_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18522_ _18522_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03171_ _14388_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03171_/X sky130_fd_sc_hd__clkbuf_16
X_12946_ _18001_/Q _13024_/B vssd1 vssd1 vccd1 vccd1 _12999_/S sky130_fd_sc_hd__and2_2
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18453_ _18921_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12877_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _18586_/Q _18300_/Q _17566_/Q _18837_/Q _14615_/X _09459_/X vssd1 vssd1 vccd1
+ vccd1 _14616_/X sky130_fd_sc_hd__mux4_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _14053_/A vssd1 vssd1 vccd1 vccd1 _13279_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18384_ _18384_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15596_ _15611_/A _15596_/B _15605_/C vssd1 vssd1 vccd1 vccd1 _15596_/X sky130_fd_sc_hd__or3_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17335_/A vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _19172_/Q _19164_/Q _19196_/Q _18331_/Q _14641_/A _14546_/X vssd1 vssd1 vccd1
+ vccd1 _14547_/X sky130_fd_sc_hd__mux4_1
X_11759_ _11759_/A vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_230_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03973_ clkbuf_0__03973_/X vssd1 vssd1 vccd1 vccd1 _15707__1001/A sky130_fd_sc_hd__clkbuf_16
XFILLER_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17266_ _17266_/A vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16217_ _18917_/Q _16098_/X _16215_/Y _16216_/X vssd1 vssd1 vccd1 vccd1 _18917_/D
+ sky130_fd_sc_hd__o211a_1
X_19005_ _19005_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13429_ _16736_/A vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__buf_4
X_17197_ _17194_/B _17195_/A _19241_/Q vssd1 vssd1 vccd1 vccd1 _17198_/C sky130_fd_sc_hd__a21o_1
XFILLER_220_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ _18744_/Q _18752_/Q _18760_/Q _18768_/Q _16127_/X _16128_/X vssd1 vssd1 vccd1
+ vccd1 _16148_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08970_ _09789_/B vssd1 vssd1 vccd1 vccd1 _09639_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_100_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19013_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03407_ clkbuf_0__03407_/X vssd1 vssd1 vccd1 vccd1 _14807__739/A sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 flash_csb vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_244_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09522_ _18998_/Q _09501_/X _09524_/S vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09453_ _09477_/C _09453_/B _09453_/C vssd1 vssd1 vccd1 vccd1 _09454_/A sky130_fd_sc_hd__and3_1
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ _19072_/Q _08952_/X _09388_/S vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03160_ clkbuf_0__03160_/X vssd1 vssd1 vccd1 vccd1 _14342__529/A sky130_fd_sc_hd__clkbuf_16
XFILLER_123_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03091_ clkbuf_0__03091_/X vssd1 vssd1 vccd1 vccd1 _14155__438/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17417__106 _17419__108/A vssd1 vssd1 vccd1 vccd1 _19319_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10090_ _18728_/Q _10069_/X _10092_/S vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03993_ clkbuf_0__03993_/X vssd1 vssd1 vccd1 vccd1 _15807__126/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12800_ _12795_/X _12800_/B vssd1 vssd1 vccd1 vccd1 _12801_/A sky130_fd_sc_hd__and2b_1
XFILLER_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308__501 _14310__503/A vssd1 vssd1 vccd1 vccd1 _18136_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ _17903_/Q _13770_/X _13779_/Y vssd1 vssd1 vccd1 vccd1 _17903_/D sky130_fd_sc_hd__o21a_1
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10992_ _18281_/Q _09127_/X _10998_/S vssd1 vssd1 vccd1 vccd1 _10993_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12731_ _12737_/C _12737_/D _12718_/X vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__o21ai_1
XFILLER_215_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12662_ _17607_/Q _12666_/C _12666_/D vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__and3_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _17567_/Q _10707_/A _11617_/S vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__mux2_1
X_15381_ _15307_/X _15377_/X _15380_/Y vssd1 vssd1 vccd1 vccd1 _15381_/X sky130_fd_sc_hd__o21a_2
X_12593_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _17782_/Q _19222_/Q _19221_/Q _19220_/Q vssd1 vssd1 vccd1 vccd1 _17133_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11544_ _11544_/A vssd1 vssd1 vccd1 vccd1 _17713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14263_/X sky130_fd_sc_hd__buf_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11475_ _11475_/A hold23/X vssd1 vssd1 vccd1 vccd1 _11491_/S sky130_fd_sc_hd__or2_2
XFILLER_137_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15421__918 _15422__919/A vssd1 vssd1 vccd1 vccd1 _18605_/CLK sky130_fd_sc_hd__inv_2
X_16002_ _18869_/Q _16002_/B _16002_/C vssd1 vssd1 vccd1 vccd1 _16007_/B sky130_fd_sc_hd__and3_1
X_13214_ _13180_/B _16054_/A _13212_/Y _13213_/X vssd1 vssd1 vccd1 vccd1 _17736_/D
+ sky130_fd_sc_hd__a211oi_1
X_10426_ _09975_/C _10424_/X _10425_/Y vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__o21a_1
X_14194_ _18069_/Q input49/X _14196_/S vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ input58/X _13431_/B vssd1 vssd1 vccd1 vccd1 _13724_/A sky130_fd_sc_hd__nand2_4
XFILLER_125_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10357_ _10357_/A vssd1 vssd1 vccd1 vccd1 _18592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _17936_/Q _17702_/Q _13076_/S vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__mux2_1
X_17953_ _17953_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14469__630 _14473__634/A vssd1 vssd1 vccd1 vccd1 _18265_/CLK sky130_fd_sc_hd__inv_2
X_10288_ _18618_/Q _10195_/X _10290_/S vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12027_ _19259_/Q vssd1 vssd1 vccd1 vccd1 _17264_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16904_ _18246_/Q _18238_/Q _18230_/Q _18222_/Q _16849_/X _16850_/X vssd1 vssd1 vccd1
+ vccd1 _16905_/B sky130_fd_sc_hd__mux4_2
XFILLER_238_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17884_ _18021_/CLK _17884_/D vssd1 vssd1 vccd1 vccd1 _17884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16835_ _18211_/Q _18195_/Q _18484_/Q _18187_/Q _16834_/X _09875_/X vssd1 vssd1 vccd1
+ vccd1 _16835_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14168__446 _14168__446/A vssd1 vssd1 vccd1 vccd1 _18054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13978_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__clkbuf_2
X_16766_ _19131_/Q _16771_/B vssd1 vssd1 vccd1 vccd1 _16766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03154_ _14306_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03154_/X sky130_fd_sc_hd__clkbuf_16
X_18505_ _18505_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_1
X_12929_ _17663_/Q _13085_/B vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15717_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15717_/X sky130_fd_sc_hd__buf_1
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18436_ _18436_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ _15579_/A _15579_/B _15584_/B vssd1 vssd1 vccd1 vccd1 _15579_/X sky130_fd_sc_hd__or3_1
X_18367_ _18367_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17318_ _17318_/A vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _18298_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17249_ _17249_/A vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__clkbuf_1
XPeripherals_180 vssd1 vssd1 vccd1 vccd1 Peripherals_180/HI wb_data_o[19] sky130_fd_sc_hd__conb_1
XFILLER_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03987_ _15779_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03987_/X sky130_fd_sc_hd__clkbuf_16
XPeripherals_191 vssd1 vssd1 vccd1 vccd1 Peripherals_191/HI wb_data_o[30] sky130_fd_sc_hd__conb_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08953_ _19272_/Q _08952_/X _08959_/S vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08884_ _19309_/Q _08883_/X _08887_/S vssd1 vssd1 vccd1 vccd1 _08885_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09505_ _19005_/Q _09504_/X _09505_/S vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14637_/A sky130_fd_sc_hd__clkbuf_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _19079_/Q _09100_/X _09369_/S vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303__497 _14305__499/A vssd1 vssd1 vccd1 vccd1 _18132_/CLK sky130_fd_sc_hd__inv_2
X_09298_ _09298_/A vssd1 vssd1 vccd1 vccd1 _19113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11260_ _11260_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11283_/S sky130_fd_sc_hd__nor2_2
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10211_ _18682_/Q _09758_/X _10211_/S vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11191_ _11191_/A vssd1 vssd1 vccd1 vccd1 _18201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10142_ _10142_/A vssd1 vssd1 vccd1 vccd1 _18710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15870__166 _15872__168/A vssd1 vssd1 vccd1 vccd1 _18841_/CLK sky130_fd_sc_hd__inv_2
XFILLER_239_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _14950_/A _14950_/B _14950_/C _14950_/D vssd1 vssd1 vccd1 vccd1 _14961_/C
+ sky130_fd_sc_hd__or4_1
X_10073_ _18735_/Q _10072_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__mux2_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03976_ clkbuf_0__03976_/X vssd1 vssd1 vccd1 vccd1 _15748_/A sky130_fd_sc_hd__clkbuf_16
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _14031_/A _16516_/D _14076_/C vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__and3_1
XFILLER_248_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16620_ _16620_/A _16620_/B vssd1 vssd1 vccd1 vccd1 _16620_/Y sky130_fd_sc_hd__nor2_1
X_13832_ input61/X _13845_/B vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__and2_1
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_207 _11820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13763_ _13707_/A _13762_/X _13701_/X vssd1 vssd1 vccd1 vccd1 _13763_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_218 _18885_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10975_ _18287_/Q _09755_/X _10977_/S vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12717_/B _12717_/C _12717_/D vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__and3_1
XFILLER_243_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15502_ _18649_/Q _15502_/B vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__xor2_1
X_19270_ _19270_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
X_16482_ _18979_/Q _18978_/Q _16482_/C vssd1 vssd1 vccd1 vccd1 _16492_/C sky130_fd_sc_hd__and3_1
XFILLER_245_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13694_ _13411_/X _13688_/X _13689_/X vssd1 vssd1 vccd1 vccd1 _13694_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14876__794 _14876__794/A vssd1 vssd1 vccd1 vccd1 _18439_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__04528_ clkbuf_0__04528_/X vssd1 vssd1 vccd1 vccd1 _16639_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18221_ _18221_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
X_12645_ _12647_/B _12647_/C _12755_/A vssd1 vssd1 vccd1 vccd1 _12645_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15364_ _15307_/X _15360_/X _15363_/Y vssd1 vssd1 vccd1 vccd1 _15364_/X sky130_fd_sc_hd__o21a_2
X_18152_ _18152_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_1
X_12576_ _17634_/Q vssd1 vssd1 vccd1 vccd1 _12758_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17103_ _13361_/X _17101_/X _12185_/X vssd1 vssd1 vccd1 vccd1 _17103_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18083_ _19337_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
X_11527_ _18032_/Q _11344_/A hold24/X vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15295_ _19000_/Q _18962_/Q _18954_/Q _17543_/Q _15273_/X _15249_/X vssd1 vssd1 vccd1
+ vccd1 _15295_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14246_ _15080_/B vssd1 vssd1 vccd1 vccd1 _16216_/A sky130_fd_sc_hd__clkbuf_2
X_11458_ _11473_/S vssd1 vssd1 vccd1 vccd1 _11467_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10409_ _10391_/X _10406_/X _10408_/Y vssd1 vssd1 vccd1 vccd1 _18568_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17526_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ _11389_/A vssd1 vssd1 vccd1 vccd1 _18121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13128_/A _11779_/A vssd1 vssd1 vccd1 vccd1 _13645_/A sky130_fd_sc_hd__or2b_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _18996_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _18024_/CLK _17936_/D vssd1 vssd1 vccd1 vccd1 _17936_/Q sky130_fd_sc_hd__dfxtp_1
X_13059_ _13059_/A vssd1 vssd1 vccd1 vccd1 _17696_/D sky130_fd_sc_hd__clkbuf_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17867_ _18031_/CLK _17867_/D vssd1 vssd1 vccd1 vccd1 _17867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16818_ _18811_/Q vssd1 vssd1 vccd1 vccd1 _16818_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17798_ _19135_/CLK _17798_/D vssd1 vssd1 vccd1 vccd1 _17798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16749_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16749_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09221_ _19148_/Q _09116_/X _09221_/S vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__mux2_1
X_14142__427 _14144__429/A vssd1 vssd1 vccd1 vccd1 _18035_/CLK sky130_fd_sc_hd__inv_2
X_18419_ _18419_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19399_ input20/X vssd1 vssd1 vccd1 vccd1 _19399_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _19179_/Q _09080_/X _09160_/S vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09083_ _08728_/X _08857_/X _11675_/A vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__a21o_4
XFILLER_238_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput70 wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_4
XFILLER_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09985_ _09985_/A vssd1 vssd1 vccd1 vccd1 _18771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17296__73 _17296__73/A vssd1 vssd1 vccd1 vccd1 _19269_/CLK sky130_fd_sc_hd__inv_2
X_08936_ _18881_/Q vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__buf_2
XFILLER_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ _08867_/A vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _18882_/Q vssd1 vssd1 vccd1 vccd1 _08798_/X sky130_fd_sc_hd__buf_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19146_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153__863 _15153__863/A vssd1 vssd1 vccd1 vccd1 _18539_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10760_ _18383_/Q _10701_/X _10762_/S vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _09419_/A vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10691_ _11529_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _10714_/S sky130_fd_sc_hd__nor2_2
XFILLER_240_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ _17613_/Q vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _17620_/Q vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ _13777_/A _14099_/X _14096_/X vssd1 vssd1 vccd1 vccd1 _14100_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_181_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11312_/A vssd1 vssd1 vccd1 vccd1 _18151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15080_ _15079_/Y _15080_/B _15080_/C vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__and3b_1
X_12292_ _12292_/A vssd1 vssd1 vccd1 vccd1 _17562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ _14031_/A _14031_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _14039_/A sky130_fd_sc_hd__and3_2
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11243_ _11142_/X _18178_/Q _11251_/S vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14763__703 _14763__703/A vssd1 vssd1 vccd1 vccd1 _18346_/CLK sky130_fd_sc_hd__inv_2
X_11174_ _11150_/X _18208_/Q _11178_/S vssd1 vssd1 vccd1 vccd1 _11175_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10125_ _10125_/A vssd1 vssd1 vccd1 vccd1 _18715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18770_ _18770_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _16010_/A vssd1 vssd1 vccd1 vccd1 _15982_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _18465_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _17721_/Q sky130_fd_sc_hd__dfxtp_4
X_15201__886 _15203__888/A vssd1 vssd1 vccd1 vccd1 _18565_/CLK sky130_fd_sc_hd__inv_2
X_14933_ _17851_/Q _14938_/A vssd1 vssd1 vccd1 vccd1 _14934_/B sky130_fd_sc_hd__and2_1
X_10056_ _10056_/A vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16675__309 _16675__309/A vssd1 vssd1 vccd1 vccd1 _19083_/CLK sky130_fd_sc_hd__inv_2
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17652_ _17991_/CLK _17652_/D vssd1 vssd1 vccd1 vccd1 _17652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14864_ _14864_/A vssd1 vssd1 vccd1 vccd1 _14864_/X sky130_fd_sc_hd__buf_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _19030_/Q _16601_/B _16602_/Y vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__o21a_1
X_17054__43 _17055__44/A vssd1 vssd1 vccd1 vccd1 _19192_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13815_ _13815_/A vssd1 vssd1 vccd1 vccd1 _13815_/X sky130_fd_sc_hd__buf_4
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17583_ _17583_/CLK _17583_/D vssd1 vssd1 vccd1 vccd1 _17583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19322_ _19322_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
X_13746_ _13746_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13746_/Y sky130_fd_sc_hd__nor2_1
X_16534_ _16534_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _16534_/X sky130_fd_sc_hd__and2_1
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ _10958_/A vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19253_ _19261_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13677_ _13244_/X _13666_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _13677_/Y sky130_fd_sc_hd__a21oi_1
X_16465_ _16466_/B _16466_/C _18976_/Q vssd1 vssd1 vccd1 vccd1 _16467_/B sky130_fd_sc_hd__a21oi_1
X_10889_ _10911_/S vssd1 vssd1 vccd1 vccd1 _10902_/S sky130_fd_sc_hd__buf_2
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ _18204_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ _12631_/B _12628_/B vssd1 vssd1 vccd1 vccd1 _17597_/D sky130_fd_sc_hd__nor2_1
X_15416_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15416_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1__f__04842_ clkbuf_0__04842_/X vssd1 vssd1 vccd1 vccd1 _17033__26/A sky130_fd_sc_hd__clkbuf_16
X_19184_ _19184_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
X_16396_ _17804_/Q _17803_/Q _16412_/B _17802_/Q vssd1 vssd1 vccd1 vccd1 _16397_/C
+ sky130_fd_sc_hd__o31ai_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ _15307_/X _15343_/X _15346_/Y vssd1 vssd1 vccd1 vccd1 _15347_/X sky130_fd_sc_hd__o21a_2
X_18135_ _18135_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
X_12559_ _12493_/X _12494_/X _12485_/X _12486_/X _12449_/S _12568_/A vssd1 vssd1 vccd1
+ vccd1 _12559_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15278_ _18673_/Q _18579_/Q _17534_/Q _17509_/Q _15262_/X _09631_/A vssd1 vssd1 vccd1
+ vccd1 _15279_/A sky130_fd_sc_hd__mux4_1
X_18066_ _18870_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_1__f__07492_ clkbuf_0__07492_/X vssd1 vssd1 vccd1 vccd1 _12319__384/A sky130_fd_sc_hd__clkbuf_16
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14229_ _18085_/Q input43/X _14229_/S vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_78_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17609_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03586_ clkbuf_0__03586_/X vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_99_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09770_ _09770_/A _09770_/B _09358_/B vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__or3b_4
XFILLER_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18968_ _18971_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17919_ _17923_/CLK _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18899_ _18899_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15821__127 _15823__129/A vssd1 vssd1 vccd1 vccd1 _18802_/CLK sky130_fd_sc_hd__inv_2
X_09204_ _09770_/A _09358_/B hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__or3b_4
XFILLER_22_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09135_ _09135_/A vssd1 vssd1 vccd1 vccd1 _19184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09066_ _09066_/A vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415__587 _14417__589/A vssd1 vssd1 vccd1 vccd1 _18222_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09968_ _18775_/Q _09967_/X _09968_/S vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15789__111 _15792__114/A vssd1 vssd1 vccd1 vccd1 _18783_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _08919_/A vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09899_ _18798_/Q _09718_/X _09907_/S vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _11980_/A vssd1 vssd1 vccd1 vccd1 _11931_/S sky130_fd_sc_hd__buf_2
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11861_ _17918_/Q _11802_/A _11812_/A _17899_/Q vssd1 vssd1 vccd1 vccd1 _11862_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13611_/S vssd1 vssd1 vccd1 vccd1 _13621_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10812_ _18987_/Q vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__buf_2
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14580_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _11840_/A vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__buf_2
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13531_ _17821_/Q _13522_/X _13530_/Y vssd1 vssd1 vccd1 vccd1 _17821_/D sky130_fd_sc_hd__o21a_1
X_16338__234 _16338__234/A vssd1 vssd1 vccd1 vccd1 _18950_/CLK sky130_fd_sc_hd__inv_2
X_10743_ _10743_/A vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16250_ _18780_/Q _18638_/Q _18788_/Q _18622_/Q _16158_/X _16182_/X vssd1 vssd1 vccd1
+ vccd1 _16250_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13462_ _13477_/B vssd1 vssd1 vccd1 vccd1 _13463_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ _18420_/Q _09718_/X _10682_/S vssd1 vssd1 vccd1 vccd1 _10675_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12413_ _12773_/B vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__buf_2
XFILLER_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16181_ _18627_/Q _18502_/Q _18908_/Q _18510_/Q _16155_/X _16156_/X vssd1 vssd1 vccd1
+ vccd1 _16181_/X sky130_fd_sc_hd__mux4_1
X_13393_ _13395_/A vssd1 vssd1 vccd1 vccd1 _13393_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16681__313 _16682__314/A vssd1 vssd1 vccd1 vccd1 _19087_/CLK sky130_fd_sc_hd__inv_2
XFILLER_153_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15062_/Y _15060_/Y _14894_/Y vssd1 vssd1 vccd1 vccd1 _18472_/D sky130_fd_sc_hd__a21boi_1
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12275_ _12263_/X _12275_/B vssd1 vssd1 vccd1 vccd1 _12276_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14014_ _17984_/Q _14011_/X _14013_/Y vssd1 vssd1 vccd1 vccd1 _17984_/D sky130_fd_sc_hd__o21a_1
XFILLER_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _11226_/A vssd1 vssd1 vccd1 vccd1 _18186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18822_ _18822_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_1
X_11157_ _11156_/X _18214_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16345__238 _16346__239/A vssd1 vssd1 vccd1 vccd1 _18954_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10108_ _18720_/Q _10069_/X _10110_/S vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18753_ _18753_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11088_ _11475_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11104_/S sky130_fd_sc_hd__or2_2
X_15965_ _18862_/Q _16025_/B _15963_/X _15964_/Y vssd1 vssd1 vccd1 vccd1 _15966_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17704_ _17704_/CLK _17704_/D vssd1 vssd1 vccd1 vccd1 _17704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14916_ _14936_/A _14916_/B vssd1 vssd1 vccd1 vccd1 _14917_/B sky130_fd_sc_hd__nand2_1
X_10039_ _10039_/A vssd1 vssd1 vccd1 vccd1 _18747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17027__21 _17028__22/A vssd1 vssd1 vccd1 vccd1 _19170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18684_ _18684_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _16010_/A vssd1 vssd1 vccd1 vccd1 _16033_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17635_ _18012_/CLK _17635_/D vssd1 vssd1 vccd1 vccd1 _17635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15687__985 _15691__989/A vssd1 vssd1 vccd1 vccd1 _18702_/CLK sky130_fd_sc_hd__inv_2
XFILLER_223_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17566_ _17566_/CLK _17566_/D vssd1 vssd1 vccd1 vccd1 _17566_/Q sky130_fd_sc_hd__dfxtp_1
X_14778_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__buf_1
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19305_ _19305_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16517_ _16532_/C vssd1 vssd1 vccd1 vccd1 _16530_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_232_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13729_ _17886_/Q _13715_/X _13728_/Y _13726_/X vssd1 vssd1 vccd1 vccd1 _17886_/D
+ sky130_fd_sc_hd__a211o_1
X_17497_ _11888_/X _17497_/B _17497_/C vssd1 vssd1 vccd1 vccd1 _17498_/A sky130_fd_sc_hd__and3b_1
X_14520__671 _14520__671/A vssd1 vssd1 vccd1 vccd1 _18306_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19236_ _19248_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16448_ _16446_/X _16447_/Y _16480_/A vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__a21oi_1
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19167_ _19167_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
X_16379_ _18981_/Q _16379_/B vssd1 vssd1 vccd1 vccd1 _16379_/X sky130_fd_sc_hd__xor2_1
XFILLER_118_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18118_ _18118_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098_ _19098_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12323__387 _12325__389/A vssd1 vssd1 vccd1 vccd1 _17568_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03807_ _15449_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03807_/X sky130_fd_sc_hd__clkbuf_16
X_18049_ _18049_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09822_ _09694_/X _18821_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09753_ _18849_/Q _09752_/X _09759_/S vssd1 vssd1 vccd1 vccd1 _09754_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09684_ _09684_/A vssd1 vssd1 vccd1 vccd1 _18903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14421__591 _14424__594/A vssd1 vssd1 vccd1 vccd1 _18226_/CLK sky130_fd_sc_hd__inv_2
XFILLER_161_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _09118_/A vssd1 vssd1 vccd1 vccd1 _19188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _18568_/Q vssd1 vssd1 vccd1 vccd1 _16291_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_0__f__04012_ clkbuf_0__04012_/X vssd1 vssd1 vccd1 vccd1 _15867__164/A sky130_fd_sc_hd__clkbuf_16
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09049_ _09049_/A vssd1 vssd1 vccd1 vccd1 _19206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _12060_/A _12060_/B vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__or2_1
XFILLER_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _11011_/A vssd1 vssd1 vccd1 vccd1 _18273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04845_ clkbuf_0__04845_/X vssd1 vssd1 vccd1 vccd1 _17049__39/A sky130_fd_sc_hd__clkbuf_16
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12962_ _17963_/Q _17674_/Q _12976_/S vssd1 vssd1 vccd1 vccd1 _12963_/B sky130_fd_sc_hd__mux2_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14463__625 _14463__625/A vssd1 vssd1 vccd1 vccd1 _18260_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_50 _17303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_61 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_72 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11913_ _19242_/Q _19243_/Q _11924_/S vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__mux2_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_83 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ _14607_/X _14694_/Y _14696_/Y _14698_/Y _14700_/Y vssd1 vssd1 vccd1 vccd1
+ _14701_/X sky130_fd_sc_hd__o32a_1
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_94 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ _12893_/A vssd1 vssd1 vccd1 vccd1 _17661_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _17923_/Q _11839_/X _11840_/X _17904_/Q vssd1 vssd1 vccd1 vccd1 _11845_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14662_/S vssd1 vssd1 vccd1 vccd1 _14732_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_205_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17351_ _17340_/X _17351_/B vssd1 vssd1 vccd1 vccd1 _17352_/A sky130_fd_sc_hd__and2b_1
X_14563_ _14594_/A vssd1 vssd1 vccd1 vccd1 _14563_/X sky130_fd_sc_hd__buf_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11775_ _11775_/A vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _18323_/Q _18324_/Q _18325_/Q _18326_/Q _18984_/Q _16511_/A vssd1 vssd1 vccd1
+ vccd1 _16302_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0__f__03589_ clkbuf_0__03589_/X vssd1 vssd1 vccd1 vccd1 _15105__824/A sky130_fd_sc_hd__clkbuf_16
X_13514_ _13240_/X _13499_/A _13513_/X vssd1 vssd1 vccd1 vccd1 _13514_/Y sky130_fd_sc_hd__a21oi_1
X_10726_ _18398_/Q _10704_/X _10726_/S vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17282_ _19264_/Q vssd1 vssd1 vccd1 vccd1 _17288_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19021_ _19027_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16233_ _16229_/X _16232_/X _16271_/S vssd1 vssd1 vccd1 vccd1 _16234_/B sky130_fd_sc_hd__mux2_1
X_13445_ _13140_/X _13437_/X _13444_/Y _13213_/X vssd1 vssd1 vccd1 vccd1 _17796_/D
+ sky130_fd_sc_hd__a211oi_1
X_10657_ _10657_/A vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13376_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13376_/X sky130_fd_sc_hd__buf_4
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16164_ _16214_/A vssd1 vssd1 vccd1 vccd1 _16164_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10588_ _09031_/X _18490_/Q _10594_/S vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__mux2_1
X_15166__873 _15167__874/A vssd1 vssd1 vccd1 vccd1 _18549_/CLK sky130_fd_sc_hd__inv_2
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12327_ _12333_/A vssd1 vssd1 vccd1 vccd1 _12327_/X sky130_fd_sc_hd__buf_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16089__202 _16090__203/A vssd1 vssd1 vccd1 vccd1 _18907_/CLK sky130_fd_sc_hd__inv_2
XFILLER_181_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15046_ _16216_/A _15046_/B vssd1 vssd1 vccd1 vccd1 _15047_/A sky130_fd_sc_hd__and2_1
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04572_ _16646_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04572_/X sky130_fd_sc_hd__clkbuf_16
X_12258_ _12258_/A vssd1 vssd1 vccd1 vccd1 _17552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11209_ _11209_/A vssd1 vssd1 vccd1 vccd1 _18193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03423_ clkbuf_0__03423_/X vssd1 vssd1 vccd1 vccd1 _14886__802/A sky130_fd_sc_hd__clkbuf_16
X_12189_ _12189_/A vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__buf_2
XFILLER_69_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18805_ _18805_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16997_ _13820_/A input77/X _16997_/S vssd1 vssd1 vccd1 vccd1 _16998_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18736_ _18736_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _18873_/Q _15948_/B vssd1 vssd1 vccd1 vccd1 _15954_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18667_ _14157_/A _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _17618_/CLK _17618_/D vssd1 vssd1 vccd1 vccd1 _17618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18598_ _18598_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__04006_ _15831_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04006_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_240_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17549_ _17772_/CLK _17549_/D vssd1 vssd1 vccd1 vccd1 _17549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19219_ _19219_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clkbuf_opt_7_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19143_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _18031_/CLK sky130_fd_sc_hd__clkbuf_16
X_14258__461 _14260__463/A vssd1 vssd1 vccd1 vccd1 _18096_/CLK sky130_fd_sc_hd__inv_2
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04839_ _17013_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04839_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__07558_ _12333_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07558_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09805_ _09805_/A vssd1 vssd1 vccd1 vccd1 _18829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09736_ _18855_/Q _09735_/X _09742_/S vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14527__677 _14527__677/A vssd1 vssd1 vccd1 vccd1 _18312_/CLK sky130_fd_sc_hd__inv_2
XFILLER_243_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09667_ _09667_/A vssd1 vssd1 vccd1 vccd1 _18909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09598_/A vssd1 vssd1 vccd1 vccd1 _18935_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021__16 _17022__17/A vssd1 vssd1 vccd1 vccd1 _19165_/CLK sky130_fd_sc_hd__inv_2
XFILLER_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11560_ _11560_/A vssd1 vssd1 vccd1 vccd1 _17706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _10526_/S vssd1 vssd1 vccd1 vccd1 _10520_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_210_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11491_ _09145_/X _18048_/Q _11491_/S vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13230_ _17738_/Q _13218_/X _13229_/Y vssd1 vssd1 vccd1 vccd1 _17738_/D sky130_fd_sc_hd__o21a_1
XFILLER_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10442_ _10117_/X _18554_/Q _10448_/S vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13161_ _13732_/A vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__buf_8
X_10373_ _10388_/S vssd1 vssd1 vccd1 vccd1 _10382_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_163_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12112_ _12112_/A vssd1 vssd1 vccd1 vccd1 _12112_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13092_ _17701_/Q _13092_/B vssd1 vssd1 vccd1 vccd1 _13096_/A sky130_fd_sc_hd__xor2_1
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15834__137 _15836__139/A vssd1 vssd1 vccd1 vccd1 _18812_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12043_ _12031_/X _12036_/X _12111_/S vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__mux2_1
X_16920_ _19208_/Q _19160_/Q _18271_/Q _18263_/Q _16882_/A _16868_/X vssd1 vssd1 vccd1
+ vccd1 _16920_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16851_ _18244_/Q _18236_/Q _18228_/Q _18220_/Q _16849_/X _16850_/X vssd1 vssd1 vccd1
+ vccd1 _16852_/B sky130_fd_sc_hd__mux4_1
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16782_ _19135_/Q _19133_/Q _16787_/S vssd1 vssd1 vccd1 vccd1 _16783_/B sky130_fd_sc_hd__mux2_1
X_13994_ _17977_/Q _13988_/X _13993_/Y vssd1 vssd1 vccd1 vccd1 _17977_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03170_ _14387_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03170_/X sky130_fd_sc_hd__clkbuf_16
X_18521_ _18521_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16084__198 _16085__199/A vssd1 vssd1 vccd1 vccd1 _18903_/CLK sky130_fd_sc_hd__inv_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12945_/A vssd1 vssd1 vccd1 vccd1 _17669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14428__597 _14430__599/A vssd1 vssd1 vccd1 vccd1 _18232_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18452_ _18452_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12876_/A vssd1 vssd1 vccd1 vccd1 _17656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17403_ _17409_/A vssd1 vssd1 vccd1 vccd1 _17403_/X sky130_fd_sc_hd__buf_1
X_14615_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__buf_4
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _13830_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _14053_/A sky130_fd_sc_hd__and2_2
XFILLER_18_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18383_ _18383_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _18653_/Q _15595_/B _15595_/C vssd1 vssd1 vccd1 vccd1 _15605_/C sky130_fd_sc_hd__and3_1
XFILLER_14_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17334_ _17323_/X _17334_/B vssd1 vssd1 vccd1 vccd1 _17335_/A sky130_fd_sc_hd__and2b_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11758_ _17863_/Q _17703_/Q _18000_/Q vssd1 vssd1 vccd1 vccd1 _11759_/A sky130_fd_sc_hd__mux2_4
X_14546_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14546_/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__03972_ clkbuf_0__03972_/X vssd1 vssd1 vccd1 vccd1 _15704__999/A sky130_fd_sc_hd__clkbuf_16
XFILLER_230_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10709_ _10709_/A vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__clkbuf_1
X_17265_ _17270_/C _17265_/B _17265_/C vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__and3b_1
XFILLER_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11689_ _19036_/Q _16613_/B vssd1 vssd1 vccd1 vccd1 _16614_/B sky130_fd_sc_hd__and2_1
XFILLER_128_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19004_ _19004_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
X_16216_ _16216_/A vssd1 vssd1 vccd1 vccd1 _16216_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13428_ _13428_/A vssd1 vssd1 vccd1 vccd1 _16736_/A sky130_fd_sc_hd__buf_4
X_17196_ _17239_/A vssd1 vssd1 vccd1 vccd1 _17235_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13359_ _16690_/A vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__buf_4
X_16147_ _10406_/A _16137_/Y _16140_/Y _16142_/Y _16146_/Y vssd1 vssd1 vccd1 vccd1
+ _16147_/X sky130_fd_sc_hd__o32a_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15029_ _15029_/A vssd1 vssd1 vccd1 vccd1 _18464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03406_ clkbuf_0__03406_/X vssd1 vssd1 vccd1 vccd1 _14799__732/A sky130_fd_sc_hd__clkbuf_16
XFILLER_110_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 flash_io0_we vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09521_ _09521_/A vssd1 vssd1 vccd1 vccd1 _18999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18719_ _18719_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _14651_/A _09456_/A vssd1 vssd1 vccd1 vccd1 _09453_/C sky130_fd_sc_hd__or2_1
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03199_ clkbuf_0__03199_/X vssd1 vssd1 vccd1 vccd1 _14744__689/A sky130_fd_sc_hd__clkbuf_16
XFILLER_240_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09383_ _09383_/A vssd1 vssd1 vccd1 vccd1 _19073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03090_ clkbuf_0__03090_/X vssd1 vssd1 vccd1 vccd1 _14150__434/A sky130_fd_sc_hd__clkbuf_16
XFILLER_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03992_ clkbuf_0__03992_/X vssd1 vssd1 vccd1 vccd1 _15801__121/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12336__397 _12338__399/A vssd1 vssd1 vccd1 vccd1 _17578_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _10833_/B _10691_/B vssd1 vssd1 vccd1 vccd1 _09742_/S sky130_fd_sc_hd__nor2_1
X_10991_ _10991_/A vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117__834 _15117__834/A vssd1 vssd1 vccd1 vccd1 _18510_/CLK sky130_fd_sc_hd__inv_2
X_12730_ _12737_/C _12737_/D vssd1 vssd1 vccd1 vccd1 _12732_/A sky130_fd_sc_hd__and2_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A vssd1 vssd1 vccd1 vccd1 _17606_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11612_ _11612_/A vssd1 vssd1 vccd1 vccd1 _17568_/D sky130_fd_sc_hd__clkbuf_1
X_14400_ _14400_/A vssd1 vssd1 vccd1 vccd1 _14400_/X sky130_fd_sc_hd__buf_1
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12592_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__clkbuf_2
X_15380_ _15281_/A _15379_/Y _15305_/A vssd1 vssd1 vccd1 vccd1 _15380_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_230_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11543_ _08883_/X _17713_/Q _11545_/S vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__mux2_1
X_14331_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14331_/X sky130_fd_sc_hd__buf_1
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ _14293_/A vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__buf_1
X_17050_ _17062_/A vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__buf_1
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ _11474_/A vssd1 vssd1 vccd1 vccd1 _18056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13213_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_125_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16001_ _16002_/B _16002_/C _18869_/Q vssd1 vssd1 vccd1 vccd1 _16003_/B sky130_fd_sc_hd__a21oi_1
XFILLER_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ _09975_/C _10424_/X _10407_/X vssd1 vssd1 vccd1 vccd1 _10425_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_183_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14193_ _14193_/A vssd1 vssd1 vccd1 vccd1 _18068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13144_ _13216_/B vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__buf_2
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _18592_/Q _09718_/X _10364_/S vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13075_ _13075_/A vssd1 vssd1 vccd1 vccd1 _17701_/D sky130_fd_sc_hd__clkbuf_1
X_17952_ _17959_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
X_15753__1039 _15753__1039/A vssd1 vssd1 vccd1 vccd1 _18756_/CLK sky130_fd_sc_hd__inv_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10287_ _10287_/A vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12026_ _11901_/X _12025_/X _12036_/S vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__mux2_1
X_16903_ _16897_/X _16901_/X _16980_/S vssd1 vssd1 vccd1 vccd1 _16903_/X sky130_fd_sc_hd__mux2_1
X_17883_ _18021_/CLK _17883_/D vssd1 vssd1 vccd1 vccd1 _17883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16834_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16834_/X sky130_fd_sc_hd__buf_4
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16765_ _19091_/Q vssd1 vssd1 vccd1 vccd1 _16765_/X sky130_fd_sc_hd__clkbuf_2
X_13977_ _17971_/Q _13967_/X _13976_/Y vssd1 vssd1 vccd1 vccd1 _17971_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03153_ _14300_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03153_/X sky130_fd_sc_hd__clkbuf_16
X_18504_ _18504_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _17659_/Q _12924_/X _12834_/X _17654_/Q _12927_/X vssd1 vssd1 vccd1 vccd1
+ _12931_/C sky130_fd_sc_hd__o221a_1
XFILLER_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18435_ _18435_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ _15535_/A _15642_/X _15615_/B _15628_/X vssd1 vssd1 vccd1 vccd1 _18670_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12859_ _12859_/A _12859_/B _12859_/C _12858_/X vssd1 vssd1 vccd1 vccd1 _12860_/D
+ sky130_fd_sc_hd__or4b_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18366_ _18366_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15578_ _15585_/B _15585_/C vssd1 vssd1 vccd1 vccd1 _15584_/B sky130_fd_sc_hd__and2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17317_ _17304_/X _17317_/B vssd1 vssd1 vccd1 vccd1 _17318_/A sky130_fd_sc_hd__and2b_1
XFILLER_222_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18297_ _18297_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
X_17248_ _17252_/B _17265_/B _17248_/C vssd1 vssd1 vccd1 vccd1 _17249_/A sky130_fd_sc_hd__and3b_1
XPeripherals_170 vssd1 vssd1 vccd1 vccd1 Peripherals_170/HI io_oeb[33] sky130_fd_sc_hd__conb_1
Xclkbuf_0__03986_ _15773_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03986_/X sky130_fd_sc_hd__clkbuf_16
XPeripherals_181 vssd1 vssd1 vccd1 vccd1 Peripherals_181/HI wb_data_o[20] sky130_fd_sc_hd__conb_1
XFILLER_175_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPeripherals_192 vssd1 vssd1 vccd1 vccd1 Peripherals_192/HI wb_data_o[31] sky130_fd_sc_hd__conb_1
XFILLER_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _19237_/Q _17179_/B vssd1 vssd1 vccd1 vccd1 _17186_/D sky130_fd_sc_hd__and2_1
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08952_ _09682_/A vssd1 vssd1 vccd1 vccd1 _08952_/X sky130_fd_sc_hd__buf_4
XFILLER_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08883_ _18988_/Q vssd1 vssd1 vccd1 vccd1 _08883_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04369_ clkbuf_0__04369_/X vssd1 vssd1 vccd1 vccd1 _16318__217/A sky130_fd_sc_hd__clkbuf_16
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659__295 _16659__295/A vssd1 vssd1 vccd1 vccd1 _19069_/CLK sky130_fd_sc_hd__inv_2
X_09504_ _18880_/Q vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09435_ _19047_/Q vssd1 vssd1 vccd1 vccd1 _14615_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09366_ _09366_/A vssd1 vssd1 vccd1 vccd1 _19080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09297_ _19113_/Q _08964_/X _09299_/S vssd1 vssd1 vccd1 vccd1 _09298_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16332__229 _16332__229/A vssd1 vssd1 vccd1 vccd1 _18945_/CLK sky130_fd_sc_hd__inv_2
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _10210_/A vssd1 vssd1 vccd1 vccd1 _18683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11190_ _18201_/Q _11047_/X _11196_/S vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10141_ _18710_/Q _10048_/X _10149_/S vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__mux2_1
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ _10135_/A vssd1 vssd1 vccd1 vccd1 _10072_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03975_ clkbuf_0__03975_/X vssd1 vssd1 vccd1 vccd1 _15720__1012/A sky130_fd_sc_hd__clkbuf_16
XFILLER_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13900_ _17943_/Q _13879_/X _13899_/Y vssd1 vssd1 vccd1 vccd1 _17943_/D sky130_fd_sc_hd__o21a_1
XFILLER_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13831_ _13847_/B vssd1 vssd1 vccd1 vccd1 _13845_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16550_ _16639_/A vssd1 vssd1 vccd1 vccd1 _16550_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_208 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ _13762_/A vssd1 vssd1 vccd1 vccd1 _13762_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10974_ _10974_/A vssd1 vssd1 vccd1 vccd1 _18288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_219 _17826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15501_ _15501_/A _15501_/B vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__nand2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12713_ _12713_/A _12713_/B vssd1 vssd1 vccd1 vccd1 _17621_/D sky130_fd_sc_hd__nor2_1
X_16481_ _18978_/Q _16482_/C _18979_/Q vssd1 vssd1 vccd1 vccd1 _16483_/B sky130_fd_sc_hd__a21oi_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13693_ _17874_/Q _13682_/X _13692_/Y vssd1 vssd1 vccd1 vccd1 _17874_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f__04527_ clkbuf_0__04527_/X vssd1 vssd1 vccd1 vccd1 _16548__259/A sky130_fd_sc_hd__clkbuf_16
XFILLER_245_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ _18220_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
X_12644_ _12647_/C _12644_/B vssd1 vssd1 vccd1 vccd1 _17601_/D sky130_fd_sc_hd__nor2_1
XFILLER_188_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _18151_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
X_12575_ _17631_/Q vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15363_ _15281_/A _15362_/Y _15285_/X vssd1 vssd1 vccd1 vccd1 _15363_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_184_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03409_ clkbuf_0__03409_/X vssd1 vssd1 vccd1 vccd1 _14813__743/A sky130_fd_sc_hd__clkbuf_16
XFILLER_196_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17102_ _12298_/A _17097_/X _17100_/X _17101_/X vssd1 vssd1 vccd1 vccd1 _17102_/Y
+ sky130_fd_sc_hd__a31oi_1
X_18082_ _19337_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
X_11526_ _11526_/A vssd1 vssd1 vccd1 vccd1 _18033_/D sky130_fd_sc_hd__clkbuf_1
X_15294_ _19319_/Q _19303_/Q _19295_/Q _19270_/Q _15293_/X _15218_/X vssd1 vssd1 vccd1
+ vccd1 _15294_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14245_ _09253_/X _14244_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _15080_/B sky130_fd_sc_hd__a21oi_4
X_11457_ _11457_/A hold23/X vssd1 vssd1 vccd1 vccd1 _11473_/S sky130_fd_sc_hd__or2_2
XFILLER_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10408_ _10391_/X _10406_/X _10407_/X vssd1 vssd1 vccd1 vccd1 _10408_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11388_ _11326_/X _18121_/Q _11394_/S vssd1 vssd1 vccd1 vccd1 _11389_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14174__451 _14177__454/A vssd1 vssd1 vccd1 vccd1 _18059_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _14113_/B vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__inv_2
X_10339_ _18477_/Q vssd1 vssd1 vccd1 vccd1 _10339_/X sky130_fd_sc_hd__buf_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _19013_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13058_ _13049_/X _13058_/B vssd1 vssd1 vccd1 vccd1 _13059_/A sky130_fd_sc_hd__and2b_1
X_17935_ _17935_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12009_ _12004_/X _12005_/X _12006_/X _12008_/X _12087_/S _12098_/S vssd1 vssd1 vccd1
+ vccd1 _12009_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17866_ _17881_/CLK _17866_/D vssd1 vssd1 vccd1 vccd1 _17866_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_226_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16817_ _16808_/X _16816_/X _16875_/S vssd1 vssd1 vccd1 vccd1 _16817_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17797_ _19135_/CLK _17797_/D vssd1 vssd1 vccd1 vccd1 _17797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16748_ _19128_/Q _16746_/X _16748_/S vssd1 vssd1 vccd1 vccd1 _16749_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16732__345 _16735__348/A vssd1 vssd1 vccd1 vccd1 _19124_/CLK sky130_fd_sc_hd__inv_2
X_09220_ _09220_/A vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__clkbuf_1
X_18418_ _18418_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19398_ input22/X vssd1 vssd1 vccd1 vccd1 _19398_/X sky130_fd_sc_hd__buf_4
XFILLER_222_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _09166_/S vssd1 vssd1 vccd1 vccd1 _09160_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18349_ _18349_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09082_ _09770_/B _10770_/B _10770_/A vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__nand3b_4
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput60 wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__03969_ _15686_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03969_/X sky130_fd_sc_hd__clkbuf_16
Xinput71 wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_6
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09984_ _18771_/Q _09951_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08935_ _08935_/A vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ _19315_/Q _08830_/X _08878_/S vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__mux2_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _08797_/A vssd1 vssd1 vccd1 vccd1 _19344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ _08917_/X _19057_/Q _09424_/S vssd1 vssd1 vccd1 vccd1 _09419_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _10690_/A vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__clkbuf_4
X_15752__1038 _15753__1039/A vssd1 vssd1 vccd1 vccd1 _18755_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _09349_/A vssd1 vssd1 vccd1 vccd1 _19087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ _12353_/X _12357_/X _12390_/S vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11311_ _11153_/X _18151_/Q _11313_/S vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__mux2_1
X_12291_ _12280_/X _12291_/B vssd1 vssd1 vccd1 vccd1 _12292_/A sky130_fd_sc_hd__and2b_1
XFILLER_181_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14030_ _17991_/Q _14012_/X _14029_/Y vssd1 vssd1 vccd1 vccd1 _17991_/D sky130_fd_sc_hd__o21a_1
XFILLER_49_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11242_ _11257_/S vssd1 vssd1 vccd1 vccd1 _11251_/S sky130_fd_sc_hd__buf_2
XFILLER_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14351__536 _14352__537/A vssd1 vssd1 vccd1 vccd1 _18171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11173_ _11173_/A vssd1 vssd1 vccd1 vccd1 _18209_/D sky130_fd_sc_hd__clkbuf_1
X_15160__868 _15161__869/A vssd1 vssd1 vccd1 vccd1 _18544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ _10123_/X _18715_/Q _10127_/S vssd1 vssd1 vccd1 vccd1 _10125_/A sky130_fd_sc_hd__mux2_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _15985_/B _15993_/B vssd1 vssd1 vccd1 vccd1 _15981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _19040_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _17720_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ _14964_/A _14962_/B _14961_/B _14961_/D vssd1 vssd1 vccd1 vccd1 _14955_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10055_ _18741_/Q _10054_/X _10064_/S vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__mux2_1
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _18013_/CLK _17651_/D vssd1 vssd1 vccd1 vccd1 _17651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _16602_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16602_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13814_ _17915_/Q _13797_/X _13813_/Y vssd1 vssd1 vccd1 vccd1 _17915_/D sky130_fd_sc_hd__o21a_1
XFILLER_235_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17582_ _17582_/CLK _17582_/D vssd1 vssd1 vccd1 vccd1 _17582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19321_ _19321_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
X_16533_ _16533_/A vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__clkbuf_1
X_13745_ _13757_/B vssd1 vssd1 vccd1 vccd1 _13755_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10957_ _08874_/X _18295_/Q _10959_/S vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19252_ _19252_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ _16464_/A _16464_/B vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__nor2_1
XFILLER_176_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13676_ _17868_/Q _13660_/X _13675_/Y vssd1 vssd1 vccd1 vccd1 _17868_/D sky130_fd_sc_hd__o21a_1
X_10888_ _10931_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _10911_/S sky130_fd_sc_hd__nor2_2
X_18203_ _18203_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ _12626_/A _12626_/B _12617_/X vssd1 vssd1 vccd1 vccd1 _12628_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_1__f__04841_ clkbuf_0__04841_/X vssd1 vssd1 vccd1 vccd1 _17030__24/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19183_ _19183_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _16393_/B _16393_/C _16466_/B vssd1 vssd1 vccd1 vccd1 _16419_/C sky130_fd_sc_hd__a21oi_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18134_ _18134_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
X_15346_ _15281_/A _15345_/Y _15285_/X vssd1 vssd1 vccd1 vccd1 _15346_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1__f__07560_ clkbuf_0__07560_/X vssd1 vssd1 vccd1 vccd1 _12348__407/A sky130_fd_sc_hd__clkbuf_16
X_12558_ _12487_/X _12489_/X _12513_/X _12557_/X _12449_/S _12504_/A vssd1 vssd1 vccd1
+ vccd1 _12558_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11509_ _18040_/Q _11344_/A _11509_/S vssd1 vssd1 vccd1 vccd1 _11510_/A sky130_fd_sc_hd__mux2_1
X_18065_ _18870_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_1__f__07491_ clkbuf_0__07491_/X vssd1 vssd1 vccd1 vccd1 _12230__375/A sky130_fd_sc_hd__clkbuf_16
X_15277_ _18830_/Q _18822_/Q _18814_/Q _18681_/Q _15214_/X _15225_/X vssd1 vssd1 vccd1
+ vccd1 _15277_/X sky130_fd_sc_hd__mux4_1
X_12489_ _12706_/B _12706_/A _17621_/Q _17622_/Q _12555_/A _12487_/S vssd1 vssd1 vccd1
+ vccd1 _12489_/X sky130_fd_sc_hd__mux4_2
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14228_ _14228_/A vssd1 vssd1 vccd1 vccd1 _18084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _14293_/A vssd1 vssd1 vccd1 vccd1 _14159_/X sky130_fd_sc_hd__buf_1
XFILLER_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03585_ clkbuf_0__03585_/X vssd1 vssd1 vccd1 vccd1 _15091__814/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252__456 _14252__456/A vssd1 vssd1 vccd1 vccd1 _18091_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18967_ _19013_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17779_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17918_ _17923_/CLK _17918_/D vssd1 vssd1 vccd1 vccd1 _17918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18898_ _18898_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434__929 _15434__929/A vssd1 vssd1 vccd1 vccd1 _18616_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17849_ _17850_/CLK _17849_/D vssd1 vssd1 vccd1 vccd1 _17849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ _09203_/A vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ _19184_/Q _09133_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ _19202_/Q _08868_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _09066_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _10135_/A vssd1 vssd1 vccd1 vccd1 _09967_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _08917_/X _19298_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 _08919_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09913_/S vssd1 vssd1 vccd1 vccd1 _09907_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _19046_/Q hold21/A vssd1 vssd1 vccd1 vccd1 _09440_/B sky130_fd_sc_hd__or2b_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11860_/A vssd1 vssd1 vccd1 vccd1 _11860_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10811_/A vssd1 vssd1 vccd1 vccd1 _18364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11791_ _13645_/B _11791_/B vssd1 vssd1 vccd1 vccd1 _11840_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__08201_ clkbuf_0__08201_/X vssd1 vssd1 vccd1 vccd1 _13120__423/A sky130_fd_sc_hd__clkbuf_16
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _13529_/X _13523_/X _13513_/X vssd1 vssd1 vccd1 vccd1 _13530_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_242_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10742_ _18391_/Q _10701_/X _10744_/S vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13461_ _13484_/S vssd1 vssd1 vccd1 vccd1 _13477_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10673_ _10688_/S vssd1 vssd1 vccd1 vccd1 _10682_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_139_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12412_ _12373_/Y _12381_/Y _12392_/Y _12405_/Y _12408_/X _12560_/S vssd1 vssd1 vccd1
+ vccd1 _12773_/B sky130_fd_sc_hd__mux4_1
XFILLER_159_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16180_ _16178_/X _16179_/X _16248_/S vssd1 vssd1 vccd1 vccd1 _16180_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13392_ _13681_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13395_/A sky130_fd_sc_hd__nor2_1
XFILLER_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15131_ _15131_/A vssd1 vssd1 vccd1 vccd1 _15131_/X sky130_fd_sc_hd__buf_1
XFILLER_103_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12274_ _17557_/Q _18020_/Q _12287_/S vssd1 vssd1 vccd1 vccd1 _12275_/B sky130_fd_sc_hd__mux2_1
XFILLER_142_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15062_ _18472_/Q vssd1 vssd1 vccd1 vccd1 _15062_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14013_ _13717_/A _14012_/X _14005_/X vssd1 vssd1 vccd1 vccd1 _14013_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_175_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11225_ _11142_/X _18186_/Q _11233_/S vssd1 vssd1 vccd1 vccd1 _11226_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11156_ _11335_/A vssd1 vssd1 vccd1 vccd1 _11156_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18821_ _18821_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10107_ _10107_/A vssd1 vssd1 vccd1 vccd1 _18721_/D sky130_fd_sc_hd__clkbuf_1
X_18752_ _18752_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ _11365_/B vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__buf_4
X_15964_ _18862_/Q _15967_/C vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _17703_/CLK _17703_/D vssd1 vssd1 vccd1 vccd1 _17703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14915_ _17851_/Q _17850_/Q _14938_/A _17849_/Q vssd1 vssd1 vccd1 vccd1 _14916_/B
+ sky130_fd_sc_hd__o31ai_1
X_10038_ _18747_/Q _09951_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18683_ _18683_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17634_ _18012_/CLK _17634_/D vssd1 vssd1 vccd1 vccd1 _17634_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14846_ _14852_/A vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__buf_1
XFILLER_64_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17565_ _17565_/CLK _17565_/D vssd1 vssd1 vccd1 vccd1 _17565_/Q sky130_fd_sc_hd__dfxtp_1
X_14777_ _14808_/A vssd1 vssd1 vccd1 vccd1 _14777_/X sky130_fd_sc_hd__buf_1
X_11989_ _11974_/X _11977_/X _11982_/X _12091_/B _12037_/S _12098_/S vssd1 vssd1 vccd1
+ vccd1 _11990_/B sky130_fd_sc_hd__mux4_1
X_19304_ _19304_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
X_16516_ _08997_/C _09252_/A _16559_/B _16516_/D vssd1 vssd1 vccd1 vccd1 _16532_/C
+ sky130_fd_sc_hd__and4bb_2
XFILLER_220_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13728_ _13783_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13728_/Y sky130_fd_sc_hd__nor2_1
XFILLER_210_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17496_ _17477_/Y _17485_/X _17495_/X _19340_/Q vssd1 vssd1 vccd1 vccd1 _17497_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19235_ _19248_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16447_ _18971_/Q _16468_/B vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__nand2_1
X_13659_ _13666_/A vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19166_ _19166_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_1
X_16378_ _16422_/B _16378_/B vssd1 vssd1 vccd1 vccd1 _16379_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18117_ _18117_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_1
X_15329_ _09614_/A _15328_/Y _15285_/X vssd1 vssd1 vccd1 vccd1 _15329_/Y sky130_fd_sc_hd__a21oi_1
X_19097_ _19097_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03806_ _15448_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03806_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_219_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _18048_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _09821_/A vssd1 vssd1 vccd1 vccd1 _18822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15751__1037 _15753__1039/A vssd1 vssd1 vccd1 vccd1 _18754_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16697__321 _16697__321/A vssd1 vssd1 vccd1 vccd1 _19096_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _18885_/Q vssd1 vssd1 vccd1 vccd1 _09752_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03599_ _15155_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03599_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09683_ _09682_/X _18903_/Q _09689_/S vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15111__829 _15111__829/A vssd1 vssd1 vccd1 vccd1 _18505_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _19188_/Q _09116_/X _09117_/S vssd1 vssd1 vccd1 vccd1 _09118_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04011_ clkbuf_0__04011_/X vssd1 vssd1 vccd1 vccd1 _15890_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_163_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09048_ _09047_/X _19206_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155__438 _14155__438/A vssd1 vssd1 vccd1 vccd1 _18046_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _09031_/X _18273_/Q _11016_/S vssd1 vssd1 vccd1 vccd1 _11011_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04844_ clkbuf_0__04844_/X vssd1 vssd1 vccd1 vccd1 _17062_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _12999_/S vssd1 vssd1 vccd1 vccd1 _12976_/S sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_40 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_51 _17454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_62 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14700_ _14640_/X _14699_/X _14604_/A vssd1 vssd1 vccd1 vccd1 _14700_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_73 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11912_ _11908_/X _11910_/X _12067_/S vssd1 vssd1 vccd1 vccd1 _11912_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_84 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15686_/A vssd1 vssd1 vccd1 vccd1 _15680_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_95 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12892_ _12877_/X _12892_/B vssd1 vssd1 vccd1 vccd1 _12893_/A sky130_fd_sc_hd__and2b_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14626_/X _14630_/X _14673_/S vssd1 vssd1 vccd1 vccd1 _14631_/X sky130_fd_sc_hd__mux2_2
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11843_/A vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17350_ _17755_/Q _19288_/Q _17350_/S vssd1 vssd1 vccd1 vccd1 _17351_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14562_ _14572_/A vssd1 vssd1 vccd1 vccd1 _14688_/S sky130_fd_sc_hd__buf_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11774_ _11774_/A input7/X vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__and2_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _18985_/Q vssd1 vssd1 vccd1 vccd1 _16511_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_0__f__03588_ clkbuf_0__03588_/X vssd1 vssd1 vccd1 vccd1 _15099__819/A sky130_fd_sc_hd__clkbuf_16
X_13513_ _13689_/A vssd1 vssd1 vccd1 vccd1 _13513_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_213_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17281_ _17288_/C _17284_/C _17280_/Y vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__a21oi_1
XFILLER_198_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10725_ _10725_/A vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14493_ _14505_/A vssd1 vssd1 vccd1 vccd1 _14493_/X sky130_fd_sc_hd__buf_1
XFILLER_207_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19020_ _19027_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
X_16232_ _16230_/X _16231_/X _18566_/Q vssd1 vssd1 vccd1 vccd1 _16232_/X sky130_fd_sc_hd__mux2_1
X_13444_ _17796_/Q _13444_/B vssd1 vssd1 vccd1 vccd1 _13444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10656_ _18428_/Q _09718_/X _10662_/S vssd1 vssd1 vccd1 vccd1 _10657_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16351__243 _16352__244/A vssd1 vssd1 vccd1 vccd1 _18959_/CLK sky130_fd_sc_hd__inv_2
X_16163_ _16234_/A _16163_/B vssd1 vssd1 vccd1 vccd1 _16163_/Y sky130_fd_sc_hd__nand2_1
X_13375_ _13414_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _13375_/Y sky130_fd_sc_hd__nor2_1
X_10587_ _10587_/A vssd1 vssd1 vccd1 vccd1 _18491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12326_ _13109_/A vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__buf_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15045_ _18467_/Q _14967_/X _15044_/Y _15026_/X vssd1 vssd1 vccd1 vccd1 _15046_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__04571_ _16645_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04571_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_79_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12257_ _12245_/X _12257_/B vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__and2b_1
XFILLER_218_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03422_ clkbuf_0__03422_/X vssd1 vssd1 vccd1 vccd1 _14881__798/A sky130_fd_sc_hd__clkbuf_16
X_11208_ _18193_/Q _11047_/X _11214_/S vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__mux2_1
X_12188_ _17530_/Q _12185_/X _12187_/X _17516_/Q vssd1 vssd1 vccd1 vccd1 _12192_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18804_ _18804_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
X_11139_ _11139_/A vssd1 vssd1 vccd1 vccd1 _18220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16996_ _16996_/A vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15947_ _15947_/A _15947_/B vssd1 vssd1 vccd1 vccd1 _15948_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18735_ _18735_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18666_ _14157_/A _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14364__546 _14364__546/A vssd1 vssd1 vccd1 vccd1 _18181_/CLK sky130_fd_sc_hd__inv_2
XFILLER_188_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17617_ _17618_/CLK _17617_/D vssd1 vssd1 vccd1 vccd1 _17617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14776__714 _14776__714/A vssd1 vssd1 vccd1 vccd1 _18357_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18597_ _18597_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17405__96 _17405__96/A vssd1 vssd1 vccd1 vccd1 _19309_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__04005_ _15830_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04005_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17548_ _17772_/CLK _17548_/D vssd1 vssd1 vccd1 vccd1 _17548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17479_ _19330_/Q _12202_/A _12212_/X _19332_/Q vssd1 vssd1 vccd1 vccd1 _17485_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19218_ _19218_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19149_ _19149_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15702__997 _15704__999/A vssd1 vssd1 vccd1 vccd1 _18714_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__04838_ _17012_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04838_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__07557_ _12327_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07557_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_62_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _17951_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_236_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09804_ _18829_/Q _09764_/X _09806_/S vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09735_ _10707_/A vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09666_ _18909_/Q _09271_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14265__466 _14265__466/A vssd1 vssd1 vccd1 vccd1 _18101_/CLK sky130_fd_sc_hd__inv_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09597_ _18935_/Q _09504_/X _09597_/S vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__mux2_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10510_ _10528_/B _10510_/B vssd1 vssd1 vccd1 vccd1 _10526_/S sky130_fd_sc_hd__nor2_2
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ _11490_/A vssd1 vssd1 vccd1 vccd1 _18049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _10441_/A vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13160_ input73/X _13210_/B vssd1 vssd1 vccd1 vccd1 _13732_/A sky130_fd_sc_hd__nand2_1
X_10372_ _10372_/A hold2/X vssd1 vssd1 vccd1 vccd1 _10388_/S sky130_fd_sc_hd__or2_2
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12111_ _12035_/X _12067_/X _12111_/S vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13091_ _17693_/Q _12924_/X _12920_/A _17695_/Q vssd1 vssd1 vccd1 vccd1 _13097_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12042_ _12023_/X _12032_/X _12111_/S vssd1 vssd1 vccd1 vccd1 _12108_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16850_ _16894_/A vssd1 vssd1 vccd1 vccd1 _16850_/X sky130_fd_sc_hd__buf_2
XFILLER_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11879__362 _11879__362/A vssd1 vssd1 vccd1 vccd1 _17509_/CLK sky130_fd_sc_hd__inv_2
X_16781_ _19134_/Q _16786_/B vssd1 vssd1 vccd1 vccd1 _16781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13993_ _13400_/A _13989_/X _13992_/X vssd1 vssd1 vccd1 vccd1 _13993_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18520_ _18520_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _16620_/A _12944_/B _12944_/C vssd1 vssd1 vccd1 vccd1 _12945_/A sky130_fd_sc_hd__and3b_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18451_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12875_ _12830_/X _12875_/B vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__and2b_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14614_ _14679_/A _14614_/B vssd1 vssd1 vccd1 vccd1 _14614_/Y sky130_fd_sc_hd__nor2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11826_/A vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18382_ _18382_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15595_/B _15595_/C _18653_/Q vssd1 vssd1 vccd1 vccd1 _15596_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17333_ _17760_/Q _19283_/Q _17333_/S vssd1 vssd1 vccd1 vccd1 _17334_/B sky130_fd_sc_hd__mux2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14545_ _14594_/A vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__buf_4
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11757_ _11757_/A vssd1 vssd1 vccd1 vccd1 _11757_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_230_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03971_ clkbuf_0__03971_/X vssd1 vssd1 vccd1 vccd1 _15696__992/A sky130_fd_sc_hd__clkbuf_16
XFILLER_187_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15750__1036 _15750__1036/A vssd1 vssd1 vccd1 vccd1 _18753_/CLK sky130_fd_sc_hd__inv_2
X_17264_ _17264_/A _17264_/B vssd1 vssd1 vccd1 vccd1 _17265_/C sky130_fd_sc_hd__or2_1
XFILLER_119_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10708_ _18405_/Q _10707_/X _10714_/S vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _19035_/Q _19034_/Q _16608_/B vssd1 vssd1 vccd1 vccd1 _16613_/B sky130_fd_sc_hd__and3_1
X_19003_ _19003_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16215_ _16190_/X _16203_/X _16213_/Y _16214_/X vssd1 vssd1 vccd1 vccd1 _16215_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_146_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13427_ _13432_/S _13709_/A _13426_/Y _13213_/X vssd1 vssd1 vccd1 vccd1 _17792_/D
+ sky130_fd_sc_hd__a211oi_1
X_17195_ _17195_/A _17203_/D vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__and2_1
X_10639_ _10654_/S vssd1 vssd1 vccd1 vccd1 _10648_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16146_ _16143_/X _16145_/X _16119_/X vssd1 vssd1 vccd1 vccd1 _16146_/Y sky130_fd_sc_hd__o21ai_1
X_13358_ _13740_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _13358_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _17552_/Q _12206_/X _12199_/X _17559_/Q _12308_/Y vssd1 vssd1 vccd1 vccd1
+ _12309_/X sky130_fd_sc_hd__o221a_1
XFILLER_142_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _13231_/X _13288_/X _13275_/X vssd1 vssd1 vccd1 vccd1 _13289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15028_ _15034_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _15029_/A sky130_fd_sc_hd__and2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03405_ clkbuf_0__03405_/X vssd1 vssd1 vccd1 vccd1 _14795__729/A sky130_fd_sc_hd__clkbuf_16
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 flash_io0_write vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_16979_ _16977_/X _16978_/X _16979_/S vssd1 vssd1 vccd1 vccd1 _16979_/X sky130_fd_sc_hd__mux2_1
X_09520_ _18999_/Q _09498_/X _09524_/S vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__mux2_1
X_18718_ _18718_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09451_ _16559_/B vssd1 vssd1 vccd1 vccd1 _09477_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18649_ _18654_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03198_ clkbuf_0__03198_/X vssd1 vssd1 vccd1 vccd1 _14532__681/A sky130_fd_sc_hd__clkbuf_16
XFILLER_224_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16358__249 _16358__249/A vssd1 vssd1 vccd1 vccd1 _18965_/CLK sky130_fd_sc_hd__inv_2
X_09382_ _19073_/Q _08949_/X _09388_/S vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14533__682 _14535__684/A vssd1 vssd1 vccd1 vccd1 _18317_/CLK sky130_fd_sc_hd__inv_2
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03991_ clkbuf_0__03991_/X vssd1 vssd1 vccd1 vccd1 _15798__119/A sky130_fd_sc_hd__clkbuf_16
XFILLER_43_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453__943 _15453__943/A vssd1 vssd1 vccd1 vccd1 _18630_/CLK sky130_fd_sc_hd__inv_2
XFILLER_142_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09718_ _10690_/A vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__buf_4
XFILLER_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10990_ _18282_/Q _09119_/X _10998_/S vssd1 vssd1 vccd1 vccd1 _10991_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _09645_/X _09649_/B _09649_/C vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__and3b_1
XFILLER_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12658_/X _12759_/A _12660_/C vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__and3b_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _17568_/Q _10704_/A _11611_/S vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12591_ _14065_/B _12527_/X _12563_/X _12574_/X _12590_/X vssd1 vssd1 vccd1 vccd1
+ _12616_/A sky130_fd_sc_hd__o2111a_2
XFILLER_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15840__142 _15840__142/A vssd1 vssd1 vccd1 vccd1 _18817_/CLK sky130_fd_sc_hd__inv_2
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11542_ _11542_/A vssd1 vssd1 vccd1 vccd1 _17714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11473_ _11344_/X _18056_/Q _11473_/S vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _15997_/Y _15999_/Y _15982_/X vssd1 vssd1 vccd1 vccd1 _18868_/D sky130_fd_sc_hd__a21oi_1
X_13212_ _17736_/Q _13212_/B vssd1 vssd1 vccd1 vccd1 _13212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10424_ _10424_/A _10424_/B _10424_/C vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__and3_1
XFILLER_171_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14192_ _18068_/Q input48/X _14196_/S vssd1 vssd1 vccd1 vccd1 _14193_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14315__507 _14317__509/A vssd1 vssd1 vccd1 vccd1 _18142_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13143_ _13135_/X _13140_/X _13142_/Y _16619_/A vssd1 vssd1 vccd1 vccd1 _17723_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10355_ _10370_/S vssd1 vssd1 vccd1 vccd1 _10364_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _13066_/X _13074_/B vssd1 vssd1 vccd1 vccd1 _13075_/A sky130_fd_sc_hd__and2b_1
X_17951_ _17951_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _18619_/Q _10192_/X _10290_/S vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12025_ _19254_/Q _19255_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16902_ _16902_/A vssd1 vssd1 vccd1 vccd1 _16980_/S sky130_fd_sc_hd__clkbuf_2
X_17882_ _18021_/CLK _17882_/D vssd1 vssd1 vccd1 vccd1 _17882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16833_ _16929_/A _16833_/B vssd1 vssd1 vccd1 vccd1 _16833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16764_ _16775_/A _16764_/B vssd1 vssd1 vccd1 vccd1 _19130_/D sky130_fd_sc_hd__nor2_1
XFILLER_219_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13976_ _13669_/X _13973_/X _13920_/X vssd1 vssd1 vccd1 vccd1 _13976_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03152_ _14294_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03152_/X sky130_fd_sc_hd__clkbuf_16
X_18503_ _18503_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ _17665_/Q _12846_/B _12838_/X _17668_/Q _12926_/Y vssd1 vssd1 vccd1 vccd1
+ _12927_/X sky130_fd_sc_hd__o221a_1
XFILLER_47_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16695_ _16707_/A vssd1 vssd1 vccd1 vccd1 _16695_/X sky130_fd_sc_hd__buf_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _18669_/D sky130_fd_sc_hd__clkbuf_1
X_18434_ _18434_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
X_12858_ _17642_/Q _12924_/A _12921_/A _17643_/Q _12857_/X vssd1 vssd1 vccd1 vccd1
+ _12858_/X sky130_fd_sc_hd__o221a_1
XFILLER_179_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11809_ _17783_/Q _11821_/B vssd1 vssd1 vccd1 vccd1 _11809_/Y sky130_fd_sc_hd__nor2_1
X_18365_ _18365_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
X_15577_ _15585_/B _15585_/C vssd1 vssd1 vccd1 vccd1 _15579_/B sky130_fd_sc_hd__nor2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12789_ _12761_/X _12789_/B vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__and2b_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17316_ _17765_/Q _19278_/Q _17381_/B vssd1 vssd1 vccd1 vccd1 _17317_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14476__636 _14476__636/A vssd1 vssd1 vccd1 vccd1 _18271_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18296_ _18296_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
X_14888__804 _14888__804/A vssd1 vssd1 vccd1 vccd1 _18449_/CLK sky130_fd_sc_hd__inv_2
X_17247_ _17250_/C _17246_/C _17250_/B vssd1 vssd1 vccd1 vccd1 _17248_/C sky130_fd_sc_hd__a21o_1
XFILLER_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03985_ _15767_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03985_/X sky130_fd_sc_hd__clkbuf_16
XPeripherals_171 vssd1 vssd1 vccd1 vccd1 Peripherals_171/HI io_oeb[34] sky130_fd_sc_hd__conb_1
XFILLER_190_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPeripherals_182 vssd1 vssd1 vccd1 vccd1 Peripherals_182/HI wb_data_o[21] sky130_fd_sc_hd__conb_1
XPeripherals_193 vssd1 vssd1 vccd1 vccd1 Peripherals_193/HI wb_error_o sky130_fd_sc_hd__conb_1
XFILLER_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17178_ _17179_/B _17180_/A _17177_/Y vssd1 vssd1 vccd1 vccd1 _19236_/D sky130_fd_sc_hd__a21oi_1
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16129_ _18625_/Q _18500_/Q _18906_/Q _18508_/Q _16127_/X _16128_/X vssd1 vssd1 vccd1
+ vccd1 _16129_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08951_ _08951_/A vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08882_ _08882_/A vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04368_ clkbuf_0__04368_/X vssd1 vssd1 vccd1 vccd1 _16314__214/A sky130_fd_sc_hd__clkbuf_16
XFILLER_229_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03419_ _14864_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03419_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09503_ _09503_/A vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09434_ _19048_/Q vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09365_ _19080_/Q _09096_/X _09369_/S vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09296_ _09296_/A vssd1 vssd1 vccd1 vccd1 _19114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789__724 _14789__724/A vssd1 vssd1 vccd1 vccd1 _18367_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10140_ _10155_/S vssd1 vssd1 vccd1 vccd1 _10149_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10071_ _10071_/A vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03974_ clkbuf_0__03974_/X vssd1 vssd1 vccd1 vccd1 _15716__1009/A sky130_fd_sc_hd__clkbuf_16
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106__412 _13106__412/A vssd1 vssd1 vccd1 vccd1 _17708_/CLK sky130_fd_sc_hd__inv_2
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13830_ _13830_/A _13855_/B _14053_/B vssd1 vssd1 vccd1 vccd1 _13847_/B sky130_fd_sc_hd__and3_1
X_17066__53 _17066__53/A vssd1 vssd1 vccd1 vccd1 _19202_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13761_ _13761_/A _13795_/B vssd1 vssd1 vccd1 vccd1 _13762_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_209 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _18288_/Q _09752_/X _10977_/S vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _17835_/Q _15505_/B vssd1 vssd1 vccd1 vccd1 _15501_/B sky130_fd_sc_hd__nand2_1
X_12712_ _12717_/C _12717_/D _12695_/X vssd1 vssd1 vccd1 vccd1 _12713_/B sky130_fd_sc_hd__o21ai_1
XFILLER_204_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _16480_/A _16480_/B vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__nor2_1
X_13692_ _13407_/X _13688_/X _13689_/X vssd1 vssd1 vccd1 vccd1 _13692_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_243_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _12383_/X _12640_/A _12617_/X vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__o21ai_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ _18150_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15362_ _15362_/A vssd1 vssd1 vccd1 vccd1 _15362_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ _18007_/Q _12574_/B _14067_/B _12574_/D vssd1 vssd1 vccd1 vccd1 _12574_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_180_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03408_ clkbuf_0__03408_/X vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__clkbuf_16
X_17101_ _17101_/A _17774_/Q _17101_/C vssd1 vssd1 vccd1 vccd1 _17101_/X sky130_fd_sc_hd__and3_1
XFILLER_184_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18081_ _19337_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_2
X_11525_ _18033_/Q _11341_/A hold24/A vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__mux2_1
X_15293_ _15301_/A vssd1 vssd1 vccd1 vccd1 _15293_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _14244_/A vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11456_ hold22/X _11456_/B _09025_/A vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__or3b_4
XFILLER_172_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ _15174_/B vssd1 vssd1 vccd1 vccd1 _10407_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11387_ _11387_/A vssd1 vssd1 vccd1 vccd1 _18122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ _13759_/A _13759_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _14113_/B sky130_fd_sc_hd__and3b_2
XFILLER_180_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _10338_/A vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__clkbuf_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _19013_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _17942_/Q _17696_/Q _13070_/S vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__mux2_1
X_17934_ _19136_/CLK _17934_/D vssd1 vssd1 vccd1 vccd1 _17934_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10269_ _10269_/A vssd1 vssd1 vccd1 vccd1 _18627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ _12007_/X _11975_/X _12008_/S vssd1 vssd1 vccd1 vccd1 _12008_/X sky130_fd_sc_hd__mux2_1
X_17865_ _17881_/CLK _17865_/D vssd1 vssd1 vccd1 vccd1 _17865_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16816_ _16811_/X _16814_/X _16984_/A vssd1 vssd1 vccd1 vccd1 _16816_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14482__640 _14484__642/A vssd1 vssd1 vccd1 vccd1 _18275_/CLK sky130_fd_sc_hd__inv_2
X_17796_ _19136_/CLK _17796_/D vssd1 vssd1 vccd1 vccd1 _17796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15847__148 _15848__149/A vssd1 vssd1 vccd1 vccd1 _18823_/CLK sky130_fd_sc_hd__inv_2
X_13959_ _13265_/X _13946_/X _13958_/Y _13951_/X vssd1 vssd1 vccd1 vccd1 _17964_/D
+ sky130_fd_sc_hd__a211oi_1
X_16747_ _19111_/Q _19110_/Q _17788_/Q vssd1 vssd1 vccd1 vccd1 _16748_/S sky130_fd_sc_hd__mux2_1
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18417_ _18417_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_1
X_15629_ _15626_/A _15622_/Y _15627_/X _15628_/X vssd1 vssd1 vccd1 vccd1 _18659_/D
+ sky130_fd_sc_hd__o211a_1
X_19397_ input28/X vssd1 vssd1 vccd1 vccd1 _19397_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09150_ _10869_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _09166_/S sky130_fd_sc_hd__nor2_2
XFILLER_188_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18348_ _18348_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18279_ _18279_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ hold12/X vssd1 vssd1 vccd1 vccd1 _10770_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput50 wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03968_ _15680_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03968_/X sky130_fd_sc_hd__clkbuf_16
Xinput61 wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput72 wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_8
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03799_ clkbuf_0__03799_/X vssd1 vssd1 vccd1 vccd1 _15429_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09983_ _09983_/A vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08934_ _08933_/X _19294_/Q _08942_/S vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08865_ _08887_/S vssd1 vssd1 vccd1 vccd1 _08878_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_111_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ _19344_/Q _08795_/X _08796_/S vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09417_ _09417_/A vssd1 vssd1 vccd1 vccd1 _19058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09348_ _19087_/Q _09268_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ _09279_/A vssd1 vssd1 vccd1 vccd1 _19121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11310_ _11310_/A vssd1 vssd1 vccd1 vccd1 _18152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12290_ _17562_/Q _18015_/Q _12293_/S vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ _11475_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11257_/S sky130_fd_sc_hd__or2_2
XFILLER_49_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11172_ _11147_/X _18209_/Q _11178_/S vssd1 vssd1 vccd1 vccd1 _11173_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _10123_/A vssd1 vssd1 vccd1 vccd1 _10123_/X sky130_fd_sc_hd__clkbuf_4
X_15980_ _15985_/B _15985_/C _15979_/Y vssd1 vssd1 vccd1 vccd1 _15980_/Y sky130_fd_sc_hd__o21ai_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _18459_/Q _14931_/B vssd1 vssd1 vccd1 vccd1 _14961_/D sky130_fd_sc_hd__xor2_1
X_10054_ _10117_/A vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17039__31 _17039__31/A vssd1 vssd1 vccd1 vccd1 _19180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _17991_/CLK _17650_/D vssd1 vssd1 vccd1 vccd1 _17650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _16613_/A _16601_/B _16601_/C vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__nor3_1
X_13813_ _13812_/X _13802_/X _13805_/X vssd1 vssd1 vccd1 vccd1 _13813_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17581_ _17581_/CLK _17581_/D vssd1 vssd1 vccd1 vccd1 _17581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15390__893 _15391__894/A vssd1 vssd1 vccd1 vccd1 _18580_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19320_ _19320_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
X_16532_ input71/X _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16533_/A sky130_fd_sc_hd__and3_1
X_13744_ _17891_/Q _13738_/X _13743_/Y _13741_/X vssd1 vssd1 vccd1 vccd1 _17891_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10956_ _10956_/A vssd1 vssd1 vccd1 vccd1 _18296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251_ _19251_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
X_16463_ _16466_/B _16440_/A _16462_/Y _16427_/X vssd1 vssd1 vccd1 vccd1 _16464_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13675_ _13240_/X _13666_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _13675_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_189_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ _18994_/Q vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__buf_4
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _18202_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _12626_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12631_/B sky130_fd_sc_hd__and2_1
X_14770__709 _14770__709/A vssd1 vssd1 vccd1 vccd1 _18352_/CLK sky130_fd_sc_hd__inv_2
X_19182_ _19182_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__04840_ clkbuf_0__04840_/X vssd1 vssd1 vccd1 vccd1 _17022__17/A sky130_fd_sc_hd__clkbuf_16
X_16394_ _18975_/Q vssd1 vssd1 vccd1 vccd1 _16466_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _18133_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _15345_/A vssd1 vssd1 vccd1 vccd1 _15345_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12557_ _12737_/C _12737_/B _12737_/A _12746_/C _12555_/X _12556_/X vssd1 vssd1 vccd1
+ vccd1 _12557_/X sky130_fd_sc_hd__mux4_2
XFILLER_157_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18064_ _18924_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
X_11508_ _11508_/A vssd1 vssd1 vccd1 vccd1 _18041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007__355 _17008__356/A vssd1 vssd1 vccd1 vccd1 _19154_/CLK sky130_fd_sc_hd__inv_2
X_15276_ _15271_/X _15272_/X _15274_/X _15275_/X _09600_/A _09625_/X vssd1 vssd1 vccd1
+ vccd1 _15276_/X sky130_fd_sc_hd__mux4_1
X_12488_ _17619_/Q vssd1 vssd1 vccd1 vccd1 _12706_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__07490_ clkbuf_0__07490_/X vssd1 vssd1 vccd1 vccd1 _12228__374/A sky130_fd_sc_hd__clkbuf_16
XFILLER_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14227_ _18084_/Q input42/X _14229_/S vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__mux2_1
X_11439_ _11454_/S vssd1 vssd1 vccd1 vccd1 _11448_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_153_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _14386_/A vssd1 vssd1 vccd1 vccd1 _14158_/X sky130_fd_sc_hd__buf_1
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15657__961 _15657__961/A vssd1 vssd1 vccd1 vccd1 _18678_/CLK sky130_fd_sc_hd__inv_2
X_13109_ _13109_/A vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__buf_1
X_18966_ _18966_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_1
X_14089_ _16516_/D vssd1 vssd1 vccd1 vccd1 _16052_/C sky130_fd_sc_hd__buf_6
XFILLER_113_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17917_ _17923_/CLK _17917_/D vssd1 vssd1 vccd1 vccd1 _17917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18897_ _18897_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17848_ _17850_/CLK _17848_/D vssd1 vssd1 vccd1 vccd1 _17848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14328__517 _14329__518/A vssd1 vssd1 vccd1 vccd1 _18152_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17779_ _17779_/CLK _17779_/D vssd1 vssd1 vccd1 vccd1 _17779_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_87_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18919_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_241_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04167_ _16092_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04167_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_wb_clk_i clkbuf_opt_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19128_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14859__780 _14862__783/A vssd1 vssd1 vccd1 vccd1 _18425_/CLK sky130_fd_sc_hd__inv_2
XFILLER_223_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17060__48 _17061__49/A vssd1 vssd1 vccd1 vccd1 _19197_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _19156_/Q _09145_/X _09202_/S vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _18665_/Q vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09064_ _09064_/A vssd1 vssd1 vccd1 vccd1 _19203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14489__646 _14490__647/A vssd1 vssd1 vccd1 vccd1 _18281_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09966_ _18473_/Q vssd1 vssd1 vccd1 vccd1 _10135_/A sky130_fd_sc_hd__buf_2
XFILLER_104_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08917_ _09679_/A vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__buf_2
XFILLER_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _11583_/B _11547_/A vssd1 vssd1 vccd1 vccd1 _09913_/S sky130_fd_sc_hd__nor2_2
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08848_ hold21/A _19046_/Q vssd1 vssd1 vccd1 vccd1 _09440_/A sky130_fd_sc_hd__or2b_1
XFILLER_100_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08779_ hold4/X vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _18364_/Q _10809_/X _10813_/S vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__08200_ clkbuf_0__08200_/X vssd1 vssd1 vccd1 vccd1 _13115__419/A sky130_fd_sc_hd__clkbuf_16
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _17826_/Q _11821_/B vssd1 vssd1 vccd1 vccd1 _11790_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _10741_/A vssd1 vssd1 vccd1 vccd1 _18392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13460_ _13623_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13484_/S sky130_fd_sc_hd__nor2_1
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10672_ _10752_/A hold8/X vssd1 vssd1 vccd1 vccd1 _10688_/S sky130_fd_sc_hd__nor2_2
XFILLER_41_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12411_ _12586_/S vssd1 vssd1 vccd1 vccd1 _12560_/S sky130_fd_sc_hd__buf_2
XFILLER_142_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13391_ _13623_/A vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__buf_4
X_15796__117 _15796__117/A vssd1 vssd1 vccd1 vccd1 _18789_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14433__601 _14434__602/A vssd1 vssd1 vccd1 vccd1 _18236_/CLK sky130_fd_sc_hd__inv_2
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _15060_/A _15060_/B _15060_/Y _14894_/Y vssd1 vssd1 vccd1 vccd1 _18471_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _12293_/S vssd1 vssd1 vccd1 vccd1 _12287_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14012_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11224_ _11239_/S vssd1 vssd1 vccd1 vccd1 _11233_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18820_ _18820_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ _11155_/A vssd1 vssd1 vccd1 vccd1 _18215_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10106_ _18721_/Q _10066_/X _10110_/S vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18751_ _18751_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ _11086_/A vssd1 vssd1 vccd1 vccd1 _18243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _15989_/A vssd1 vssd1 vccd1 vccd1 _15963_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _17951_/CLK _17702_/D vssd1 vssd1 vccd1 vccd1 _17702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14914_ _14914_/A _14914_/B vssd1 vssd1 vccd1 vccd1 _14963_/A sky130_fd_sc_hd__or2_1
X_10037_ _10037_/A vssd1 vssd1 vccd1 vccd1 _18748_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18682_ _18682_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17633_ _18012_/CLK _17633_/D vssd1 vssd1 vccd1 vccd1 _17633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17564_ _18027_/CLK _17564_/D vssd1 vssd1 vccd1 vccd1 _17564_/Q sky130_fd_sc_hd__dfxtp_2
X_11988_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12098_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19303_ _19303_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13727_ _17885_/Q _13715_/X _13724_/Y _13726_/X vssd1 vssd1 vccd1 vccd1 _17885_/D
+ sky130_fd_sc_hd__a211o_1
X_16515_ _14623_/A _16534_/B _16514_/Y _16364_/Y _18986_/Q vssd1 vssd1 vccd1 vccd1
+ _18986_/D sky130_fd_sc_hd__a32o_1
XFILLER_189_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10939_ _18303_/Q _10898_/X _10941_/S vssd1 vssd1 vccd1 vccd1 _10940_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17495_ _19338_/Q _12298_/X _12182_/X _19327_/Q _17494_/X vssd1 vssd1 vccd1 vccd1
+ _17495_/X sky130_fd_sc_hd__o221a_1
X_13119__422 _13120__423/A vssd1 vssd1 vccd1 vccd1 _17718_/CLK sky130_fd_sc_hd__inv_2
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19234_ _19251_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13658_ _13769_/A _13681_/B vssd1 vssd1 vccd1 vccd1 _13666_/A sky130_fd_sc_hd__nor2_2
X_16446_ _16467_/A _16446_/B _16453_/C vssd1 vssd1 vccd1 vccd1 _16446_/X sky130_fd_sc_hd__or3_1
XFILLER_220_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ _12610_/B _12610_/C _12608_/Y vssd1 vssd1 vccd1 vccd1 _17592_/D sky130_fd_sc_hd__a21oi_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19165_ _19165_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16377_ _17796_/Q _16383_/A _17795_/Q vssd1 vssd1 vccd1 vccd1 _16378_/B sky130_fd_sc_hd__o21ai_1
X_13589_ _17842_/Q _16520_/A _13589_/S vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15328_ _15328_/A vssd1 vssd1 vccd1 vccd1 _15328_/Y sky130_fd_sc_hd__inv_2
X_18116_ _18116_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19096_ _19096_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03805_ _15447_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03805_/X sky130_fd_sc_hd__clkbuf_16
X_15440__934 _15440__934/A vssd1 vssd1 vccd1 vccd1 _18621_/CLK sky130_fd_sc_hd__inv_2
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _15281_/A _15258_/Y _15305_/A vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__a21oi_1
X_18047_ _18047_/CLK _18047_/D vssd1 vssd1 vccd1 vccd1 _18047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _09691_/X _18822_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15397__899 _15397__899/A vssd1 vssd1 vccd1 vccd1 _18586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09751_ _09751_/A vssd1 vssd1 vccd1 vccd1 _18850_/D sky130_fd_sc_hd__clkbuf_1
X_18949_ _18949_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03598_ _15149_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03598_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _09682_/A vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_227_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15766__1049 _15766__1049/A vssd1 vssd1 vccd1 vccd1 _18766_/CLK sky130_fd_sc_hd__inv_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033__26 _17033__26/A vssd1 vssd1 vccd1 vccd1 _19175_/CLK sky130_fd_sc_hd__inv_2
XFILLER_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12341__401 _12342__402/A vssd1 vssd1 vccd1 vccd1 _17582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _10713_/A vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__buf_2
XFILLER_182_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__04010_ clkbuf_0__04010_/X vssd1 vssd1 vccd1 vccd1 _15860__159/A sky130_fd_sc_hd__clkbuf_16
XFILLER_198_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _11338_/A vssd1 vssd1 vccd1 vccd1 _09047_/X sky130_fd_sc_hd__buf_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16706__329 _16706__329/A vssd1 vssd1 vccd1 vccd1 _19104_/CLK sky130_fd_sc_hd__inv_2
XFILLER_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _18780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04843_ clkbuf_0__04843_/X vssd1 vssd1 vccd1 vccd1 _17039__31/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12960_/A vssd1 vssd1 vccd1 vccd1 _17673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_30 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_41 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_52 _13161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11911_ _17780_/Q vssd1 vssd1 vccd1 vccd1 _12067_/S sky130_fd_sc_hd__buf_2
XFILLER_219_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_63 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_74 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12891_ _17975_/Q _17661_/Q _12891_/S vssd1 vssd1 vccd1 vccd1 _12892_/B sky130_fd_sc_hd__mux2_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_85 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_96 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14628_/X _14629_/X _14734_/A vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11848_/A _11842_/B vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__and2_2
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _19049_/Q vssd1 vssd1 vccd1 vccd1 _14561_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11773_ _11773_/A vssd1 vssd1 vccd1 vccd1 _11773_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__buf_2
XFILLER_14_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03587_ clkbuf_0__03587_/X vssd1 vssd1 vccd1 vccd1 _15118_/A sky130_fd_sc_hd__clkbuf_16
X_16300_ _18995_/Q vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17280_ _17288_/C _17284_/C _17112_/B vssd1 vssd1 vccd1 vccd1 _17280_/Y sky130_fd_sc_hd__o21ai_1
X_10724_ _18399_/Q _10701_/X _10726_/S vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15804__124 _15804__124/A vssd1 vssd1 vccd1 vccd1 _18796_/CLK sky130_fd_sc_hd__inv_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16231_ _18629_/Q _18504_/Q _18910_/Q _18512_/Q _16182_/A _16117_/A vssd1 vssd1 vccd1
+ vccd1 _16231_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13443_ _13441_/X _13437_/X _13442_/Y _13213_/X vssd1 vssd1 vccd1 vccd1 _17795_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_201_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10655_ _10655_/A vssd1 vssd1 vccd1 vccd1 _18429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16162_ _16154_/X _16161_/X _16162_/S vssd1 vssd1 vccd1 vccd1 _16163_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13374_ _13374_/A vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__buf_4
XFILLER_126_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ _08991_/X _18491_/Q _10594_/S vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15044_ _15044_/A _15049_/B vssd1 vssd1 vccd1 vccd1 _15044_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04570_ _16639_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04570_/X sky130_fd_sc_hd__clkbuf_16
X_12256_ _17552_/Q _18025_/Q _12270_/S vssd1 vssd1 vccd1 vccd1 _12257_/B sky130_fd_sc_hd__mux2_1
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_1_1__f__03421_ clkbuf_0__03421_/X vssd1 vssd1 vccd1 vccd1 _14876__794/A sky130_fd_sc_hd__clkbuf_16
X_11207_ _11207_/A vssd1 vssd1 vccd1 vccd1 _18194_/D sky130_fd_sc_hd__clkbuf_1
X_12187_ _12187_/A vssd1 vssd1 vccd1 vccd1 _12187_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_214_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18803_ _18803_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ _18220_/Q _11062_/X _11140_/S vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16995_ _13830_/A input76/X _16997_/S vssd1 vssd1 vccd1 vccd1 _16996_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18734_ _18734_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _11223_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11085_/S sky130_fd_sc_hd__or2_2
X_15946_ _17814_/Q _15943_/B _17813_/Q vssd1 vssd1 vccd1 vccd1 _15947_/B sky130_fd_sc_hd__o21ai_1
XFILLER_237_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18665_ _14157_/A _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17616_ _17618_/CLK _17616_/D vssd1 vssd1 vccd1 vccd1 _17616_/Q sky130_fd_sc_hd__dfxtp_1
X_15173__879 _15173__879/A vssd1 vssd1 vccd1 vccd1 _18555_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18596_ _18596_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04004_ _15824_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04004_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_225_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17547_ _17547_/CLK _17547_/D vssd1 vssd1 vccd1 vccd1 _17547_/Q sky130_fd_sc_hd__dfxtp_1
X_14759_ _14759_/A vssd1 vssd1 vccd1 vccd1 _14759_/X sky130_fd_sc_hd__buf_1
X_16096__208 _16096__208/A vssd1 vssd1 vccd1 vccd1 _18913_/CLK sky130_fd_sc_hd__inv_2
XFILLER_225_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17478_ _19329_/Q _17478_/B vssd1 vssd1 vccd1 vccd1 _17485_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19217_ _19217_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16429_ _16475_/A vssd1 vssd1 vccd1 vccd1 _16429_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19148_ _19148_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04837_ _17006_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04837_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19079_ _19079_/CLK _19079_/D vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__07556_ _12326_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07556_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_246_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14783__719 _14783__719/A vssd1 vssd1 vccd1 vccd1 _18362_/CLK sky130_fd_sc_hd__inv_2
XFILLER_236_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03619_ clkbuf_0__03619_/X vssd1 vssd1 vccd1 vccd1 _15198__884/A sky130_fd_sc_hd__clkbuf_16
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _09734_/A vssd1 vssd1 vccd1 vccd1 _18856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19327_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09665_ _09665_/A vssd1 vssd1 vccd1 vccd1 _18910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09596_/A vssd1 vssd1 vccd1 vccd1 _18936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10440_ _10112_/X _18555_/Q _10448_/S vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10371_/A vssd1 vssd1 vccd1 vccd1 _18585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12110_ _12110_/A vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_123_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ _17700_/Q _13090_/B vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__xnor2_1
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _12115_/S vssd1 vssd1 vccd1 vccd1 _12111_/S sky130_fd_sc_hd__buf_2
XFILLER_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13992_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16780_ _16795_/A _16780_/B vssd1 vssd1 vccd1 vccd1 _19133_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12943_ _12931_/X _12933_/X _12942_/X _17669_/Q vssd1 vssd1 vccd1 vccd1 _12944_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18450_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
X_12874_ _17980_/Q _17656_/Q _12944_/B vssd1 vssd1 vccd1 vccd1 _12875_/B sky130_fd_sc_hd__mux2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15668_/A vssd1 vssd1 vccd1 vccd1 _15662_/X sky130_fd_sc_hd__buf_1
XFILLER_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12348__407 _12348__407/A vssd1 vssd1 vccd1 vccd1 _17588_/CLK sky130_fd_sc_hd__inv_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11825_ _19146_/Q vssd1 vssd1 vccd1 vccd1 _13830_/A sky130_fd_sc_hd__clkbuf_2
X_14613_ _17582_/Q _18380_/Q _18388_/Q _18422_/Q _14554_/X _09444_/A vssd1 vssd1 vccd1
+ vccd1 _14614_/B sky130_fd_sc_hd__mux4_1
X_15593_ _15591_/Y _15592_/Y _15581_/X vssd1 vssd1 vccd1 vccd1 _18652_/D sky130_fd_sc_hd__a21oi_1
X_18381_ _18381_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17332_ _17332_/A vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14544_/A vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11756_ _18000_/Q _17882_/Q vssd1 vssd1 vccd1 vccd1 _11757_/A sky130_fd_sc_hd__and2b_2
XFILLER_198_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03970_ clkbuf_0__03970_/X vssd1 vssd1 vccd1 vccd1 _15717_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10707_ _10707_/A vssd1 vssd1 vccd1 vccd1 _10707_/X sky130_fd_sc_hd__clkbuf_2
X_17263_ _17274_/D vssd1 vssd1 vccd1 vccd1 _17270_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11687_ _19033_/Q _16607_/B vssd1 vssd1 vccd1 vccd1 _16608_/B sky130_fd_sc_hd__and2_1
X_19002_ _19002_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_1
X_16214_ _16214_/A vssd1 vssd1 vccd1 vccd1 _16214_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13426_ _17792_/Q _13432_/S vssd1 vssd1 vccd1 vccd1 _13426_/Y sky130_fd_sc_hd__nor2_1
X_17194_ _19241_/Q _17194_/B vssd1 vssd1 vccd1 vccd1 _17203_/D sky130_fd_sc_hd__and2_1
X_10638_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10654_/S sky130_fd_sc_hd__or2_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886__367 _11886__367/A vssd1 vssd1 vccd1 vccd1 _17514_/CLK sky130_fd_sc_hd__inv_2
X_16145_ _18446_/Q _19084_/Q _19121_/Q _18430_/Q _16144_/X _10420_/X vssd1 vssd1 vccd1
+ vccd1 _16145_/X sky130_fd_sc_hd__mux4_2
X_13357_ _13357_/A vssd1 vssd1 vccd1 vccd1 _13375_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ _10569_/A vssd1 vssd1 vccd1 vccd1 _18498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12308_ _17552_/Q _12206_/X _12212_/A _17556_/Q _12307_/X vssd1 vssd1 vccd1 vccd1
+ _12308_/Y sky130_fd_sc_hd__a221oi_1
X_15765__1048 _15766__1049/A vssd1 vssd1 vccd1 vccd1 _18765_/CLK sky130_fd_sc_hd__inv_2
X_13288_ _13288_/A vssd1 vssd1 vccd1 vccd1 _13288_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14370__551 _14370__551/A vssd1 vssd1 vccd1 vccd1 _18186_/CLK sky130_fd_sc_hd__inv_2
X_15027_ _18464_/Q _14967_/X _15025_/X _15026_/X vssd1 vssd1 vccd1 vccd1 _15028_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03404_ clkbuf_0__03404_/X vssd1 vssd1 vccd1 vccd1 _14786__721/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__07172_ clkbuf_0__07172_/X vssd1 vssd1 vccd1 vccd1 _12222__369/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16978_ _18063_/Q _18055_/Q _18047_/Q _18039_/Q _16868_/A _16834_/X vssd1 vssd1 vccd1
+ vccd1 _16978_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 flash_io1_we vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
XFILLER_65_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18717_ _18717_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_1
X_15929_ _17822_/Q _15929_/B vssd1 vssd1 vccd1 vccd1 _15930_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09450_ _09446_/A _09453_/B _09449_/X vssd1 vssd1 vccd1 vccd1 _19049_/D sky130_fd_sc_hd__a21oi_1
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18648_ _18654_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03197_ clkbuf_0__03197_/X vssd1 vssd1 vccd1 vccd1 _14527__677/A sky130_fd_sc_hd__clkbuf_16
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09381_ _09381_/A vssd1 vssd1 vccd1 vccd1 _19074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18579_ _18579_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12225__371 _12226__372/A vssd1 vssd1 vccd1 vccd1 _17535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16629__271 _16632__274/A vssd1 vssd1 vccd1 vccd1 _19045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14271__471 _14271__471/A vssd1 vssd1 vccd1 vccd1 _18106_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03990_ clkbuf_0__03990_/X vssd1 vssd1 vccd1 vccd1 _15792__114/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17078__62 _17078__62/A vssd1 vssd1 vccd1 vccd1 _19211_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _18890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__or2_1
XFILLER_167_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09579_ _09579_/A vssd1 vssd1 vccd1 vccd1 _18943_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11610_ _11610_/A vssd1 vssd1 vccd1 vccd1 _17569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12590_ _12574_/B _14067_/B _14065_/B _12589_/X vssd1 vssd1 vccd1 vccd1 _12590_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03424_ clkbuf_0__03424_/X vssd1 vssd1 vccd1 vccd1 _14892__807/A sky130_fd_sc_hd__clkbuf_16
XFILLER_212_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11541_ _08880_/X _17714_/Q _11545_/S vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _11472_/A vssd1 vssd1 vccd1 vccd1 _18057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13211_ _13815_/A vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__buf_12
XFILLER_87_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10423_ _10423_/A vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__clkbuf_1
X_14191_ _14191_/A vssd1 vssd1 vccd1 vccd1 _18067_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _17723_/Q _13147_/B vssd1 vssd1 vccd1 vccd1 _13142_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _11565_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _10370_/S sky130_fd_sc_hd__nor2_2
XFILLER_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13073_ _17937_/Q _17701_/Q _13076_/S vssd1 vssd1 vccd1 vccd1 _13074_/B sky130_fd_sc_hd__mux2_1
X_17950_ _17951_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10285_ _10285_/A vssd1 vssd1 vccd1 vccd1 _18620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12024_ _11895_/X _11900_/X _12036_/S vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16901_ _16898_/X _16899_/X _16979_/S vssd1 vssd1 vccd1 vccd1 _16901_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17881_ _17881_/CLK _17881_/D vssd1 vssd1 vccd1 vccd1 _17881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16832_ _18179_/Q _18171_/Q _18163_/Q _18155_/Q _16813_/X _09869_/A vssd1 vssd1 vccd1
+ vccd1 _16833_/B sky130_fd_sc_hd__mux4_1
X_15651__956 _15651__956/A vssd1 vssd1 vccd1 vccd1 _18673_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ _16687_/B _16758_/Y _16761_/Y _13755_/A _16762_/X vssd1 vssd1 vccd1 vccd1
+ _16764_/B sky130_fd_sc_hd__o32a_1
X_13975_ _17970_/Q _13967_/X _13974_/Y vssd1 vssd1 vccd1 vccd1 _17970_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03151_ _14293_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03151_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18502_ _18502_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12926_ _17664_/Q _12835_/X _12834_/A _17654_/Q _12925_/X vssd1 vssd1 vccd1 vccd1
+ _12926_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_234_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18433_ _18433_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15645_ _15642_/X _15645_/B _16915_/A vssd1 vssd1 vccd1 vccd1 _15646_/A sky130_fd_sc_hd__and3b_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12857_ _17644_/Q _12920_/A _12835_/A _17647_/Q vssd1 vssd1 vccd1 vccd1 _12857_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ _17933_/Q _11785_/X _11800_/X _11807_/X vssd1 vssd1 vccd1 vccd1 _11808_/X
+ sky130_fd_sc_hd__o211a_4
X_18364_ _18364_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12788_ _17639_/Q _17996_/Q _12862_/B vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__mux2_1
X_15576_ _15573_/X _15575_/Y _15553_/X vssd1 vssd1 vccd1 vccd1 _18649_/D sky130_fd_sc_hd__a21oi_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17315_/A vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__clkbuf_1
X_11739_ _11739_/A vssd1 vssd1 vccd1 vccd1 _11739_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_230_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14853__775 _14853__775/A vssd1 vssd1 vccd1 vccd1 _18420_/CLK sky130_fd_sc_hd__inv_2
X_18295_ _18295_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17246_ _17250_/B _17250_/C _17246_/C vssd1 vssd1 vccd1 vccd1 _17252_/B sky130_fd_sc_hd__and3_1
Xclkbuf_0__03984_ _15761_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03984_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPeripherals_172 vssd1 vssd1 vccd1 vccd1 Peripherals_172/HI io_oeb[35] sky130_fd_sc_hd__conb_1
XPeripherals_183 vssd1 vssd1 vccd1 vccd1 Peripherals_183/HI wb_data_o[22] sky130_fd_sc_hd__conb_1
XFILLER_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPeripherals_194 vssd1 vssd1 vccd1 vccd1 io_oeb[0] Peripherals_194/LO sky130_fd_sc_hd__conb_1
X_13409_ _13407_/X _13395_/X _13408_/X vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__a21oi_1
X_17177_ _17179_/B _17180_/A _17126_/X vssd1 vssd1 vccd1 vccd1 _17177_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16128_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16128_/X sky130_fd_sc_hd__buf_2
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08950_ _19273_/Q _08949_/X _08959_/S vssd1 vssd1 vccd1 vccd1 _08951_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16059_ _16059_/A _16061_/B vssd1 vssd1 vccd1 vccd1 _18885_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08881_ _19310_/Q _08880_/X _08887_/S vssd1 vssd1 vccd1 vccd1 _08882_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04367_ clkbuf_0__04367_/X vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__03418_ _14858_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03418_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ _19006_/Q _09501_/X _09505_/S vssd1 vssd1 vccd1 vccd1 _09503_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09433_ _14544_/A vssd1 vssd1 vccd1 vccd1 _09433_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09364_/A vssd1 vssd1 vccd1 vccd1 _19081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09295_ _19114_/Q _08961_/X _09299_/S vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377__557 _14378__558/A vssd1 vssd1 vccd1 vccd1 _18192_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14754__695 _14758__699/A vssd1 vssd1 vccd1 vccd1 _18338_/CLK sky130_fd_sc_hd__inv_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput160 _11830_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10070_ _18736_/Q _10069_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__mux2_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03973_ clkbuf_0__03973_/X vssd1 vssd1 vccd1 vccd1 _15710__1004/A sky130_fd_sc_hd__clkbuf_16
XFILLER_88_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _13855_/B _16688_/B vssd1 vssd1 vccd1 vccd1 _13795_/B sky130_fd_sc_hd__nand2_2
X_10972_ _10972_/A vssd1 vssd1 vccd1 vccd1 _18289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12711_ _12717_/C _12717_/D vssd1 vssd1 vccd1 vccd1 _12713_/A sky130_fd_sc_hd__and2_1
XFILLER_243_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13691_ _17873_/Q _13682_/X _13690_/Y vssd1 vssd1 vccd1 vccd1 _17873_/D sky130_fd_sc_hd__o21a_1
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15764__1047 _15766__1049/A vssd1 vssd1 vccd1 vccd1 _18764_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12642_ _12651_/D vssd1 vssd1 vccd1 vccd1 _12647_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321__512 _14323__514/A vssd1 vssd1 vccd1 vccd1 _18147_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15361_ _19073_/Q _19065_/Q _19057_/Q _19011_/Q _15208_/A _09605_/A vssd1 vssd1 vccd1
+ vccd1 _15362_/A sky130_fd_sc_hd__mux4_1
X_15130__844 _15130__844/A vssd1 vssd1 vccd1 vccd1 _18520_/CLK sky130_fd_sc_hd__inv_2
XFILLER_212_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12573_ _18004_/Q _12834_/A _12470_/A vssd1 vssd1 vccd1 vccd1 _12574_/D sky130_fd_sc_hd__o21ba_1
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03407_ clkbuf_0__03407_/X vssd1 vssd1 vccd1 vccd1 _14806__738/A sky130_fd_sc_hd__clkbuf_16
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17100_ _13346_/B _17101_/C _17098_/Y _17099_/X vssd1 vssd1 vccd1 vccd1 _17100_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11524_ _11524_/A vssd1 vssd1 vccd1 vccd1 _18034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14312_ _14318_/A vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__buf_1
X_18080_ _19146_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
X_15292_ _19115_/Q _18946_/Q _18604_/Q _19344_/Q _15245_/X _15291_/X vssd1 vssd1 vccd1
+ vccd1 _15292_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113__417 _13115__419/A vssd1 vssd1 vccd1 vccd1 _17713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _17037_/A vssd1 vssd1 vccd1 vccd1 _17031_/X sky130_fd_sc_hd__buf_1
X_14278__477 _14280__479/A vssd1 vssd1 vccd1 vccd1 _18112_/CLK sky130_fd_sc_hd__inv_2
X_14243_ _14243_/A input65/X _14243_/C vssd1 vssd1 vccd1 vccd1 _14244_/A sky130_fd_sc_hd__and3_2
X_11455_ _11455_/A vssd1 vssd1 vccd1 vccd1 _18091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10406_ _10406_/A _10406_/B _10417_/A vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__and3_1
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ _11321_/X _18122_/Q _11394_/S vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ _18080_/Q vssd1 vssd1 vccd1 vccd1 _13759_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10337_ _18598_/Q _10336_/X _10343_/S vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18982_ _18987_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13076_/S vssd1 vssd1 vccd1 vccd1 _13070_/S sky130_fd_sc_hd__clkbuf_2
X_17933_ _19136_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _18627_/Q _10192_/X _10272_/S vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _19237_/Q _19238_/Q _12007_/S vssd1 vssd1 vccd1 vccd1 _12007_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17864_ _17881_/CLK _17864_/D vssd1 vssd1 vccd1 vccd1 _17864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10199_ _18687_/Q _10198_/X _10199_/S vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16815_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16984_/A sky130_fd_sc_hd__buf_2
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ _19014_/CLK _17795_/D vssd1 vssd1 vccd1 vccd1 _17795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16746_ _16741_/X _16743_/X _16786_/B vssd1 vssd1 vccd1 vccd1 _16746_/X sky130_fd_sc_hd__mux2_1
X_13958_ _17964_/Q _13962_/B vssd1 vssd1 vccd1 vccd1 _13958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_235_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12909_ _12894_/X _12909_/B vssd1 vssd1 vccd1 vccd1 _12910_/A sky130_fd_sc_hd__and2b_1
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16677_/X sky130_fd_sc_hd__buf_1
X_13889_ _17939_/Q _13878_/X _13888_/Y vssd1 vssd1 vccd1 vccd1 _17939_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18416_ _18416_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15628_ _16915_/A vssd1 vssd1 vccd1 vccd1 _15628_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ input31/X vssd1 vssd1 vccd1 vccd1 _19396_/X sky130_fd_sc_hd__buf_2
XFILLER_195_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18347_ _18347_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15559_ _18646_/Q _15569_/B vssd1 vssd1 vccd1 vccd1 _15559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09080_ _10690_/A vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__buf_2
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _18278_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17229_ _17229_/A vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__clkbuf_1
Xinput40 wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__03967_ _15674_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03967_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput51 wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_2
XFILLER_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput73 wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_8
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03798_ clkbuf_0__03798_/X vssd1 vssd1 vccd1 vccd1 _15413__912/A sky130_fd_sc_hd__clkbuf_16
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09982_ _18772_/Q _09947_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08933_ _09691_/A vssd1 vssd1 vccd1 vccd1 _08933_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08864_ _11529_/A _10851_/A vssd1 vssd1 vccd1 vccd1 _08887_/S sky130_fd_sc_hd__nor2_2
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _18883_/Q vssd1 vssd1 vccd1 vccd1 _08795_/X sky130_fd_sc_hd__buf_2
XFILLER_244_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__07169_ _11875_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07169_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09416_ _08910_/X _19058_/Q _09424_/S vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09347_ _09347_/A vssd1 vssd1 vccd1 vccd1 _19088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _19121_/Q _09277_/X _09281_/S vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ _11240_/A vssd1 vssd1 vccd1 vccd1 _18179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11171_ _11171_/A vssd1 vssd1 vccd1 vccd1 _18210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10122_/A vssd1 vssd1 vccd1 vccd1 _18716_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _14930_/A _14930_/B vssd1 vssd1 vccd1 vccd1 _14931_/B sky130_fd_sc_hd__nand2_1
X_10053_ _10053_/A vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804__736 _14807__739/A vssd1 vssd1 vccd1 vccd1 _18379_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _19028_/Q _16596_/B _19029_/Q vssd1 vssd1 vccd1 vccd1 _16601_/C sky130_fd_sc_hd__a21oi_1
XFILLER_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _13812_/A vssd1 vssd1 vccd1 vccd1 _13812_/X sky130_fd_sc_hd__buf_4
XFILLER_95_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17580_ _17580_/CLK _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16531_ _16531_/A vssd1 vssd1 vccd1 vccd1 _18993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13743_ _14074_/A _13743_/B vssd1 vssd1 vccd1 vccd1 _13743_/Y sky130_fd_sc_hd__nor2_1
X_10955_ _08871_/X _18296_/Q _10959_/S vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19250_ _19251_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16462_ _16466_/B _16466_/C vssd1 vssd1 vccd1 vccd1 _16462_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_177_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13674_ _13689_/A vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__clkbuf_2
X_10886_ _10886_/A vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18201_ _18201_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12625_ _12625_/A vssd1 vssd1 vccd1 vccd1 _17596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19181_ _19181_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16393_ _18975_/Q _16393_/B _16393_/C vssd1 vssd1 vccd1 vccd1 _16419_/B sky130_fd_sc_hd__and3_1
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _18132_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_1
X_12556_ _12556_/A vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15344_ _19072_/Q _19064_/Q _19056_/Q _19010_/Q _15232_/X _15233_/X vssd1 vssd1 vccd1
+ vccd1 _15345_/A sky130_fd_sc_hd__mux4_1
XFILLER_196_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ _18041_/Q _11341_/A _11509_/S vssd1 vssd1 vccd1 vccd1 _11508_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18063_ _18063_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
X_12487_ _12432_/X _12415_/X _12487_/S vssd1 vssd1 vccd1 vccd1 _12487_/X sky130_fd_sc_hd__mux2_2
X_15275_ _18937_/Q _18900_/Q _18892_/Q _18846_/Q _15251_/X _15252_/X vssd1 vssd1 vccd1
+ vccd1 _15275_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14226_ _14226_/A vssd1 vssd1 vccd1 vccd1 _18083_/D sky130_fd_sc_hd__clkbuf_1
X_11438_ _11511_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11454_/S sky130_fd_sc_hd__nor2_2
XFILLER_208_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14157_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14157_/X sky130_fd_sc_hd__buf_1
X_11369_ _11326_/X _18129_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _11370_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15853__153 _15854__154/A vssd1 vssd1 vccd1 vccd1 _18828_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14088_ _18013_/Q _14077_/S _14087_/Y vssd1 vssd1 vccd1 vccd1 _18013_/D sky130_fd_sc_hd__o21a_1
X_18965_ _18965_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13039_ _13076_/S vssd1 vssd1 vccd1 vccd1 _13053_/S sky130_fd_sc_hd__clkbuf_2
X_17916_ _19128_/CLK _17916_/D vssd1 vssd1 vccd1 vccd1 _17916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18896_ _18896_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17847_ _17850_/CLK _17847_/D vssd1 vssd1 vccd1 vccd1 _17847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17778_ _18021_/CLK _17778_/D vssd1 vssd1 vccd1 vccd1 _17778_/Q sky130_fd_sc_hd__dfxtp_1
X_17045__35 _17048__38/A vssd1 vssd1 vccd1 vccd1 _19184_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04166_ _16086_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04166_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_223_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09201_ _09201_/A vssd1 vssd1 vccd1 vccd1 _19157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15664__966 _15664__966/A vssd1 vssd1 vccd1 vccd1 _18683_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_56_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18010_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09132_ _09132_/A vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ _19203_/Q _08830_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _09064_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15763__1046 _15763__1046/A vssd1 vssd1 vccd1 vccd1 _18763_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09965_ _09965_/A vssd1 vssd1 vccd1 vccd1 _18776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08916_ _18886_/Q vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_246_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _09896_/A vssd1 vssd1 vccd1 vccd1 _18802_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _09446_/A hold12/A _08844_/A _08842_/Y vssd1 vssd1 vccd1 vccd1 _08847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_246_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ hold10/X vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10740_ _18392_/Q _10698_/X _10744_/S vssd1 vssd1 vccd1 vccd1 _10741_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _10671_/A vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12410_ _12515_/A vssd1 vssd1 vccd1 vccd1 _12586_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13390_ _11717_/X _13388_/Y _13389_/Y vssd1 vssd1 vccd1 vccd1 _17783_/D sky130_fd_sc_hd__o21a_1
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ _15060_/A _15060_/B vssd1 vssd1 vccd1 vccd1 _15060_/Y sky130_fd_sc_hd__nand2_1
X_12272_ _12272_/A vssd1 vssd1 vccd1 vccd1 _17556_/D sky130_fd_sc_hd__clkbuf_1
X_14810__740 _14814__744/A vssd1 vssd1 vccd1 vccd1 _18383_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11223_ _11223_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11239_/S sky130_fd_sc_hd__or2_2
XFILLER_181_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _11153_/X _18215_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ _10105_/A vssd1 vssd1 vccd1 vccd1 _18722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18750_ _18750_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11085_ _09055_/X _18243_/Q _11085_/S vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__mux2_1
X_15962_ _15962_/A vssd1 vssd1 vccd1 vccd1 _16025_/B sky130_fd_sc_hd__clkinv_2
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _17951_/CLK _17701_/D vssd1 vssd1 vccd1 vccd1 _17701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ _18467_/Q _14913_/B _14913_/C vssd1 vssd1 vccd1 vccd1 _14914_/B sky130_fd_sc_hd__and3_1
X_10036_ _18748_/Q _09947_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__mux2_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _18681_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17632_ _18012_/CLK _17632_/D vssd1 vssd1 vccd1 vccd1 _17632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17563_ _18021_/CLK _17563_/D vssd1 vssd1 vccd1 vccd1 _17563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11987_ _12109_/S vssd1 vssd1 vccd1 vccd1 _12037_/S sky130_fd_sc_hd__clkbuf_2
X_19302_ _19302_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16514_ _16514_/A _16534_/A _16514_/C vssd1 vssd1 vccd1 vccd1 _16514_/Y sky130_fd_sc_hd__nor3_1
X_13726_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13726_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17494_ _17494_/A _17494_/B _17494_/C _17494_/D vssd1 vssd1 vccd1 vccd1 _17494_/X
+ sky130_fd_sc_hd__and4_1
X_10938_ _10938_/A vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19233_ _19251_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _18971_/Q _16445_/B vssd1 vssd1 vccd1 vccd1 _16453_/C sky130_fd_sc_hd__and2_1
X_13657_ _17862_/Q _13649_/X _13656_/Y vssd1 vssd1 vccd1 vccd1 _17862_/D sky130_fd_sc_hd__o21a_1
X_10869_ _10869_/A _11547_/A vssd1 vssd1 vccd1 vccd1 _10885_/S sky130_fd_sc_hd__nor2_2
XFILLER_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12608_ _12610_/B _12610_/C _12607_/X vssd1 vssd1 vccd1 vccd1 _12608_/Y sky130_fd_sc_hd__o21ai_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _19164_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _18982_/Q _16376_/B vssd1 vssd1 vccd1 vccd1 _16376_/X sky130_fd_sc_hd__or2_1
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _17841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18115_ _18115_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _19071_/Q _19063_/Q _19055_/Q _19009_/Q _15232_/X _15233_/X vssd1 vssd1 vccd1
+ vccd1 _15328_/A sky130_fd_sc_hd__mux4_1
Xclkbuf_0__04853_ _17087_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04853_/X sky130_fd_sc_hd__clkbuf_16
X_12539_ _12568_/A _12539_/B vssd1 vssd1 vccd1 vccd1 _12539_/Y sky130_fd_sc_hd__nand2_1
X_19095_ _19095_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03804_ _15441_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03804_/X sky130_fd_sc_hd__clkbuf_16
X_18046_ _18046_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
X_15258_ _15258_/A vssd1 vssd1 vccd1 vccd1 _15258_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334__522 _14334__522/A vssd1 vssd1 vccd1 vccd1 _18157_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _14231_/A vssd1 vssd1 vccd1 vccd1 _14218_/S sky130_fd_sc_hd__buf_2
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15189_ _15626_/A _15186_/X _15188_/X _18660_/Q vssd1 vssd1 vccd1 vccd1 _15189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_103_wb_clk_i clkbuf_opt_1_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18924_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09750_ _18850_/Q _09749_/X _09759_/S vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__mux2_1
X_18948_ _18948_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03597_ _15143_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03597_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_227_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09681_ _09681_/A vssd1 vssd1 vccd1 vccd1 _18904_/D sky130_fd_sc_hd__clkbuf_1
X_18879_ _18879_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14495__651 _14498__654/A vssd1 vssd1 vccd1 vccd1 _18286_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09115_ _18987_/Q vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09046_ _18663_/Q vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_191_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09948_ _18780_/Q _09947_/X _09956_/S vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__04842_ clkbuf_0__04842_/X vssd1 vssd1 vccd1 vccd1 _17036__29/A sky130_fd_sc_hd__clkbuf_16
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_20 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_31 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09879_/A vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_42 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11910_ _17194_/B _19241_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_53 _13165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_64 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_75 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _12890_/A vssd1 vssd1 vccd1 vccd1 _17660_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_86 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__07492_ clkbuf_0__07492_/X vssd1 vssd1 vccd1 vccd1 _12239__383/A sky130_fd_sc_hd__clkbuf_16
XFILLER_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_97 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _17924_/Q _11839_/X _11840_/X _17905_/Q vssd1 vssd1 vccd1 vccd1 _11842_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11772_ _11772_/A input8/X vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__and2_4
XFILLER_199_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14560_ _14551_/X _14558_/X _14730_/S vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__mux2_2
XFILLER_54_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03586_ clkbuf_0__03586_/X vssd1 vssd1 vccd1 vccd1 _15416_/A sky130_fd_sc_hd__clkbuf_16
X_13511_ _17815_/Q _13499_/X _13510_/Y vssd1 vssd1 vccd1 vccd1 _17815_/D sky130_fd_sc_hd__o21a_1
X_10723_ _10723_/A vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _18779_/Q _18637_/Q _18787_/Q _18621_/Q _16117_/A _16138_/A vssd1 vssd1 vccd1
+ vccd1 _16230_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13442_ _17795_/Q _13444_/B vssd1 vssd1 vccd1 vccd1 _13442_/Y sky130_fd_sc_hd__nor2_1
X_10654_ _09280_/X _18429_/Q _10654_/S vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14396__571 _14396__571/A vssd1 vssd1 vccd1 vccd1 _18206_/CLK sky130_fd_sc_hd__inv_2
X_13373_ _11907_/S _13355_/X _13372_/Y _13359_/X vssd1 vssd1 vccd1 vccd1 _17779_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16161_ _16157_/X _16159_/X _16286_/S vssd1 vssd1 vccd1 vccd1 _16161_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ hold19/A vssd1 vssd1 vccd1 vccd1 _10594_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_166_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15112_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__buf_1
X_16092_ _16092_/A vssd1 vssd1 vccd1 vccd1 _16092_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18879_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12255_ _12293_/S vssd1 vssd1 vccd1 vccd1 _12270_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_181_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15043_ _18467_/Q _18466_/Q _15043_/C vssd1 vssd1 vccd1 vccd1 _15049_/B sky130_fd_sc_hd__and3_1
XFILLER_126_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _18194_/Q _11042_/X _11214_/S vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03420_ clkbuf_0__03420_/X vssd1 vssd1 vccd1 vccd1 _15086_/A sky130_fd_sc_hd__clkbuf_16
X_12186_ _12186_/A vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__buf_2
XFILLER_122_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18802_ _18802_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_1
X_11137_ _11137_/A vssd1 vssd1 vccd1 vccd1 _18221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16994_ _16994_/A vssd1 vssd1 vccd1 vccd1 _19145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18733_ _18733_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ _11222_/A _11068_/B _11383_/B vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__or3_2
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15945_ _15945_/A _15945_/B _15945_/C _15945_/D vssd1 vssd1 vccd1 vccd1 _15945_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _10019_/A vssd1 vssd1 vccd1 vccd1 _18756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18664_ _14157_/A _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17615_ _17618_/CLK _17615_/D vssd1 vssd1 vccd1 vccd1 _17615_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14827_ _14833_/A vssd1 vssd1 vccd1 vccd1 _14827_/X sky130_fd_sc_hd__buf_1
XFILLER_92_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18595_ _18595_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _17546_/CLK _17546_/D vssd1 vssd1 vccd1 vccd1 _17546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15762__1045 _15763__1046/A vssd1 vssd1 vccd1 vccd1 _18762_/CLK sky130_fd_sc_hd__inv_2
X_13709_ _13709_/A _13709_/B vssd1 vssd1 vccd1 vccd1 _13709_/Y sky130_fd_sc_hd__nor2_1
X_17477_ _19324_/Q _12180_/X _12298_/X _19338_/Q vssd1 vssd1 vccd1 vccd1 _17477_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14689_ _18368_/Q _18320_/Q _18376_/Q _17709_/Q _14599_/X _14627_/X vssd1 vssd1 vccd1
+ vccd1 _14689_/X sky130_fd_sc_hd__mux4_1
X_14817__746 _14818__747/A vssd1 vssd1 vccd1 vccd1 _18389_/CLK sky130_fd_sc_hd__inv_2
XFILLER_225_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19216_ _19216_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16428_ _16506_/A _16534_/A _16428_/C vssd1 vssd1 vccd1 vccd1 _16475_/A sky130_fd_sc_hd__and3_1
XFILLER_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19147_ _19147_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
X_16359_ _16359_/A vssd1 vssd1 vccd1 vccd1 _16359_/X sky130_fd_sc_hd__buf_1
XFILLER_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04836_ _17000_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04836_/X sky130_fd_sc_hd__clkbuf_16
X_19078_ _19078_/CLK _19078_/D vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18029_ _18029_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__07555_ _12320_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07555_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328__225 _16329__226/A vssd1 vssd1 vccd1 vccd1 _18941_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09802_ _18830_/Q _09761_/X _09806_/S vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09733_ _18856_/Q _09732_/X _09733_/S vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09664_ _18910_/Q _09268_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15866__163 _15867__164/A vssd1 vssd1 vccd1 vccd1 _18838_/CLK sky130_fd_sc_hd__inv_2
X_09595_ _18936_/Q _09501_/X _09597_/S vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19039_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_190 _09223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10370_ _18585_/Q _09741_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09029_ _09029_/A vssd1 vssd1 vccd1 vccd1 _19211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _12201_/A _12207_/A vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ _17976_/Q _13988_/X _13990_/Y vssd1 vssd1 vccd1 vccd1 _17976_/D sky130_fd_sc_hd__o21a_1
XFILLER_246_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _15730_/A vssd1 vssd1 vccd1 vccd1 _15730_/X sky130_fd_sc_hd__buf_1
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12942_ _12942_/A _12942_/B _12942_/C _12942_/D vssd1 vssd1 vccd1 vccd1 _12942_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_74_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__buf_1
XFILLER_234_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12873_ _12873_/A vssd1 vssd1 vccd1 vccd1 _17655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14662_/S vssd1 vssd1 vccd1 vccd1 _14679_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _17908_/Q _11812_/X _11821_/Y input17/X _11796_/X vssd1 vssd1 vccd1 vccd1
+ _11824_/X sky130_fd_sc_hd__a221o_2
X_18380_ _18380_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15595_/B _15597_/B vssd1 vssd1 vccd1 vccd1 _15592_/Y sky130_fd_sc_hd__nand2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17323_/X _17331_/B vssd1 vssd1 vccd1 vccd1 _17332_/A sky130_fd_sc_hd__and2b_1
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14543_/A vssd1 vssd1 vccd1 vccd1 _14543_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11755_ _11755_/A vssd1 vssd1 vccd1 vccd1 _11755_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17262_ _17264_/A _17262_/B _17262_/C _17262_/D vssd1 vssd1 vccd1 vccd1 _17274_/D
+ sky130_fd_sc_hd__and4_1
X_10706_ _10706_/A vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14474_ _14474_/A vssd1 vssd1 vccd1 vccd1 _14474_/X sky130_fd_sc_hd__buf_1
XFILLER_201_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11686_ _19032_/Q _19031_/Q _16602_/B vssd1 vssd1 vccd1 vccd1 _16607_/B sky130_fd_sc_hd__and3_1
X_19001_ _19001_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16213_ _16234_/A _16213_/B vssd1 vssd1 vccd1 vccd1 _16213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ _13425_/A vssd1 vssd1 vccd1 vccd1 _13709_/A sky130_fd_sc_hd__buf_4
X_17193_ _17194_/B _17195_/A _17192_/Y vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__a21oi_1
X_10637_ _10637_/A vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16144_ _16195_/A vssd1 vssd1 vccd1 vccd1 _16144_/X sky130_fd_sc_hd__clkbuf_4
X_13356_ _14072_/A vssd1 vssd1 vccd1 vccd1 _13740_/A sky130_fd_sc_hd__buf_4
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10568_ _10117_/X _18498_/Q _10574_/S vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _17563_/Q _12185_/A _12204_/A _17555_/Q vssd1 vssd1 vccd1 vccd1 _12307_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14138__424 _14138__424/A vssd1 vssd1 vccd1 vccd1 _18032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13287_ _17754_/Q _13280_/X _13286_/Y vssd1 vssd1 vccd1 vccd1 _17754_/D sky130_fd_sc_hd__o21a_1
X_10499_ _10499_/A vssd1 vssd1 vccd1 vccd1 _18529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _15026_/A vssd1 vssd1 vccd1 vccd1 _15026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03403_ clkbuf_0__03403_/X vssd1 vssd1 vccd1 vccd1 _14783__719/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _12169_/A vssd1 vssd1 vccd1 vccd1 _17527_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__07171_ clkbuf_0__07171_/X vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16977_ _19211_/Q _19163_/Q _18274_/Q _18266_/Q _16828_/A _16813_/X vssd1 vssd1 vccd1
+ vccd1 _16977_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14446__612 _14447__613/A vssd1 vssd1 vccd1 vccd1 _18247_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 flash_io1_write vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18716_ _18716_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_1
X_15928_ _15967_/C _15926_/Y _15927_/X vssd1 vssd1 vccd1 vccd1 _15928_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_209_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18647_ _18657_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03196_ clkbuf_0__03196_/X vssd1 vssd1 vccd1 vccd1 _14523__674/A sky130_fd_sc_hd__clkbuf_16
XFILLER_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09380_ _19074_/Q _08944_/X _09388_/S vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18578_ _18578_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17529_ _18031_/CLK _17529_/D vssd1 vssd1 vccd1 vccd1 _17529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17499__6 _17501__8/A vssd1 vssd1 vccd1 vccd1 _19341_/CLK sky130_fd_sc_hd__inv_2
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09716_ _09697_/X _18890_/Q _09716_/S vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _18926_/D sky130_fd_sc_hd__nor2_1
XFILLER_216_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09578_ _18943_/Q _09504_/X _09578_/S vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__mux2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03423_ clkbuf_0__03423_/X vssd1 vssd1 vccd1 vccd1 _14888__804/A sky130_fd_sc_hd__clkbuf_16
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17396__89 _17396__89/A vssd1 vssd1 vccd1 vccd1 _19302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11540_ _11540_/A vssd1 vssd1 vccd1 vccd1 _17715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _11341_/X _18057_/Q _11473_/S vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ input55/X _13210_/B vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__nand2_4
X_10422_ _10405_/B _10422_/B _10433_/C vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__and3b_1
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15460__949 _15460__949/A vssd1 vssd1 vccd1 vccd1 _18636_/CLK sky130_fd_sc_hd__inv_2
XFILLER_167_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14190_ _13873_/A input47/X _14196_/S vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13141_ _14136_/B vssd1 vssd1 vccd1 vccd1 _13147_/B sky130_fd_sc_hd__clkbuf_2
X_10353_ _10353_/A vssd1 vssd1 vccd1 vccd1 _18593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _13072_/A vssd1 vssd1 vccd1 vccd1 _17700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10284_ _18620_/Q _10189_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10285_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12023_ _11916_/X _11892_/X _12032_/S vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16900_ _16900_/A vssd1 vssd1 vccd1 vccd1 _16979_/S sky130_fd_sc_hd__clkbuf_2
X_17880_ _17881_/CLK _17880_/D vssd1 vssd1 vccd1 vccd1 _17880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16831_ _16900_/A vssd1 vssd1 vccd1 vccd1 _16929_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16762_ _16762_/A vssd1 vssd1 vccd1 vccd1 _16762_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13974_ _13777_/X _13973_/X _13920_/X vssd1 vssd1 vccd1 vccd1 _13974_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03150_ _14287_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03150_/X sky130_fd_sc_hd__clkbuf_16
X_18501_ _18501_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12925_ _17655_/Q _13081_/B vssd1 vssd1 vccd1 vccd1 _12925_/X sky130_fd_sc_hd__xor2_1
XFILLER_246_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18432_ _18432_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15644_ _15642_/B _15619_/X _16860_/A _15642_/A vssd1 vssd1 vccd1 vccd1 _15645_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _17638_/Q _13081_/B vssd1 vssd1 vccd1 vccd1 _12859_/C sky130_fd_sc_hd__xor2_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _17914_/Q _11793_/X _11806_/X _11802_/X vssd1 vssd1 vccd1 vccd1 _11807_/X
+ sky130_fd_sc_hd__a211o_1
X_18363_ _18363_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15575_ _18649_/Q _15597_/B vssd1 vssd1 vccd1 vccd1 _15575_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12787_ _12787_/A vssd1 vssd1 vccd1 vccd1 _17638_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17314_ _17304_/X _17314_/B vssd1 vssd1 vccd1 vccd1 _17315_/A sky130_fd_sc_hd__and2b_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11738_ _17934_/Q _11742_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__and2_4
X_18294_ _18294_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ _17250_/C _17246_/C _17244_/Y vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__a21oi_1
XFILLER_187_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03983_ _15755_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03983_/X sky130_fd_sc_hd__clkbuf_16
X_11669_ _17508_/Q _09694_/A _11671_/S vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__mux2_1
XPeripherals_173 vssd1 vssd1 vccd1 vccd1 Peripherals_173/HI io_oeb[36] sky130_fd_sc_hd__conb_1
XFILLER_70_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13408_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17176_ _17180_/A _17176_/B vssd1 vssd1 vccd1 vccd1 _19235_/D sky130_fd_sc_hd__nor2_1
XPeripherals_184 vssd1 vssd1 vccd1 vccd1 Peripherals_184/HI wb_data_o[23] sky130_fd_sc_hd__conb_1
XFILLER_122_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPeripherals_195 vssd1 vssd1 vccd1 vccd1 io_oeb[2] Peripherals_195/LO sky130_fd_sc_hd__conb_1
XFILLER_155_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14388_ _14400_/A vssd1 vssd1 vccd1 vccd1 _14388_/X sky130_fd_sc_hd__buf_1
XFILLER_127_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16127_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16127_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13339_ _17772_/Q _13329_/X _13338_/Y vssd1 vssd1 vccd1 vccd1 _17772_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ _16058_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _18884_/D sky130_fd_sc_hd__nor2_1
XFILLER_233_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15009_ _15009_/A vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__clkbuf_1
X_08880_ _18989_/Q vssd1 vssd1 vccd1 vccd1 _08880_/X sky130_fd_sc_hd__buf_6
XFILLER_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03417_ _14852_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03417_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_244_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09501_ _18881_/Q vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__buf_2
XFILLER_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ _19050_/Q vssd1 vssd1 vccd1 vccd1 _14544_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_240_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03179_ clkbuf_0__03179_/X vssd1 vssd1 vccd1 vccd1 _14436__604/A sky130_fd_sc_hd__clkbuf_16
XFILLER_197_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _19081_/Q _09092_/X _09369_/S vssd1 vssd1 vccd1 vccd1 _09364_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09294_ _09294_/A vssd1 vssd1 vccd1 vccd1 _19115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput150 _11860_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_134_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput161 _11833_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_133_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17302__78 _17302__78/A vssd1 vssd1 vccd1 vccd1 _19274_/CLK sky130_fd_sc_hd__inv_2
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03972_ clkbuf_0__03972_/X vssd1 vssd1 vccd1 vccd1 _15701__996/A sky130_fd_sc_hd__clkbuf_16
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _18289_/Q _09749_/X _10977_/S vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12710_ _12710_/A vssd1 vssd1 vccd1 vccd1 _17620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13690_ _13529_/X _13688_/X _13689_/X vssd1 vssd1 vccd1 vccd1 _13690_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_204_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12641_ _17601_/Q _17600_/Q _17599_/Q _12641_/D vssd1 vssd1 vccd1 vccd1 _12651_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _19218_/Q _19106_/Q _18289_/Q _19098_/Q _15308_/X _09613_/A vssd1 vssd1 vccd1
+ vccd1 _15360_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12572_ _12774_/D vssd1 vssd1 vccd1 vccd1 _12834_/A sky130_fd_sc_hd__buf_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03406_ clkbuf_0__03406_/X vssd1 vssd1 vccd1 vccd1 _14801__734/A sky130_fd_sc_hd__clkbuf_16
XFILLER_212_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11523_ _18034_/Q _11338_/A hold24/A vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15291_ _15291_/A vssd1 vssd1 vccd1 vccd1 _15291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _15076_/A _14241_/X _18482_/Q vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11454_ _18091_/Q _11282_/X _11454_/S vssd1 vssd1 vccd1 vccd1 _11455_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10405_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10417_/A sky130_fd_sc_hd__and2_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11385_ _11400_/S vssd1 vssd1 vccd1 vccd1 _11394_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03199_ clkbuf_0__03199_/X vssd1 vssd1 vccd1 vccd1 _14539__687/A sky130_fd_sc_hd__clkbuf_16
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13124_ _13845_/A _11707_/S _16715_/B vssd1 vssd1 vccd1 vccd1 _17722_/D sky130_fd_sc_hd__a21o_1
X_10336_ _18478_/Q vssd1 vssd1 vccd1 vccd1 _10336_/X sky130_fd_sc_hd__clkbuf_4
X_18981_ _19014_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13055_ _13055_/A vssd1 vssd1 vccd1 vccd1 _17695_/D sky130_fd_sc_hd__clkbuf_1
X_17932_ _19136_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10267_/A vssd1 vssd1 vccd1 vccd1 _18628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12006_ _19233_/Q _17173_/B _19235_/Q _19236_/Q _11924_/S _12008_/S vssd1 vssd1 vccd1
+ vccd1 _12006_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17863_ _17881_/CLK _17863_/D vssd1 vssd1 vccd1 vccd1 _17863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ _18473_/Q vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__buf_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319__384 _12319__384/A vssd1 vssd1 vccd1 vccd1 _17565_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16814_ _19204_/Q _19156_/Q _18267_/Q _18259_/Q _16828_/A _16813_/X vssd1 vssd1 vccd1
+ vccd1 _16814_/X sky130_fd_sc_hd__mux4_1
X_17794_ _19135_/CLK _17794_/D vssd1 vssd1 vccd1 vccd1 _17794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16745_ _19110_/Q _17788_/Q _16744_/X vssd1 vssd1 vccd1 vccd1 _16786_/B sky130_fd_sc_hd__o21a_2
X_13957_ _13192_/X _13946_/X _13956_/Y _13951_/X vssd1 vssd1 vccd1 vccd1 _17963_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12908_ _17970_/Q _17666_/Q _12908_/S vssd1 vssd1 vccd1 vccd1 _12909_/B sky130_fd_sc_hd__mux2_1
X_17072__58 _17073__59/A vssd1 vssd1 vccd1 vccd1 _19207_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16676_ _16718_/A vssd1 vssd1 vccd1 vccd1 _16676_/X sky130_fd_sc_hd__buf_1
X_13888_ _13669_/X _13885_/X _13880_/X vssd1 vssd1 vccd1 vccd1 _13888_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15627_ _15535_/A _15630_/B _15626_/X _15622_/B _15642_/A vssd1 vssd1 vccd1 vccd1
+ _15627_/X sky130_fd_sc_hd__a311o_1
X_18415_ _18415_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
X_19395_ input25/X vssd1 vssd1 vccd1 vccd1 _19395_/X sky130_fd_sc_hd__clkbuf_1
X_12839_ _17651_/Q _12838_/X _12834_/X _17637_/Q vssd1 vssd1 vccd1 vccd1 _12843_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18346_ _18346_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15558_ _15579_/A _15558_/B _15561_/B vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__or3_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18277_ _18277_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _17830_/Q _15489_/B vssd1 vssd1 vccd1 vccd1 _15490_/B sky130_fd_sc_hd__xor2_1
X_17228_ _17233_/C _17235_/B _17228_/C vssd1 vssd1 vccd1 vccd1 _17229_/A sky130_fd_sc_hd__and3b_1
Xinput30 vga_r[1] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__03966_ _15668_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03966_/X sky130_fd_sc_hd__clkbuf_16
Xinput41 wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput52 wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
XFILLER_238_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput63 wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17159_ _17159_/A _17159_/B vssd1 vssd1 vccd1 vccd1 _17160_/C sky130_fd_sc_hd__or2_1
XFILLER_128_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput74 wb_rst_i vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_6
Xclkbuf_1_1__f__03797_ clkbuf_0__03797_/X vssd1 vssd1 vccd1 vccd1 _15409__909/A sky130_fd_sc_hd__clkbuf_16
XFILLER_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15107__825 _15109__827/A vssd1 vssd1 vccd1 vccd1 _18501_/CLK sky130_fd_sc_hd__inv_2
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _09981_/A vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08932_ _18882_/Q vssd1 vssd1 vccd1 vccd1 _09691_/A sky130_fd_sc_hd__buf_2
XFILLER_233_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08863_ _10931_/A vssd1 vssd1 vccd1 vccd1 _10851_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08794_ _08794_/A vssd1 vssd1 vccd1 vccd1 _19345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__07168_ _11874_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07168_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14383__562 _14385__564/A vssd1 vssd1 vccd1 vccd1 _18197_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09415_ _09430_/S vssd1 vssd1 vccd1 vccd1 _09424_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09346_ _19088_/Q _09265_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _09347_/A sky130_fd_sc_hd__mux2_1
X_14459__622 _14460__623/A vssd1 vssd1 vccd1 vccd1 _18257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_200_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09277_ _18474_/Q vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__buf_2
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14390__566 _14391__567/A vssd1 vssd1 vccd1 vccd1 _18201_/CLK sky130_fd_sc_hd__inv_2
X_11170_ _11142_/X _18210_/Q _11178_/S vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10121_ _10120_/X _18716_/Q _10127_/S vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ _18742_/Q _10048_/X _10064_/S vssd1 vssd1 vccd1 vccd1 _10053_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238__382 _12239__383/A vssd1 vssd1 vccd1 vccd1 _17546_/CLK sky130_fd_sc_hd__inv_2
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _17914_/Q _13797_/X _13810_/Y vssd1 vssd1 vccd1 vccd1 _17914_/D sky130_fd_sc_hd__o21a_1
XFILLER_217_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _16530_/A _16530_/B vssd1 vssd1 vccd1 vccd1 _16531_/A sky130_fd_sc_hd__and2_1
XFILLER_232_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13742_ _17890_/Q _13738_/X _13740_/Y _13741_/X vssd1 vssd1 vccd1 vccd1 _17890_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10954_ _10954_/A vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14284__482 _14284__482/A vssd1 vssd1 vccd1 vccd1 _18117_/CLK sky130_fd_sc_hd__inv_2
XFILLER_244_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _16459_/X _16460_/Y _16480_/A vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__a21oi_1
X_13673_ _17867_/Q _13659_/X _13672_/Y vssd1 vssd1 vccd1 vccd1 _17867_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ _18331_/Q _10812_/X _10885_/S vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18200_ _18200_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12624_ _12626_/B _12624_/B _12695_/A vssd1 vssd1 vccd1 vccd1 _12625_/A sky130_fd_sc_hd__and3b_1
X_19180_ _19180_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16392_ _17801_/Q _16397_/B vssd1 vssd1 vccd1 vccd1 _16393_/C sky130_fd_sc_hd__nand2_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17505__3 _17506__4/A vssd1 vssd1 vccd1 vccd1 _19347_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18131_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15343_ _19217_/Q _19105_/Q _18288_/Q _19097_/Q _15308_/X _09613_/A vssd1 vssd1 vccd1
+ vccd1 _15343_/X sky130_fd_sc_hd__mux4_1
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _12555_/A vssd1 vssd1 vccd1 vccd1 _12555_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04369_ clkbuf_0__04369_/X vssd1 vssd1 vccd1 vccd1 _16320__219/A sky130_fd_sc_hd__clkbuf_16
XFILLER_145_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11506_ _11506_/A vssd1 vssd1 vccd1 vccd1 _18042_/D sky130_fd_sc_hd__clkbuf_1
X_18062_ _18062_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
X_15274_ _19318_/Q _19302_/Q _19294_/Q _19269_/Q _15273_/X _15249_/X vssd1 vssd1 vccd1
+ vccd1 _15274_/X sky130_fd_sc_hd__mux4_1
X_12486_ _12428_/X _12431_/X _12487_/S vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__mux2_2
XFILLER_157_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _17013_/X sky130_fd_sc_hd__buf_1
XFILLER_156_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14225_ _18083_/Q input41/X _14229_/S vssd1 vssd1 vccd1 vccd1 _14226_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ _11437_/A vssd1 vssd1 vccd1 vccd1 _18099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15892__181 _15893__182/A vssd1 vssd1 vccd1 vccd1 _18857_/CLK sky130_fd_sc_hd__inv_2
X_11368_ _11368_/A vssd1 vssd1 vccd1 vccd1 _18130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10319_ _10319_/A vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14087_ _13815_/X _14077_/S _14060_/X vssd1 vssd1 vccd1 vccd1 _14087_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18964_ _18964_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_1
X_11299_ _18156_/Q _11279_/X _11301_/S vssd1 vssd1 vccd1 vccd1 _11300_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13038_ _13038_/A vssd1 vssd1 vccd1 vccd1 _17690_/D sky130_fd_sc_hd__clkbuf_1
X_17915_ _19128_/CLK _17915_/D vssd1 vssd1 vccd1 vccd1 _17915_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _18895_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17846_ _17850_/CLK _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17777_ _18021_/CLK _17777_/D vssd1 vssd1 vccd1 vccd1 _17777_/Q sky130_fd_sc_hd__dfxtp_1
X_14989_ _15001_/A _14989_/B vssd1 vssd1 vccd1 vccd1 _14990_/A sky130_fd_sc_hd__and2_1
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04165_ _16080_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04165_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_235_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09200_ _19157_/Q _09142_/X _09202_/S vssd1 vssd1 vccd1 vccd1 _09201_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ _19185_/Q _09130_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09132_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18329_ _18996_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _09077_/S vssd1 vssd1 vccd1 vccd1 _09071_/S sky130_fd_sc_hd__buf_2
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_96_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _15785_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19147_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14866__786 _14866__786/A vssd1 vssd1 vccd1 vccd1 _18431_/CLK sky130_fd_sc_hd__inv_2
X_09964_ _18776_/Q _09963_/X _09968_/S vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08915_ _08915_/A vssd1 vssd1 vccd1 vccd1 _19299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _09891_/B _09895_/B _09895_/C vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__and3b_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _08838_/A _09442_/A _09441_/A _09441_/B vssd1 vssd1 vccd1 vccd1 _08846_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _11655_/A vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__buf_4
XFILLER_100_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _18421_/Q _09741_/X _10670_/S vssd1 vssd1 vccd1 vccd1 _10671_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09329_/A vssd1 vssd1 vccd1 vccd1 _19096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12271_ _12263_/X _12271_/B vssd1 vssd1 vccd1 vccd1 _12272_/A sky130_fd_sc_hd__and2b_1
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14010_ _14090_/A _14031_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__and3_2
X_11222_ _11222_/A _11456_/B _11383_/B vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__or3_4
XFILLER_175_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ _11332_/A vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10104_ _18722_/Q _10063_/X _10104_/S vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__mux2_1
X_11084_ _11084_/A vssd1 vssd1 vccd1 vccd1 _18244_/D sky130_fd_sc_hd__clkbuf_1
X_15961_ _16033_/A _15961_/B vssd1 vssd1 vccd1 vccd1 _18861_/D sky130_fd_sc_hd__nor2_1
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17700_ _17951_/CLK _17700_/D vssd1 vssd1 vccd1 vccd1 _17700_/Q sky130_fd_sc_hd__dfxtp_1
X_14912_ _14913_/B _14913_/C _18467_/Q vssd1 vssd1 vccd1 vccd1 _14914_/A sky130_fd_sc_hd__a21oi_1
X_10035_ _10035_/A vssd1 vssd1 vccd1 vccd1 _18749_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18680_ _18680_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17631_ _18012_/CLK _17631_/D vssd1 vssd1 vccd1 vccd1 _17631_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17562_ _18021_/CLK _17562_/D vssd1 vssd1 vccd1 vccd1 _17562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11986_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12109_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440__607 _14440__607/A vssd1 vssd1 vccd1 vccd1 _18242_/CLK sky130_fd_sc_hd__inv_2
XFILLER_189_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19301_ _19301_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
X_16513_ _16511_/A _16505_/X _16512_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18985_/D
+ sky130_fd_sc_hd__o211a_1
X_13725_ _17454_/A vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__buf_2
X_17493_ _17493_/A _17493_/B _17493_/C _17493_/D vssd1 vssd1 vccd1 vccd1 _17494_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_56_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10937_ _18304_/Q _10895_/X _10941_/S vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19232_ _19251_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _18971_/Q _16445_/B vssd1 vssd1 vccd1 vccd1 _16446_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13656_ _13712_/A _13649_/A _13532_/X vssd1 vssd1 vccd1 vccd1 _13656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_204_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ _10868_/A vssd1 vssd1 vccd1 vccd1 _18339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _19163_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _18982_/Q _16376_/B vssd1 vssd1 vccd1 vccd1 _16375_/Y sky130_fd_sc_hd__nand2_1
X_13587_ _13629_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__or2_1
XFILLER_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10799_ _10799_/A vssd1 vssd1 vccd1 vccd1 _18368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18114_ _18114_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__04852_ _17081_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04852_/X sky130_fd_sc_hd__clkbuf_16
X_15326_ _19216_/Q _19104_/Q _18287_/Q _19096_/Q _15308_/X _09631_/X vssd1 vssd1 vccd1
+ vccd1 _15326_/X sky130_fd_sc_hd__mux4_1
X_12538_ _12538_/A vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__clkbuf_2
X_19094_ _19094_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03803_ _15435_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03803_/X sky130_fd_sc_hd__clkbuf_16
X_18045_ _18045_/CLK _18045_/D vssd1 vssd1 vccd1 vccd1 _18045_/Q sky130_fd_sc_hd__dfxtp_1
X_15257_ _19068_/Q _19060_/Q _19052_/Q _19006_/Q _15208_/A _09605_/A vssd1 vssd1 vccd1
+ vccd1 _15258_/A sky130_fd_sc_hd__mux4_1
X_12469_ _12462_/X _12467_/X _12469_/S vssd1 vssd1 vccd1 vccd1 _12470_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _14208_/A vssd1 vssd1 vccd1 vccd1 _18075_/D sky130_fd_sc_hd__clkbuf_1
X_15188_ _15188_/A _18659_/Q vssd1 vssd1 vccd1 vccd1 _15188_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ _14151_/A vssd1 vssd1 vccd1 vccd1 _14139_/X sky130_fd_sc_hd__buf_1
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03596_ _15137_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03596_/X sky130_fd_sc_hd__clkbuf_16
X_18947_ _18947_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09680_ _09679_/X _18904_/Q _09689_/S vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__mux2_1
X_15670__971 _15671__972/A vssd1 vssd1 vccd1 vccd1 _18688_/CLK sky130_fd_sc_hd__inv_2
X_18878_ _18888_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17018__14 _17018__14/A vssd1 vssd1 vccd1 vccd1 _19163_/CLK sky130_fd_sc_hd__inv_2
X_17829_ _18919_/CLK _17829_/D vssd1 vssd1 vccd1 vccd1 _17829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14872__790 _14873__791/A vssd1 vssd1 vccd1 vccd1 _18435_/CLK sky130_fd_sc_hd__inv_2
XFILLER_241_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ _09114_/A vssd1 vssd1 vccd1 vccd1 _19189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09045_ _09045_/A vssd1 vssd1 vccd1 vccd1 _19207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16999__349 _16999__349/A vssd1 vssd1 vccd1 vccd1 _19148_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09947_ _10120_/A vssd1 vssd1 vccd1 vccd1 _09947_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__04841_ clkbuf_0__04841_/X vssd1 vssd1 vccd1 vccd1 _17028__22/A sky130_fd_sc_hd__clkbuf_16
XFILLER_213_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_10 _10180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09878_/A vssd1 vssd1 vccd1 vccd1 _18807_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07560_ clkbuf_0__07560_/X vssd1 vssd1 vccd1 vccd1 _13102__409/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_32 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_43 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_54 _13265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _08829_/A vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_65 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_76 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__07491_ clkbuf_0__07491_/X vssd1 vssd1 vccd1 vccd1 _12234__379/A sky130_fd_sc_hd__clkbuf_16
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_87 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_98 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11840_ _11840_/A vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504__659 _14504__659/A vssd1 vssd1 vccd1 vccd1 _18294_/CLK sky130_fd_sc_hd__inv_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_242_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13510_ _13237_/X _13499_/A _13494_/X vssd1 vssd1 vccd1 vccd1 _13510_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03585_ clkbuf_0__03585_/X vssd1 vssd1 vccd1 vccd1 _15089__812/A sky130_fd_sc_hd__clkbuf_16
XFILLER_241_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ _18400_/Q _10698_/X _10726_/S vssd1 vssd1 vccd1 vccd1 _10723_/A sky130_fd_sc_hd__mux2_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13441_ _13441_/A vssd1 vssd1 vccd1 vccd1 _13441_/X sky130_fd_sc_hd__buf_6
X_10653_ _10653_/A vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16160_ _16289_/S vssd1 vssd1 vccd1 vccd1 _16286_/S sky130_fd_sc_hd__clkbuf_2
X_13372_ _13750_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _13372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ hold18/X _11365_/B vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__or2_2
XFILLER_220_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15042_ _18467_/Q _15042_/B vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12254_ _12254_/A vssd1 vssd1 vccd1 vccd1 _17551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ _11220_/S vssd1 vssd1 vccd1 vccd1 _11214_/S sky130_fd_sc_hd__clkbuf_2
X_12185_ _12185_/A vssd1 vssd1 vccd1 vccd1 _12185_/X sky130_fd_sc_hd__buf_2
X_18801_ _19251_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11136_ _18221_/Q _11059_/X _11140_/S vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16993_ _14243_/A input75/X _16997_/S vssd1 vssd1 vccd1 vccd1 _16994_/A sky130_fd_sc_hd__mux2_1
X_16542__254 _16542__254/A vssd1 vssd1 vccd1 vccd1 _19000_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18732_ _18732_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _11067_/A vssd1 vssd1 vccd1 vccd1 _18251_/D sky130_fd_sc_hd__clkbuf_1
X_15944_ _15939_/Y _15940_/X _15942_/Y _15943_/X vssd1 vssd1 vccd1 vccd1 _15945_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _18756_/Q _09947_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18663_ _14157_/A _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _17618_/CLK _17614_/D vssd1 vssd1 vccd1 vccd1 _17614_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18594_ _18594_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _17545_/CLK _17545_/D vssd1 vssd1 vccd1 vccd1 _17545_/Q sky130_fd_sc_hd__dfxtp_1
X_11969_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12034_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13708_ _17879_/Q _13709_/B _13707_/Y _13376_/X vssd1 vssd1 vccd1 vccd1 _17879_/D
+ sky130_fd_sc_hd__a211o_1
X_14405__579 _14405__579/A vssd1 vssd1 vccd1 vccd1 _18214_/CLK sky130_fd_sc_hd__inv_2
X_17476_ _17476_/A vssd1 vssd1 vccd1 vccd1 _19339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14688_ _14686_/X _14687_/X _14688_/S vssd1 vssd1 vccd1 vccd1 _14688_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _19215_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_1
X_13639_ _13710_/A _13639_/B vssd1 vssd1 vccd1 vccd1 _13640_/A sky130_fd_sc_hd__or2_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16427_ _16471_/A vssd1 vssd1 vccd1 vccd1 _16427_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19146_ _19146_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15309_ _19215_/Q _19103_/Q _18286_/Q _19095_/Q _15308_/X _09631_/X vssd1 vssd1 vccd1
+ vccd1 _15309_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14297__492 _14297__492/A vssd1 vssd1 vccd1 vccd1 _18127_/CLK sky130_fd_sc_hd__inv_2
XFILLER_195_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19077_ _19077_/CLK _19077_/D vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfxtp_1
X_16289_ _16287_/X _16288_/X _16289_/S vssd1 vssd1 vccd1 vccd1 _16289_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18028_ _18029_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09801_/A vssd1 vssd1 vccd1 vccd1 _18831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09732_ _10704_/A vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _09663_/A vssd1 vssd1 vccd1 vccd1 _18911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09594_ _09594_/A vssd1 vssd1 vccd1 vccd1 _18937_/D sky130_fd_sc_hd__clkbuf_1
X_16671__305 _16674__308/A vssd1 vssd1 vccd1 vccd1 _19079_/CLK sky130_fd_sc_hd__inv_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_180 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_191 _09262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19287_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09028_ _08991_/X _19211_/Q _09044_/S vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15677__977 _15677__977/A vssd1 vssd1 vccd1 vccd1 _18694_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13990_ _13740_/A _13989_/X _13978_/X vssd1 vssd1 vccd1 vccd1 _13990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_213_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12941_ _12941_/A _12941_/B _12941_/C _12941_/D vssd1 vssd1 vccd1 vccd1 _12942_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12830_/X _12872_/B vssd1 vssd1 vccd1 vccd1 _12873_/A sky130_fd_sc_hd__and2b_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14696_/A _14611_/B vssd1 vssd1 vccd1 vccd1 _14611_/Y sky130_fd_sc_hd__nor2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14879__796 _14881__798/A vssd1 vssd1 vccd1 vccd1 _18441_/CLK sky130_fd_sc_hd__inv_2
X_11823_ _17928_/Q _11815_/X _11816_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _11823_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15595_/B _15595_/C _15590_/Y vssd1 vssd1 vccd1 vccd1 _15591_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17761_/Q _19282_/Q _17333_/S vssd1 vssd1 vccd1 vccd1 _17331_/B sky130_fd_sc_hd__mux2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14619_/A vssd1 vssd1 vccd1 vccd1 _14543_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _17862_/Q _19291_/Q _17772_/Q vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__mux2_4
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17261_/A vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__clkbuf_1
X_10705_ _18406_/Q _10704_/X _10705_/S vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__mux2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11685_ _19030_/Q _16601_/B vssd1 vssd1 vccd1 vccd1 _16602_/B sky130_fd_sc_hd__and2_1
XFILLER_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16212_ _16208_/X _16211_/X _16271_/S vssd1 vssd1 vccd1 vccd1 _16213_/B sky130_fd_sc_hd__mux2_1
X_19000_ _19000_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_1
X_13424_ input63/X _13431_/B vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__nand2_2
X_17192_ _17194_/B _17195_/A _17191_/X vssd1 vssd1 vccd1 vccd1 _17192_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10636_ _18437_/Q _10135_/A _10636_/S vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16143_ _16194_/A vssd1 vssd1 vccd1 vccd1 _16143_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13355_ _13357_/A vssd1 vssd1 vccd1 vccd1 _13355_/X sky130_fd_sc_hd__clkbuf_2
X_10567_ _10567_/A vssd1 vssd1 vccd1 vccd1 _18499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16728__342 _16728__342/A vssd1 vssd1 vccd1 vccd1 _19121_/CLK sky130_fd_sc_hd__inv_2
X_12306_ _12306_/A _12306_/B _12306_/C _12306_/D vssd1 vssd1 vccd1 vccd1 _12316_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_170_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16074_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16074_/X sky130_fd_sc_hd__buf_1
X_13286_ _13285_/X _13282_/X _13275_/X vssd1 vssd1 vccd1 vccd1 _13286_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ _10120_/X _18529_/Q _10502_/S vssd1 vssd1 vccd1 vccd1 _10499_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15025_ _18464_/Q _15031_/C vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__xor2_1
XFILLER_108_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03402_ clkbuf_0__03402_/X vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12168_ _12166_/X _12168_/B vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__07170_ clkbuf_0__07170_/X vssd1 vssd1 vccd1 vccd1 _11879__362/A sky130_fd_sc_hd__clkbuf_16
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _11119_/A vssd1 vssd1 vccd1 vccd1 _18229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12099_ _12097_/X _12098_/X _12099_/S vssd1 vssd1 vccd1 vccd1 _12195_/A sky130_fd_sc_hd__mux2_1
X_16976_ _16974_/X _16975_/X _16976_/S vssd1 vssd1 vccd1 vccd1 _16976_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ _18715_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_1
X_14823__751 _14824__752/A vssd1 vssd1 vccd1 vccd1 _18394_/CLK sky130_fd_sc_hd__inv_2
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _15927_/A _15927_/B _18861_/Q vssd1 vssd1 vccd1 vccd1 _15927_/X sky130_fd_sc_hd__or3b_1
Xinput6 flash_sck vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18646_ _18657_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03195_ clkbuf_0__03195_/X vssd1 vssd1 vccd1 vccd1 _14514__666/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14809_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14809_/X sky130_fd_sc_hd__buf_1
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18577_ _18577_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17528_ _17878_/CLK _17528_/D vssd1 vssd1 vccd1 vccd1 _17528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17459_ _17742_/Q _19334_/Q _17468_/S vssd1 vssd1 vccd1 vccd1 _17460_/B sky130_fd_sc_hd__mux2_1
XFILLER_220_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16334__230 _16338__234/A vssd1 vssd1 vccd1 vccd1 _18946_/CLK sky130_fd_sc_hd__inv_2
XFILLER_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19129_ _19136_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
X_14453__617 _14455__619/A vssd1 vssd1 vccd1 vccd1 _18252_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09715_ _09715_/A vssd1 vssd1 vccd1 vccd1 _18891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14347__533 _14347__533/A vssd1 vssd1 vccd1 vccd1 _18168_/CLK sky130_fd_sc_hd__inv_2
X_15195__881 _15195__881/A vssd1 vssd1 vccd1 vccd1 _18560_/CLK sky130_fd_sc_hd__inv_2
XFILLER_216_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09646_ _08889_/B _09645_/X _09616_/X vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__o21ai_1
XFILLER_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12232__377 _12234__379/A vssd1 vssd1 vccd1 vccd1 _17541_/CLK sky130_fd_sc_hd__inv_2
XFILLER_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09577_ _09577_/A vssd1 vssd1 vccd1 vccd1 _18944_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16636__277 _16638__279/A vssd1 vssd1 vccd1 vccd1 _19051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03422_ clkbuf_0__03422_/X vssd1 vssd1 vccd1 vccd1 _14882__799/A sky130_fd_sc_hd__clkbuf_16
XFILLER_243_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11470_ _11470_/A vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10421_ _18556_/Q _16097_/A _10420_/X vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13140_ _13777_/A vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__buf_6
X_10352_ _18593_/Q _10351_/X _10352_/S vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14766__705 _14768__707/A vssd1 vssd1 vccd1 vccd1 _18348_/CLK sky130_fd_sc_hd__inv_2
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ _13066_/X _13071_/B vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__and2b_1
X_10283_ _10283_/A vssd1 vssd1 vccd1 vccd1 _18621_/D sky130_fd_sc_hd__clkbuf_1
X_12022_ _12022_/A vssd1 vssd1 vccd1 vccd1 _12099_/S sky130_fd_sc_hd__buf_2
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16830_ _16927_/A _16830_/B vssd1 vssd1 vccd1 vccd1 _16830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13973_ _13973_/A vssd1 vssd1 vccd1 vccd1 _13973_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16761_ _16783_/A _16761_/B vssd1 vssd1 vccd1 vccd1 _16761_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17084__67 _17086__69/A vssd1 vssd1 vccd1 vccd1 _19216_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18500_ _18500_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12924_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_234_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18431_ _18431_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12855_ _17642_/Q _12924_/A _12853_/Y _12854_/X vssd1 vssd1 vccd1 vccd1 _12859_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_185_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15643_ _15808_/C _15643_/B vssd1 vssd1 vccd1 vccd1 _16860_/A sky130_fd_sc_hd__and2_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _17769_/Q input11/X _11831_/C vssd1 vssd1 vccd1 vccd1 _11806_/X sky130_fd_sc_hd__and3b_1
X_15574_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15597_/B sky130_fd_sc_hd__clkbuf_2
X_18362_ _18362_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ _12761_/X _12786_/B vssd1 vssd1 vccd1 vccd1 _12787_/A sky130_fd_sc_hd__and2b_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _17766_/Q _19277_/Q _17381_/B vssd1 vssd1 vccd1 vccd1 _17314_/B sky130_fd_sc_hd__mux2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _17826_/Q vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__inv_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18293_ _18293_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17244_ _17250_/C _17246_/C _17191_/X vssd1 vssd1 vccd1 vccd1 _17244_/Y sky130_fd_sc_hd__o21ai_1
X_14456_ _14456_/A vssd1 vssd1 vccd1 vccd1 _14456_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__03982_ _15754_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03982_/X sky130_fd_sc_hd__clkbuf_16
X_11668_ _11668_/A vssd1 vssd1 vccd1 vccd1 _17509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPeripherals_163 vssd1 vssd1 vccd1 vccd1 Peripherals_163/HI io_oeb[1] sky130_fd_sc_hd__conb_1
X_13407_ _14079_/A vssd1 vssd1 vccd1 vccd1 _13407_/X sky130_fd_sc_hd__clkbuf_4
XPeripherals_174 vssd1 vssd1 vccd1 vccd1 Peripherals_174/HI io_oeb[37] sky130_fd_sc_hd__conb_1
X_17175_ _19235_/Q _17169_/X _17164_/X vssd1 vssd1 vccd1 vccd1 _17176_/B sky130_fd_sc_hd__o21ai_1
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10619_ _10619_/A vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__clkbuf_1
XPeripherals_185 vssd1 vssd1 vccd1 vccd1 Peripherals_185/HI wb_data_o[24] sky130_fd_sc_hd__conb_1
X_14387_ _14449_/A vssd1 vssd1 vccd1 vccd1 _14387_/X sky130_fd_sc_hd__buf_1
XPeripherals_196 vssd1 vssd1 vccd1 vccd1 io_oeb[3] Peripherals_196/LO sky130_fd_sc_hd__conb_1
X_11599_ _17573_/Q _10713_/A _11599_/S vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14517__669 _14517__669/A vssd1 vssd1 vccd1 vccd1 _18304_/CLK sky130_fd_sc_hd__inv_2
X_16126_ _18775_/Q _18633_/Q _18783_/Q _18617_/Q _16117_/A _16138_/A vssd1 vssd1 vccd1
+ vccd1 _16126_/X sky130_fd_sc_hd__mux4_1
X_13338_ _13240_/X _13330_/X _13337_/X vssd1 vssd1 vccd1 vccd1 _13338_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _16057_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _18883_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _13268_/X _13259_/X _13260_/X vssd1 vssd1 vccd1 vccd1 _13269_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15008_ _15034_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _15009_/A sky130_fd_sc_hd__and2_1
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15099__819 _15099__819/A vssd1 vssd1 vccd1 vccd1 _18495_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03416_ _14846_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03416_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_238_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16959_ _18062_/Q _18054_/Q _18046_/Q _18038_/Q _16870_/X _16871_/X vssd1 vssd1 vccd1
+ vccd1 _16959_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09500_ _09500_/A vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09431_ _09431_/A vssd1 vssd1 vccd1 vccd1 _19051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18629_ _18629_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03178_ clkbuf_0__03178_/X vssd1 vssd1 vccd1 vccd1 _14427__596/A sky130_fd_sc_hd__clkbuf_16
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _09362_/A vssd1 vssd1 vccd1 vccd1 _19082_/D sky130_fd_sc_hd__clkbuf_1
X_16555__264 _16555__264/A vssd1 vssd1 vccd1 vccd1 _19010_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09293_ _19115_/Q _08958_/X _09293_/S vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput140 _17720_/Q vssd1 vssd1 vccd1 vccd1 probe_blink[0] sky130_fd_sc_hd__buf_2
Xoutput151 _11863_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[17] sky130_fd_sc_hd__buf_2
X_17299__75 _17302__78/A vssd1 vssd1 vccd1 vccd1 _19271_/CLK sky130_fd_sc_hd__inv_2
Xoutput162 _18065_/Q vssd1 vssd1 vccd1 vccd1 wb_stall_o sky130_fd_sc_hd__buf_2
XFILLER_88_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03971_ clkbuf_0__03971_/X vssd1 vssd1 vccd1 vccd1 _15698__994/A sky130_fd_sc_hd__clkbuf_16
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _10970_/A vssd1 vssd1 vccd1 vccd1 _18290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09629_ _09626_/A _09626_/B _09616_/X vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__o21ai_1
XFILLER_216_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12640_ _12640_/A _12640_/B vssd1 vssd1 vccd1 vccd1 _17600_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12571_ _12469_/S _12566_/X _12568_/Y _12570_/Y vssd1 vssd1 vccd1 vccd1 _12774_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03405_ clkbuf_0__03405_/X vssd1 vssd1 vccd1 vccd1 _14793__727/A sky130_fd_sc_hd__clkbuf_16
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11522_/A vssd1 vssd1 vccd1 vccd1 _18035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15290_ _18571_/Q _15207_/X _15270_/X _15289_/X vssd1 vssd1 vccd1 vccd1 _18571_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14241_ _14239_/X _14240_/X _18472_/Q vssd1 vssd1 vccd1 vccd1 _14241_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15879__174 _15879__174/A vssd1 vssd1 vccd1 vccd1 _18849_/CLK sky130_fd_sc_hd__inv_2
X_16684__315 _16685__316/A vssd1 vssd1 vccd1 vccd1 _19089_/CLK sky130_fd_sc_hd__inv_2
X_11453_ _11453_/A vssd1 vssd1 vccd1 vccd1 _18092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _10404_/A _18556_/Q _16097_/A vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__and3_1
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _14256_/A vssd1 vssd1 vccd1 vccd1 _14172_/X sky130_fd_sc_hd__buf_1
XFILLER_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11384_ _11457_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11400_/S sky130_fd_sc_hd__or2_2
XFILLER_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13123_ _13710_/A vssd1 vssd1 vccd1 vccd1 _16715_/B sky130_fd_sc_hd__buf_6
Xclkbuf_1_0__f__03198_ clkbuf_0__03198_/X vssd1 vssd1 vccd1 vccd1 _14535__684/A sky130_fd_sc_hd__clkbuf_16
XFILLER_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10335_ _10335_/A vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__clkbuf_1
X_18980_ _19014_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13054_ _13049_/X _13054_/B vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__and2b_1
XFILLER_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17931_ _19136_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10266_ _18628_/Q _10189_/X _10266_/S vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12005_ _11950_/X _11954_/X _12005_/S vssd1 vssd1 vccd1 vccd1 _12005_/X sky130_fd_sc_hd__mux2_1
X_17862_ _18031_/CLK _17862_/D vssd1 vssd1 vccd1 vccd1 _17862_/Q sky130_fd_sc_hd__dfxtp_1
X_10197_ _10197_/A vssd1 vssd1 vccd1 vccd1 _18688_/D sky130_fd_sc_hd__clkbuf_1
X_15436__930 _15440__934/A vssd1 vssd1 vccd1 vccd1 _18617_/CLK sky130_fd_sc_hd__inv_2
XFILLER_227_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16813_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16813_/X sky130_fd_sc_hd__buf_4
X_17793_ _19136_/CLK _17793_/D vssd1 vssd1 vccd1 vccd1 _17793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17057__45 _17058__46/A vssd1 vssd1 vccd1 vccd1 _19194_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _19111_/Q _17788_/Q vssd1 vssd1 vccd1 vccd1 _16744_/X sky130_fd_sc_hd__or2b_1
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13956_ _17963_/Q _13962_/B vssd1 vssd1 vccd1 vccd1 _13956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12907_ _12907_/A vssd1 vssd1 vccd1 vccd1 _17665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13887_ _17938_/Q _13878_/X _13886_/Y vssd1 vssd1 vccd1 vccd1 _17938_/D sky130_fd_sc_hd__o21a_1
XFILLER_235_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18414_ _18414_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
X_12838_ _12838_/A vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__buf_2
X_15626_ _15626_/A _15626_/B vssd1 vssd1 vccd1 vccd1 _15626_/X sky130_fd_sc_hd__or2_1
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ input24/X vssd1 vssd1 vccd1 vccd1 _19394_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18345_ _18345_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12769_ _12769_/A vssd1 vssd1 vccd1 vccd1 _12769_/Y sky130_fd_sc_hd__inv_2
X_15557_ _18646_/Q _15557_/B _15557_/C vssd1 vssd1 vccd1 vccd1 _15561_/B sky130_fd_sc_hd__and3_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15488_ _18653_/Q _15489_/B _15488_/C vssd1 vssd1 vccd1 vccd1 _15528_/B sky130_fd_sc_hd__and3_1
X_18276_ _18276_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput20 io_in[2] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_12
X_17227_ _17225_/B _17225_/C _17225_/D _19250_/Q vssd1 vssd1 vccd1 vccd1 _17228_/C
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_0__03965_ _15662_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03965_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_174_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 vga_vsync vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_8
Xinput42 wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_4
X_17158_ _17159_/A _17158_/B _17162_/D vssd1 vssd1 vccd1 vccd1 _17158_/X sky130_fd_sc_hd__and3_1
XFILLER_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput75 wb_sel_i[0] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_4
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03796_ clkbuf_0__03796_/X vssd1 vssd1 vccd1 vccd1 _15400__901/A sky130_fd_sc_hd__clkbuf_16
X_16109_ _18593_/Q _18609_/Q _18735_/Q _18516_/Q _16106_/X _16108_/X vssd1 vssd1 vccd1
+ vccd1 _16110_/B sky130_fd_sc_hd__mux4_1
X_17089_ _13361_/X _17101_/A _12182_/A vssd1 vssd1 vccd1 vccd1 _17089_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09980_ _18773_/Q _09943_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08931_ _08931_/A vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08862_ _09148_/B _09148_/C _09476_/A vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__or3b_4
XFILLER_112_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08793_ _19345_/Q _08792_/X _08796_/S vssd1 vssd1 vccd1 vccd1 _08794_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__07167_ _11873_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__07167_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09414_ _09826_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09430_/S sky130_fd_sc_hd__or2_2
XFILLER_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09345_ _09345_/A vssd1 vssd1 vccd1 vccd1 _19089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15760__1044 _15760__1044/A vssd1 vssd1 vccd1 vccd1 _18761_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09276_ _09276_/A vssd1 vssd1 vccd1 vccd1 _19122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10120_ _10120_/A vssd1 vssd1 vccd1 vccd1 _10120_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_164_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10051_ _10073_/S vssd1 vssd1 vccd1 vccd1 _10064_/S sky130_fd_sc_hd__buf_2
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _13268_/X _13802_/X _13805_/X vssd1 vssd1 vccd1 vccd1 _13810_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _14802_/A vssd1 vssd1 vccd1 vccd1 _14790_/X sky130_fd_sc_hd__buf_1
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13741_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10953_ _08868_/X _18297_/Q _10959_/S vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13672_ _13237_/X _13666_/X _13661_/X vssd1 vssd1 vccd1 vccd1 _13672_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16460_ _18974_/Q _16468_/B vssd1 vssd1 vccd1 vccd1 _16460_/Y sky130_fd_sc_hd__nand2_1
X_10884_ _10884_/A vssd1 vssd1 vccd1 vccd1 _18332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _12622_/B _12622_/C _12622_/A vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16391_ _18976_/Q _16391_/B vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__xnor2_1
XFILLER_223_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18130_ _18130_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_1
X_15342_ _15298_/X _15339_/X _15341_/X _15305_/X vssd1 vssd1 vccd1 vccd1 _15342_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12554_ _17630_/Q vssd1 vssd1 vccd1 vccd1 _12746_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_185_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04368_ clkbuf_0__04368_/X vssd1 vssd1 vccd1 vccd1 _16313__213/A sky130_fd_sc_hd__clkbuf_16
X_11505_ _18042_/Q _11338_/A _11509_/S vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169__875 _15173__879/A vssd1 vssd1 vccd1 vccd1 _18551_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18061_ _18061_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
X_15273_ _15273_/A vssd1 vssd1 vccd1 vccd1 _15273_/X sky130_fd_sc_hd__clkbuf_4
X_12485_ _12440_/X _12426_/X _12556_/A vssd1 vssd1 vccd1 vccd1 _12485_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14224_ _14224_/A vssd1 vssd1 vccd1 vccd1 _18082_/D sky130_fd_sc_hd__clkbuf_1
X_17012_ _17043_/A vssd1 vssd1 vccd1 vccd1 _17012_/X sky130_fd_sc_hd__buf_1
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _18099_/Q _11282_/X _11436_/S vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16649__287 _16649__287/A vssd1 vssd1 vccd1 vccd1 _19061_/CLK sky130_fd_sc_hd__inv_2
XFILLER_138_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11367_ _11321_/X _18130_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _11368_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _09685_/X _18605_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__mux2_1
X_14086_ _12555_/X _14077_/S _14085_/Y vssd1 vssd1 vccd1 vccd1 _18012_/D sky130_fd_sc_hd__o21a_1
XFILLER_180_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18963_ _18963_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11298_ _11298_/A vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__clkbuf_1
X_17413__103 _17414__104/A vssd1 vssd1 vccd1 vccd1 _19316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13037_ _13032_/X _13037_/B vssd1 vssd1 vccd1 vccd1 _13038_/A sky130_fd_sc_hd__and2b_1
X_17914_ _19128_/CLK _17914_/D vssd1 vssd1 vccd1 vccd1 _17914_/Q sky130_fd_sc_hd__dfxtp_2
X_10249_ _10249_/A vssd1 vssd1 vccd1 vccd1 _18636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18894_ _18894_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17845_ _18921_/CLK _17845_/D vssd1 vssd1 vccd1 vccd1 _17845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17776_ _17776_/CLK _17776_/D vssd1 vssd1 vccd1 vccd1 _17776_/Q sky130_fd_sc_hd__dfxtp_1
X_14779__715 _14783__719/A vssd1 vssd1 vccd1 vccd1 _18358_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14988_ _18457_/Q _14978_/X _14987_/Y _15057_/A vssd1 vssd1 vccd1 vccd1 _14989_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__04164_ _16074_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04164_/X sky130_fd_sc_hd__clkbuf_16
X_13939_ _17957_/Q _13941_/B vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16658_ _16658_/A vssd1 vssd1 vccd1 vccd1 _16658_/X sky130_fd_sc_hd__buf_1
XFILLER_90_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15609_ _18656_/Q _15610_/B vssd1 vssd1 vccd1 vccd1 _15615_/C sky130_fd_sc_hd__and2_1
X_15113__830 _15114__831/A vssd1 vssd1 vccd1 vccd1 _18506_/CLK sky130_fd_sc_hd__inv_2
X_15860__159 _15860__159/A vssd1 vssd1 vccd1 vccd1 _18834_/CLK sky130_fd_sc_hd__inv_2
X_16589_ _16602_/A _16593_/C vssd1 vssd1 vccd1 vccd1 _16589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09130_ _18666_/Q vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__clkbuf_4
X_18328_ _18996_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09061_ _10851_/A _10869_/A vssd1 vssd1 vccd1 vccd1 _09077_/S sky130_fd_sc_hd__nor2_2
XFILLER_148_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18259_ _18259_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09963_ _10132_/A vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_65_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17963_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08914_ _08910_/X _19299_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 _08915_/A sky130_fd_sc_hd__mux2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09894_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09895_/B sky130_fd_sc_hd__or2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _09446_/A hold12/A vssd1 vssd1 vccd1 vccd1 _09441_/B sky130_fd_sc_hd__nor2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778__1059 _15778__1059/A vssd1 vssd1 vccd1 vccd1 _18776_/CLK sky130_fd_sc_hd__inv_2
XFILLER_217_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__08199_ _13109_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__08199_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_73_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08776_ _16294_/B _09647_/A vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__nand2_4
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14164__443 _14165__444/A vssd1 vssd1 vccd1 vccd1 _18051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09328_ _19096_/Q _08955_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _09281_/S vssd1 vssd1 vccd1 vccd1 _09272_/S sky130_fd_sc_hd__buf_2
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ _17556_/Q _18021_/Q _12270_/S vssd1 vssd1 vccd1 vccd1 _12271_/B sky130_fd_sc_hd__mux2_1
XFILLER_154_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11221_ _11221_/A vssd1 vssd1 vccd1 vccd1 _18187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11152_ _11152_/A vssd1 vssd1 vccd1 vccd1 _18216_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16722__337 _16724__339/A vssd1 vssd1 vccd1 vccd1 _19116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ _10103_/A vssd1 vssd1 vccd1 vccd1 _18723_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11083_ _09051_/X _18244_/Q _11085_/S vssd1 vssd1 vccd1 vccd1 _11084_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15960_ _15986_/A _16035_/B _15967_/C vssd1 vssd1 vccd1 vccd1 _15961_/B sky130_fd_sc_hd__mux2_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ _14922_/B _17847_/Q _14936_/A _17846_/Q vssd1 vssd1 vccd1 vccd1 _14913_/C
+ sky130_fd_sc_hd__o31ai_1
X_10034_ _18749_/Q _09943_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__mux2_1
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17630_ _18012_/CLK _17630_/D vssd1 vssd1 vccd1 vccd1 _17630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ _18027_/CLK _17561_/D vssd1 vssd1 vccd1 vccd1 _17561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11985_ _17159_/A _19232_/Q _17169_/B _17173_/B _11961_/X _11957_/S vssd1 vssd1 vccd1
+ vccd1 _12091_/B sky130_fd_sc_hd__mux4_2
XFILLER_216_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19300_ _19300_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03799_ clkbuf_0__03799_/X vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__clkbuf_16
X_16512_ _16506_/A _16298_/Y _16514_/C _16511_/X _16507_/X vssd1 vssd1 vccd1 vccd1
+ _16512_/X sky130_fd_sc_hd__a41o_1
X_13724_ _13724_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13724_/Y sky130_fd_sc_hd__nor2_1
X_10936_ _10936_/A vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17492_ _19336_/Q _17492_/B vssd1 vssd1 vccd1 vccd1 _17493_/D sky130_fd_sc_hd__xnor2_1
XFILLER_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19231_ _19251_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16443_ _16439_/X _16441_/Y _16480_/A vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__a21oi_1
X_13655_ _17861_/Q _13649_/X _13654_/Y vssd1 vssd1 vccd1 vccd1 _17861_/D sky130_fd_sc_hd__o21a_1
X_10867_ _18339_/Q _10812_/X _10867_/S vssd1 vssd1 vccd1 vccd1 _10868_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A vssd1 vssd1 vccd1 vccd1 _17591_/D sky130_fd_sc_hd__clkbuf_1
X_19162_ _19162_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _17841_/Q _16522_/A _13589_/S vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__mux2_1
X_16374_ _17794_/Q _16422_/B vssd1 vssd1 vccd1 vccd1 _16376_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _18368_/Q _10797_/X _10804_/S vssd1 vssd1 vccd1 vccd1 _10799_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18113_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_1
X_12537_ _12360_/X _12369_/X _12473_/X _12535_/X _12569_/S _12502_/A vssd1 vssd1 vccd1
+ vccd1 _12537_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04851_ _17075_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04851_/X sky130_fd_sc_hd__clkbuf_16
X_15325_ _15298_/X _15322_/X _15324_/X _15305_/X vssd1 vssd1 vccd1 vccd1 _15325_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19093_ _19093_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03802_ _15429_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03802_/X sky130_fd_sc_hd__clkbuf_16
X_18044_ _18044_/CLK _18044_/D vssd1 vssd1 vccd1 vccd1 _18044_/Q sky130_fd_sc_hd__dfxtp_1
X_12468_ _12515_/A vssd1 vssd1 vccd1 vccd1 _12469_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_145_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15256_ _18932_/Q vssd1 vssd1 vccd1 vccd1 _15281_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11419_ _11419_/A vssd1 vssd1 vccd1 vccd1 _18107_/D sky130_fd_sc_hd__clkbuf_1
X_14207_ _18075_/Q input33/X _14207_/S vssd1 vssd1 vccd1 vccd1 _14208_/A sky130_fd_sc_hd__mux2_1
X_15187_ _19143_/Q _19144_/Q _18658_/Q vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__mux2_1
X_12399_ _17596_/Q vssd1 vssd1 vccd1 vccd1 _12622_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_235_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14069_ _14069_/A _14069_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__or3b_2
X_18946_ _18946_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03595_ _15131_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03595_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18877_ _18889_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17828_ _18482_/CLK _17828_/D vssd1 vssd1 vccd1 vccd1 _17828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17759_ _19327_/CLK _17759_/D vssd1 vssd1 vccd1 vccd1 _17759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341__528 _14342__529/A vssd1 vssd1 vccd1 vccd1 _18163_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09113_ _19189_/Q _09112_/X _09117_/S vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ _09043_/X _19207_/Q _09044_/S vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09946_ _18478_/Q vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__buf_4
XFILLER_131_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04840_ clkbuf_0__04840_/X vssd1 vssd1 vccd1 vccd1 _17024__19/A sky130_fd_sc_hd__clkbuf_16
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09877_ _09869_/B _09877_/B _09895_/C vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__and3b_1
XINSDIODE2_11 _10180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_22 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_33 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_44 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _19316_/Q _08804_/X _08828_/S vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_55 _13493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_66 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__07490_ clkbuf_0__07490_/X vssd1 vssd1 vccd1 vccd1 _12226__372/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_77 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_88 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08759_ hold1/X vssd1 vssd1 vccd1 vccd1 _10219_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_99 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _17866_/Q _17652_/Q _18003_/Q vssd1 vssd1 vccd1 vccd1 _11771_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10721_ _10721_/A vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ _13434_/X _13437_/X _13439_/Y _13213_/X vssd1 vssd1 vccd1 vccd1 _17794_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10652_ _09277_/X _18430_/Q _10654_/S vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13750_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_210_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10583_ _10583_/A _10583_/B _09894_/A vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__or3b_4
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ _15041_/A vssd1 vssd1 vccd1 vccd1 _18466_/D sky130_fd_sc_hd__clkbuf_1
X_12253_ _12245_/X _12253_/B vssd1 vssd1 vccd1 vccd1 _12254_/A sky130_fd_sc_hd__and2b_1
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ hold18/X _11204_/B vssd1 vssd1 vccd1 vccd1 _11220_/S sky130_fd_sc_hd__nor2_2
X_12184_ _12184_/A vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__buf_2
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18800_ _18993_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _11135_/A vssd1 vssd1 vccd1 vccd1 _18222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16992_ _19144_/Q _16797_/A _16991_/X _16915_/X vssd1 vssd1 vccd1 vccd1 _19144_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18731_ _18731_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11066_ _18251_/Q _11065_/X _11066_/S vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__mux2_1
X_15943_ _18871_/Q _15943_/B _15943_/C vssd1 vssd1 vccd1 vccd1 _15943_/X sky130_fd_sc_hd__and3_1
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _10017_/A vssd1 vssd1 vccd1 vccd1 _18757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18662_ _14157_/A _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15874_ _15880_/A vssd1 vssd1 vccd1 vccd1 _15874_/X sky130_fd_sc_hd__buf_1
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _17618_/CLK _17613_/D vssd1 vssd1 vccd1 vccd1 _17613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _18593_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _17544_/CLK _17544_/D vssd1 vssd1 vccd1 vccd1 _17544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11968_ _17778_/Q vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_205_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13707_ _13707_/A _13709_/B vssd1 vssd1 vccd1 vccd1 _13707_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17475_ _16736_/A _17475_/B vssd1 vssd1 vccd1 vccd1 _17476_/A sky130_fd_sc_hd__and2b_1
X_10919_ _18312_/Q _10895_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10920_/A sky130_fd_sc_hd__mux2_1
X_11899_ _11975_/S vssd1 vssd1 vccd1 vccd1 _11956_/S sky130_fd_sc_hd__buf_2
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14687_ _18408_/Q _18400_/Q _19313_/Q _17717_/Q _14594_/X _14595_/X vssd1 vssd1 vccd1
+ vccd1 _14687_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19214_ _19214_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _16426_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _16471_/A sky130_fd_sc_hd__or2_1
X_13638_ _17858_/Q _16522_/A _13642_/S vssd1 vssd1 vccd1 vccd1 _13639_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19145_ _19146_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13569_ _13636_/A vssd1 vssd1 vccd1 vccd1 _13569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15308_ _15308_/A vssd1 vssd1 vccd1 vccd1 _15308_/X sky130_fd_sc_hd__buf_2
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ _19076_/CLK _19076_/D vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16288_ _18782_/Q _18640_/Q _18790_/Q _18624_/Q _16195_/A _16182_/X vssd1 vssd1 vccd1
+ vccd1 _16288_/X sky130_fd_sc_hd__mux4_1
X_15777__1058 _15778__1059/A vssd1 vssd1 vccd1 vccd1 _18775_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18027_ _18027_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15239_ _15244_/A _15223_/X _15267_/A _15238_/X vssd1 vssd1 vccd1 vccd1 _15239_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09800_ _18831_/Q _09758_/X _09800_/S vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09731_ _09731_/A vssd1 vssd1 vccd1 vccd1 _18857_/D sky130_fd_sc_hd__clkbuf_1
X_18929_ _18929_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09662_ _18911_/Q _09265_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09593_ _18937_/Q _09498_/X _09597_/S vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__05079_ clkbuf_0__05079_/X vssd1 vssd1 vccd1 vccd1 _17402__94/A sky130_fd_sc_hd__clkbuf_16
XFILLER_242_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_170 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_181 _11753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_192 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17611_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09027_ _09056_/S vssd1 vssd1 vccd1 vccd1 _09044_/S sky130_fd_sc_hd__buf_2
XFILLER_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126__840 _15128__842/A vssd1 vssd1 vccd1 vccd1 _18516_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15873__169 _15873__169/A vssd1 vssd1 vccd1 vccd1 _18844_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14510__664 _14510__664/A vssd1 vssd1 vccd1 vccd1 _18299_/CLK sky130_fd_sc_hd__inv_2
X_09929_ _09929_/A vssd1 vssd1 vccd1 vccd1 _18785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12940_ _17667_/Q _13092_/B vssd1 vssd1 vccd1 vccd1 _12941_/D sky130_fd_sc_hd__xor2_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12871_ _17981_/Q _17655_/Q _12944_/B vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__mux2_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15430__925 _15434__929/A vssd1 vssd1 vccd1 vccd1 _18612_/CLK sky130_fd_sc_hd__inv_2
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _19076_/Q _18340_/Q _17574_/Q _18792_/Q _14579_/X _14580_/X vssd1 vssd1 vccd1
+ vccd1 _14611_/B sky130_fd_sc_hd__mux4_2
XFILLER_57_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ _17909_/Q _11812_/X _11821_/Y input16/X _11796_/X vssd1 vssd1 vccd1 vccd1
+ _11822_/X sky130_fd_sc_hd__a221o_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15595_/B _15595_/C _15551_/A vssd1 vssd1 vccd1 vccd1 _15590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11753_ _11753_/A vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _16559_/C _16426_/A vssd1 vssd1 vccd1 vccd1 _14619_/A sky130_fd_sc_hd__and2_2
XFILLER_242_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10704_ _10704_/A vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17264_/B _17265_/B _17260_/C vssd1 vssd1 vccd1 vccd1 _17261_/A sky130_fd_sc_hd__and3b_1
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _19029_/Q _19028_/Q _16596_/B vssd1 vssd1 vccd1 vccd1 _16601_/B sky130_fd_sc_hd__and3_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _16209_/X _16210_/X _16286_/S vssd1 vssd1 vccd1 vccd1 _16211_/X sky130_fd_sc_hd__mux2_1
X_13423_ _13761_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13432_/S sky130_fd_sc_hd__nor2_1
X_10635_ _10635_/A vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__clkbuf_1
X_17191_ _17191_/A vssd1 vssd1 vccd1 vccd1 _17191_/X sky130_fd_sc_hd__buf_2
XFILLER_174_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ _14069_/A _13354_/B _14069_/B vssd1 vssd1 vccd1 vccd1 _13357_/A sky130_fd_sc_hd__or3_4
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16142_ _16223_/A _16142_/B vssd1 vssd1 vccd1 vccd1 _16142_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10566_ _10112_/X _18499_/Q _10574_/S vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _17561_/Q _17489_/B vssd1 vssd1 vccd1 vccd1 _12306_/D sky130_fd_sc_hd__xnor2_1
XFILLER_182_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13285_ _13441_/A vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__buf_4
XFILLER_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10497_ _10497_/A vssd1 vssd1 vccd1 vccd1 _18530_/D sky130_fd_sc_hd__clkbuf_1
X_15024_ _15024_/A vssd1 vssd1 vccd1 vccd1 _18463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03401_ clkbuf_0__03401_/X vssd1 vssd1 vccd1 vccd1 _14776__714/A sky130_fd_sc_hd__clkbuf_16
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12167_ _17527_/Q _17724_/Q _12170_/S vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ _18229_/Q _11059_/X _11122_/S vssd1 vssd1 vccd1 vccd1 _11119_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12098_ _11918_/X _11927_/X _12098_/S vssd1 vssd1 vccd1 vccd1 _12098_/X sky130_fd_sc_hd__mux2_1
X_16975_ _18154_/Q _18146_/Q _18138_/Q _18282_/Q _16809_/X _16810_/X vssd1 vssd1 vccd1
+ vccd1 _16975_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14411__584 _14411__584/A vssd1 vssd1 vccd1 vccd1 _18219_/CLK sky130_fd_sc_hd__inv_2
X_18714_ _18714_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15926_ _15927_/A _15927_/B vssd1 vssd1 vccd1 vccd1 _15926_/Y sky130_fd_sc_hd__nand2_1
X_11049_ _11049_/A vssd1 vssd1 vccd1 vccd1 _18257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 io_in[10] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_232_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18645_ _18657_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03194_ clkbuf_0__03194_/X vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14808_ _14808_/A vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__buf_1
XFILLER_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18576_ _18922_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17527_ _17878_/CLK _17527_/D vssd1 vssd1 vccd1 vccd1 _17527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14739_ _14561_/X _14732_/Y _14734_/Y _14736_/Y _14738_/Y vssd1 vssd1 vccd1 vccd1
+ _14739_/X sky130_fd_sc_hd__o32a_1
XFILLER_178_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ _17458_/A vssd1 vssd1 vccd1 vccd1 _19333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16409_ _18969_/Q _17807_/Q vssd1 vssd1 vccd1 vccd1 _16410_/S sky130_fd_sc_hd__xnor2_1
XFILLER_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19128_ _19128_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19059_ _19059_/CLK _19059_/D vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04579_ clkbuf_0__04579_/X vssd1 vssd1 vccd1 vccd1 _16685__316/A sky130_fd_sc_hd__clkbuf_16
XFILLER_102_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _09694_/X _18891_/Q _09716_/S vssd1 vssd1 vccd1 vccd1 _09715_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__and2_1
XFILLER_228_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _18944_/Q _09501_/X _09578_/S vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__mux2_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_196_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03421_ clkbuf_0__03421_/X vssd1 vssd1 vccd1 vccd1 _14873__791/A sky130_fd_sc_hd__clkbuf_16
XFILLER_51_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15683__982 _15685__984/A vssd1 vssd1 vccd1 vccd1 _18699_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10420_ _10420_/A vssd1 vssd1 vccd1 vccd1 _10420_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ _18473_/Q vssd1 vssd1 vccd1 vccd1 _10351_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13070_ _17938_/Q _17700_/Q _13070_/S vssd1 vssd1 vccd1 vccd1 _13071_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10282_ _18621_/Q _10186_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _11945_/X _12016_/X _12020_/X vssd1 vssd1 vccd1 vccd1 _12201_/A sky130_fd_sc_hd__o21ai_1
XFILLER_2_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15204__889 _15204__889/A vssd1 vssd1 vccd1 vccd1 _18568_/CLK sky130_fd_sc_hd__inv_2
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ _19131_/Q _19129_/Q _16767_/S vssd1 vssd1 vccd1 vccd1 _16761_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13972_ _17969_/Q _13967_/X _13971_/Y vssd1 vssd1 vccd1 vccd1 _17969_/D sky130_fd_sc_hd__o21a_1
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15711_/X sky130_fd_sc_hd__buf_1
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _17665_/Q _12846_/B _12835_/X _17664_/Q vssd1 vssd1 vccd1 vccd1 _12931_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16691_ _16687_/X _16689_/X _16795_/A vssd1 vssd1 vccd1 vccd1 _19091_/D sky130_fd_sc_hd__o21ba_1
XFILLER_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15776__1057 _15776__1057/A vssd1 vssd1 vccd1 vccd1 _18774_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18430_ _18430_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
X_15642_ _15642_/A _15642_/B vssd1 vssd1 vccd1 vccd1 _15642_/X sky130_fd_sc_hd__and2_1
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _17643_/Q _12921_/A _12838_/A _17651_/Q vssd1 vssd1 vccd1 vccd1 _12854_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11805_ _11837_/A _13278_/B vssd1 vssd1 vccd1 vccd1 _11831_/C sky130_fd_sc_hd__nor2_1
X_18361_ _18361_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15579_/A _15573_/B _15585_/C vssd1 vssd1 vccd1 vccd1 _15573_/X sky130_fd_sc_hd__or3_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _17638_/Q _17997_/Q _12862_/B vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__mux2_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03619_ clkbuf_0__03619_/X vssd1 vssd1 vccd1 vccd1 _15195__881/A sky130_fd_sc_hd__clkbuf_16
XFILLER_214_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17312_/A vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14524_/A vssd1 vssd1 vccd1 vccd1 _14524_/X sky130_fd_sc_hd__buf_1
X_11736_ _11736_/A vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _18292_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ _19254_/Q vssd1 vssd1 vccd1 vccd1 _17250_/C sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03981_ _15748_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03981_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _17509_/Q _09691_/A _11671_/S vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPeripherals_164 vssd1 vssd1 vccd1 vccd1 Peripherals_164/HI io_oeb[6] sky130_fd_sc_hd__conb_1
X_13406_ _16767_/S _13405_/B _13405_/Y _13376_/X vssd1 vssd1 vccd1 vccd1 _17786_/D
+ sky130_fd_sc_hd__a211o_1
X_17174_ _17186_/C vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10618_ _10135_/X _18445_/Q _10618_/S vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__mux2_1
XPeripherals_175 vssd1 vssd1 vccd1 vccd1 Peripherals_175/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ _11598_/A vssd1 vssd1 vccd1 vccd1 _17574_/D sky130_fd_sc_hd__clkbuf_1
X_14386_ _14386_/A vssd1 vssd1 vccd1 vccd1 _14386_/X sky130_fd_sc_hd__buf_1
XPeripherals_186 vssd1 vssd1 vccd1 vccd1 Peripherals_186/HI wb_data_o[25] sky130_fd_sc_hd__conb_1
XPeripherals_197 vssd1 vssd1 vccd1 vccd1 io_oeb[4] Peripherals_197/LO sky130_fd_sc_hd__conb_1
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ _16123_/X _16124_/X _16276_/A vssd1 vssd1 vccd1 vccd1 _16125_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13337_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13337_/X sky130_fd_sc_hd__clkbuf_4
X_10549_ _10549_/A vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16056_ _16056_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _18882_/D sky130_fd_sc_hd__nor2_1
X_13268_ _14083_/A vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__buf_4
XFILLER_108_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15007_ _15005_/A _14991_/X _15006_/Y _14993_/X vssd1 vssd1 vccd1 vccd1 _15008_/B
+ sky130_fd_sc_hd__a22o_1
X_12219_ _13951_/A vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _16057_/A _13180_/B _13198_/Y _13187_/X vssd1 vssd1 vccd1 vccd1 _17733_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_243_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03415_ _14840_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03415_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16958_ _19210_/Q _19162_/Q _18273_/Q _18265_/Q _16828_/A _16868_/X vssd1 vssd1 vccd1
+ vccd1 _16958_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15909_ _18868_/Q _15937_/B _15909_/C vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__and3_1
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16889_ _16818_/X _16888_/X _16860_/X vssd1 vssd1 vccd1 vccd1 _16889_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09430_ _08941_/X _19051_/Q _09430_/S vssd1 vssd1 vccd1 vccd1 _09431_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18628_ _18628_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03177_ clkbuf_0__03177_/X vssd1 vssd1 vccd1 vccd1 _14424__594/A sky130_fd_sc_hd__clkbuf_16
XFILLER_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _19082_/Q _09080_/X _09369_/S vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18559_ _18559_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _09292_/A vssd1 vssd1 vccd1 vccd1 _19116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput130 _19395_/X vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__buf_2
XFILLER_217_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput141 _17721_/Q vssd1 vssd1 vccd1 vccd1 probe_blink[1] sky130_fd_sc_hd__buf_2
Xoutput152 _11866_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_161_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03970_ clkbuf_0__03970_/X vssd1 vssd1 vccd1 vccd1 _15705_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16642__282 _16643__283/A vssd1 vssd1 vccd1 vccd1 _19056_/CLK sky130_fd_sc_hd__inv_2
XFILLER_247_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09628_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _18932_/D sky130_fd_sc_hd__nor2_1
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09559_ _09559_/A vssd1 vssd1 vccd1 vccd1 _18952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ _12408_/X _12569_/X _12580_/A vssd1 vssd1 vccd1 vccd1 _12570_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14772__710 _14773__711/A vssd1 vssd1 vccd1 vccd1 _18353_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03404_ clkbuf_0__03404_/X vssd1 vssd1 vccd1 vccd1 _14789__724/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f__07172_ clkbuf_0__07172_/X vssd1 vssd1 vccd1 vccd1 _11886__367/A sky130_fd_sc_hd__clkbuf_16
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11521_ _18035_/Q _11335_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ _18918_/Q _18919_/Q _18920_/Q _18921_/Q _18470_/Q _18471_/Q vssd1 vssd1 vccd1
+ vccd1 _14240_/X sky130_fd_sc_hd__mux4_1
X_11452_ _18092_/Q _11279_/X _11454_/S vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10403_ _10403_/A _10403_/B _10403_/C _10403_/D vssd1 vssd1 vccd1 vccd1 _16097_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ _11383_/A _11383_/B _09025_/A vssd1 vssd1 vccd1 vccd1 _11438_/B sky130_fd_sc_hd__or3b_4
XFILLER_178_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03197_ clkbuf_0__03197_/X vssd1 vssd1 vccd1 vccd1 _14529__679/A sky130_fd_sc_hd__clkbuf_16
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13122_ _17454_/A vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__clkbuf_4
X_10334_ _18599_/Q _10333_/X _10343_/S vssd1 vssd1 vccd1 vccd1 _10335_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13053_ _17943_/Q _17695_/Q _13053_/S vssd1 vssd1 vccd1 vccd1 _13054_/B sky130_fd_sc_hd__mux2_1
X_17930_ _19136_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10265_ _10265_/A vssd1 vssd1 vccd1 vccd1 _18629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12004_ _11976_/X _11949_/X _12008_/S vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17861_ _18031_/CLK _17861_/D vssd1 vssd1 vccd1 vccd1 _17861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10196_ _18688_/Q _10195_/X _10199_/S vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _18808_/Q vssd1 vssd1 vccd1 vccd1 _16828_/A sky130_fd_sc_hd__clkbuf_4
X_17792_ _19135_/CLK _17792_/D vssd1 vssd1 vccd1 vccd1 _17792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16743_ _19135_/Q _16741_/S _16742_/X vssd1 vssd1 vccd1 vccd1 _16743_/X sky130_fd_sc_hd__a21o_1
X_13955_ _13184_/X _13946_/X _13954_/Y _13951_/X vssd1 vssd1 vccd1 vccd1 _17962_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _12894_/X _12906_/B vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__and2b_1
XFILLER_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13886_ _13777_/X _13885_/X _13880_/X vssd1 vssd1 vccd1 vccd1 _13886_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18413_ _18413_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15625_ _15626_/A _15626_/B vssd1 vssd1 vccd1 vccd1 _15630_/B sky130_fd_sc_hd__nand2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19393_ input27/X vssd1 vssd1 vccd1 vccd1 _19393_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_234_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12837_ _17636_/Q _12850_/A _12932_/A _17639_/Q vssd1 vssd1 vccd1 vccd1 _12843_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14523__674 _14523__674/A vssd1 vssd1 vccd1 vccd1 _18309_/CLK sky130_fd_sc_hd__inv_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18344_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
X_15556_ _18646_/Q _15562_/C vssd1 vssd1 vccd1 vccd1 _15558_/B sky130_fd_sc_hd__nor2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12767_/X _12446_/X _12768_/S vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__mux2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11719_ _11719_/A vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__clkbuf_1
X_18275_ _18275_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_15487_ _15489_/B _15488_/C _18653_/Q vssd1 vssd1 vccd1 vccd1 _15528_/A sky130_fd_sc_hd__a21oi_1
X_12699_ _12707_/B _12707_/C _12695_/X vssd1 vssd1 vccd1 vccd1 _12700_/B sky130_fd_sc_hd__o21ai_1
XFILLER_238_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _17237_/D vssd1 vssd1 vccd1 vccd1 _17233_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 io_in[20] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
XFILLER_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03964_ _15661_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03964_/X sky130_fd_sc_hd__clkbuf_16
Xinput21 io_in[3] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_6
XFILLER_163_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput32 wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput54 wb_cyc_i vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_4
X_17157_ _17157_/A vssd1 vssd1 vccd1 vccd1 _19230_/D sky130_fd_sc_hd__clkbuf_1
Xinput65 wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_6
Xinput76 wb_sel_i[1] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__03795_ clkbuf_0__03795_/X vssd1 vssd1 vccd1 vccd1 _15397__899/A sky130_fd_sc_hd__clkbuf_16
XFILLER_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16108_ _16138_/A vssd1 vssd1 vccd1 vccd1 _16108_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08930_ _08929_/X _19295_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 _08931_/A sky130_fd_sc_hd__mux2_1
X_16039_ _18879_/Q _18878_/Q _18877_/Q vssd1 vssd1 vccd1 vccd1 _16049_/C sky130_fd_sc_hd__and3_1
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08861_ hold20/X vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_229_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08792_ _18884_/Q vssd1 vssd1 vccd1 vccd1 _08792_/X sky130_fd_sc_hd__buf_2
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04378_ _16359_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04378_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_77_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _09413_/A vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09344_ _19089_/Q _09262_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _09345_/A sky130_fd_sc_hd__mux2_1
X_14424__594 _14424__594/A vssd1 vssd1 vccd1 vccd1 _18229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_240_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14836__762 _14838__764/A vssd1 vssd1 vccd1 vccd1 _18405_/CLK sky130_fd_sc_hd__inv_2
XFILLER_244_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ _19122_/Q _09274_/X _09281_/S vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15775__1056 _15776__1057/A vssd1 vssd1 vccd1 vccd1 _18773_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _10094_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10073_/S sky130_fd_sc_hd__nor2_2
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466__628 _14467__629/A vssd1 vssd1 vccd1 vccd1 _18263_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13740_ _13740_/A _13743_/B vssd1 vssd1 vccd1 vccd1 _13740_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952_ _10952_/A vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13671_ _17866_/Q _13659_/X _13670_/Y vssd1 vssd1 vccd1 vccd1 _17866_/D sky130_fd_sc_hd__o21a_1
X_10883_ _18332_/Q _10809_/X _10885_/S vssd1 vssd1 vccd1 vccd1 _10884_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _15410_/A vssd1 vssd1 vccd1 vccd1 _15410_/X sky130_fd_sc_hd__buf_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _12622_/A _12622_/B _12622_/C vssd1 vssd1 vccd1 vccd1 _12626_/B sky130_fd_sc_hd__and3_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _17800_/Q _16393_/B vssd1 vssd1 vccd1 vccd1 _16391_/B sky130_fd_sc_hd__xor2_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ _15341_/A _15303_/X vssd1 vssd1 vccd1 vccd1 _15341_/X sky130_fd_sc_hd__or2b_1
X_12553_ _17627_/Q vssd1 vssd1 vccd1 vccd1 _12737_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16354__245 _16355__246/A vssd1 vssd1 vccd1 vccd1 _18961_/CLK sky130_fd_sc_hd__inv_2
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04367_ clkbuf_0__04367_/X vssd1 vssd1 vccd1 vccd1 _16333_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18060_ _18060_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
X_11504_ _11504_/A vssd1 vssd1 vccd1 vccd1 _18043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ _18999_/Q _18961_/Q _18953_/Q _17542_/Q _15209_/X _15218_/X vssd1 vssd1 vccd1
+ vccd1 _15272_/X sky130_fd_sc_hd__mux4_1
X_12484_ _18005_/Q _12351_/X _12762_/A vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__a21o_1
XFILLER_185_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ _18082_/Q input40/X _14229_/S vssd1 vssd1 vccd1 vccd1 _14224_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11435_ _11435_/A vssd1 vssd1 vccd1 vccd1 _18100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11366_ _11381_/S vssd1 vssd1 vccd1 vccd1 _11375_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15696__992 _15696__992/A vssd1 vssd1 vccd1 vccd1 _18709_/CLK sky130_fd_sc_hd__inv_2
X_10317_ _10317_/A vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__clkbuf_1
X_14291__488 _14292__489/A vssd1 vssd1 vccd1 vccd1 _18123_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14085_ _13812_/X _14077_/S _14060_/X vssd1 vssd1 vccd1 vccd1 _14085_/Y sky130_fd_sc_hd__a21oi_1
X_18962_ _18962_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_1
X_11297_ _18157_/Q _11276_/X _11301_/S vssd1 vssd1 vccd1 vccd1 _11298_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13036_ _17948_/Q _17690_/Q _13099_/B vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__mux2_1
X_17913_ _19128_/CLK _17913_/D vssd1 vssd1 vccd1 vccd1 _17913_/Q sky130_fd_sc_hd__dfxtp_1
X_10248_ _18636_/Q _10189_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _10249_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18893_ _18893_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17844_ _19136_/CLK _17844_/D vssd1 vssd1 vccd1 vccd1 _17844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10179_ _10179_/A vssd1 vssd1 vccd1 vccd1 _18694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17775_ _17779_/CLK _17775_/D vssd1 vssd1 vccd1 vccd1 _17775_/Q sky130_fd_sc_hd__dfxtp_1
X_14987_ _14987_/A _14998_/C vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_219_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04163_ _16068_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04163_/X sky130_fd_sc_hd__clkbuf_16
X_13938_ _13150_/X _13925_/X _13936_/Y _13937_/X vssd1 vssd1 vccd1 vccd1 _17956_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12332__394 _12332__394/A vssd1 vssd1 vccd1 vccd1 _17575_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13869_ _17934_/Q _13863_/B _13867_/X _13868_/X vssd1 vssd1 vccd1 vccd1 _17934_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15608_ _15606_/X _15607_/Y _15581_/A vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__a21oi_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16588_ _16588_/A vssd1 vssd1 vccd1 vccd1 _16593_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18327_ _19013_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15612_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _09358_/B _10770_/C _10770_/A vssd1 vssd1 vccd1 vccd1 _10869_/A sky130_fd_sc_hd__nand3b_4
X_18258_ _18258_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _19245_/Q _17209_/B vssd1 vssd1 vccd1 vccd1 _17216_/D sky130_fd_sc_hd__and2_1
XFILLER_190_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18189_ _18189_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16708__330 _16710__332/A vssd1 vssd1 vccd1 vccd1 _19105_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09962_ _18474_/Q vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__buf_2
XFILLER_44_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08913_ _08942_/S vssd1 vssd1 vccd1 vccd1 _08930_/S sky130_fd_sc_hd__clkbuf_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09893_/A vssd1 vssd1 vccd1 vccd1 _18803_/D sky130_fd_sc_hd__clkbuf_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08844_/A vssd1 vssd1 vccd1 vccd1 _08844_/Y sky130_fd_sc_hd__inv_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__08198_ _13103_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__08198_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08775_ _08889_/B _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__and3_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _09327_/A vssd1 vssd1 vccd1 vccd1 _19097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09258_ _10638_/A _10094_/A vssd1 vssd1 vccd1 vccd1 _09281_/S sky130_fd_sc_hd__nor2_2
XFILLER_193_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09189_ _09189_/A vssd1 vssd1 vccd1 vccd1 _19163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14884__800 _14886__802/A vssd1 vssd1 vccd1 vccd1 _18445_/CLK sky130_fd_sc_hd__inv_2
X_11220_ _18187_/Q _11065_/X _11220_/S vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11151_ _11150_/X _18216_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _11152_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ _18723_/Q _10060_/X _10104_/S vssd1 vssd1 vccd1 vccd1 _10103_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _11082_/A vssd1 vssd1 vccd1 vccd1 _18245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14910_ _18466_/Q _14910_/B vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__xnor2_1
X_10033_ _10033_/A vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _15890_/A vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__buf_1
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ _18021_/CLK _17560_/D vssd1 vssd1 vccd1 vccd1 _17560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11984_ _19234_/Q vssd1 vssd1 vccd1 vccd1 _17173_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_217_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03798_ clkbuf_0__03798_/X vssd1 vssd1 vccd1 vccd1 _15415__914/A sky130_fd_sc_hd__clkbuf_16
X_16511_ _16511_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16511_/X sky130_fd_sc_hd__or2_1
X_13723_ _17884_/Q _13715_/X _13722_/Y _13710_/X vssd1 vssd1 vccd1 vccd1 _17884_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17491_ _19334_/Q _17491_/B vssd1 vssd1 vccd1 vccd1 _17493_/C sky130_fd_sc_hd__xnor2_1
XFILLER_17_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10935_ _18305_/Q _10892_/X _10941_/S vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19230_ _19251_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _16469_/A vssd1 vssd1 vccd1 vccd1 _16480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13654_ _13709_/A _13649_/X _13532_/X vssd1 vssd1 vccd1 vccd1 _13654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16655__292 _16655__292/A vssd1 vssd1 vccd1 vccd1 _19066_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10866_ _10866_/A vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _12610_/C _12605_/B _12709_/B vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__and3b_1
XFILLER_176_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ _19161_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _17796_/Q _17795_/Q _16383_/A vssd1 vssd1 vccd1 vccd1 _16422_/B sky130_fd_sc_hd__or3_1
X_13585_ _13265_/X _13574_/B _13584_/Y _13569_/X vssd1 vssd1 vccd1 vccd1 _17840_/D
+ sky130_fd_sc_hd__a211oi_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10797_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__buf_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18112_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__04850_ _17074_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04850_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15324_ _15324_/A _15303_/X vssd1 vssd1 vccd1 vccd1 _15324_/X sky130_fd_sc_hd__or2b_1
X_12536_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12569_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_223_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19092_ _19092_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03801_ _15423_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03801_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_185_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18043_ _18043_/CLK _18043_/D vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
X_15255_ _19213_/Q _19101_/Q _18284_/Q _19093_/Q _15291_/A _09613_/A vssd1 vssd1 vccd1
+ vccd1 _15255_/X sky130_fd_sc_hd__mux4_1
X_12467_ _12463_/X _12464_/X _12465_/X _12466_/X _12567_/S _12408_/A vssd1 vssd1 vccd1
+ vccd1 _12467_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ _14206_/A vssd1 vssd1 vccd1 vccd1 _18074_/D sky130_fd_sc_hd__clkbuf_1
X_11418_ _11344_/X _18107_/Q _11418_/S vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15186_ _19141_/Q _19142_/Q _15626_/B vssd1 vssd1 vccd1 vccd1 _15186_/X sky130_fd_sc_hd__mux2_1
X_12398_ _17592_/Q _12610_/A _12394_/X _12622_/B _12396_/X _12397_/X vssd1 vssd1 vccd1
+ vccd1 _12398_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14785__720 _14786__721/A vssd1 vssd1 vccd1 vccd1 _18363_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14137_ _13147_/B _13441_/X _14136_/Y _11697_/X vssd1 vssd1 vccd1 vccd1 _18031_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11349_ _18138_/Q _11259_/X _11357_/S vssd1 vssd1 vccd1 vccd1 _11350_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14068_ input72/X _16518_/B _14055_/X _14067_/X _15083_/B vssd1 vssd1 vccd1 vccd1
+ _18005_/D sky130_fd_sc_hd__a311o_1
X_18945_ _18945_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03594_ _15125_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03594_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_239_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13019_ _13019_/A _13019_/B _13019_/C _13019_/D vssd1 vssd1 vccd1 vccd1 _13020_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_140_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18876_ _18876_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17827_ _19136_/CLK _17827_/D vssd1 vssd1 vccd1 vccd1 _17827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17758_ _19290_/CLK _17758_/D vssd1 vssd1 vccd1 vccd1 _17758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15774__1055 _15776__1057/A vssd1 vssd1 vccd1 vccd1 _18772_/CLK sky130_fd_sc_hd__inv_2
X_17689_ _17945_/CLK _17689_/D vssd1 vssd1 vccd1 vccd1 _17689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09112_ _10710_/A vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__buf_2
XFILLER_202_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09043_ _11335_/A vssd1 vssd1 vccd1 vccd1 _09043_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ _09945_/A vssd1 vssd1 vccd1 vccd1 _18781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15456__945 _15457__946/A vssd1 vssd1 vccd1 vccd1 _18632_/CLK sky130_fd_sc_hd__inv_2
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _18799_/Q _15808_/C _09875_/X vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_12 _10189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_34 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08827_/A vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_45 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_56 _13434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_67 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_78 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_89 _19389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ _18933_/Q vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__inv_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17024__19 _17024__19/A vssd1 vssd1 vccd1 vccd1 _19168_/CLK sky130_fd_sc_hd__inv_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10720_ _18401_/Q _10695_/X _10726_/S vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__mux2_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10651_ _10651_/A vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13370_ _12034_/A _13355_/X _13369_/Y _13359_/X vssd1 vssd1 vccd1 vccd1 _17778_/D
+ sky130_fd_sc_hd__a211o_1
X_10582_ _11222_/A _11456_/B _10987_/B vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__or3_4
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _16216_/A _15040_/B vssd1 vssd1 vccd1 vccd1 _15041_/A sky130_fd_sc_hd__and2_1
X_12252_ _17551_/Q _18026_/Q _12318_/B vssd1 vssd1 vccd1 vccd1 _12253_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _11203_/A vssd1 vssd1 vccd1 vccd1 _18195_/D sky130_fd_sc_hd__clkbuf_1
X_12183_ _17515_/Q _12180_/X _12182_/X _17518_/Q vssd1 vssd1 vccd1 vccd1 _12192_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_14849__772 _14850__773/A vssd1 vssd1 vccd1 vccd1 _18417_/CLK sky130_fd_sc_hd__inv_2
X_11134_ _18222_/Q _11056_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _11135_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16991_ _16892_/X _16980_/X _16990_/Y vssd1 vssd1 vccd1 vccd1 _16991_/X sky130_fd_sc_hd__a21o_1
XFILLER_150_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18730_ _18730_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
X_11065_ _18661_/Q vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__buf_2
X_15942_ _15943_/B _15943_/C _18871_/Q vssd1 vssd1 vccd1 vccd1 _15942_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ _18757_/Q _09943_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__mux2_1
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _14157_/A _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17612_ _17618_/CLK _17612_/D vssd1 vssd1 vccd1 vccd1 _17612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_7_1_wb_clk_i clkbuf_opt_7_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_7_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_221_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18592_ _18592_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _17543_/CLK _17543_/D vssd1 vssd1 vccd1 vccd1 _17543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11967_ _11962_/X _11966_/X _12091_/A vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__mux2_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13706_ _13712_/B vssd1 vssd1 vccd1 vccd1 _13709_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17474_ _17737_/Q _19339_/Q _17474_/S vssd1 vssd1 vccd1 vccd1 _17475_/B sky130_fd_sc_hd__mux2_1
X_10918_ _10918_/A vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__clkbuf_1
X_14686_ _19177_/Q _19169_/Q _19201_/Q _18336_/Q _14591_/X _14592_/X vssd1 vssd1 vccd1
+ vccd1 _14686_/X sky130_fd_sc_hd__mux4_2
X_11898_ _11892_/X _11895_/X _12032_/S vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19213_ _19213_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
X_16425_ _16428_/C vssd1 vssd1 vccd1 vccd1 _16534_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13637_ _13265_/X _13626_/B _13635_/Y _13636_/X vssd1 vssd1 vccd1 vccd1 _17857_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10849_ _18347_/Q _10812_/X _10849_/S vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19144_ _19144_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13568_ _17835_/Q _13568_/B vssd1 vssd1 vccd1 vccd1 _13568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15307_ _15307_/A vssd1 vssd1 vccd1 vccd1 _15307_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12519_ _12394_/X _17595_/Q _17596_/Q _17597_/Q _12426_/S _12359_/A vssd1 vssd1 vccd1
+ vccd1 _12519_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19075_ _19075_/CLK _19075_/D vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16287_ _18632_/Q _18507_/Q _18913_/Q _18515_/Q _16182_/A _16117_/A vssd1 vssd1 vccd1
+ vccd1 _16287_/X sky130_fd_sc_hd__mux4_2
X_13499_ _13499_/A vssd1 vssd1 vccd1 vccd1 _13499_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18026_ _18029_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15238_ _15229_/X _15237_/X _09615_/A vssd1 vssd1 vccd1 vccd1 _15238_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09730_ _18857_/Q _09729_/X _09733_/S vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18928_ _18928_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_228_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ _09661_/A vssd1 vssd1 vccd1 vccd1 _18912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18859_ _18859_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ _09592_/A vssd1 vssd1 vccd1 vccd1 _18938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__05078_ clkbuf_0__05078_/X vssd1 vssd1 vccd1 vccd1 _17395__88/A sky130_fd_sc_hd__clkbuf_16
XFILLER_78_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_160 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_171 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_182 _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_193 _10120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09026_ _11223_/A _11024_/A vssd1 vssd1 vccd1 vccd1 _09056_/S sky130_fd_sc_hd__or2_2
XFILLER_152_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09928_ _18785_/Q _09274_/X _09932_/S vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09859_ _09859_/A _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__and3_1
XFILLER_86_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _12870_/A vssd1 vssd1 vccd1 vccd1 _17654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _17843_/Q _11821_/B vssd1 vssd1 vccd1 vccd1 _11821_/Y sky130_fd_sc_hd__nor2_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _18996_/Q _18995_/Q vssd1 vssd1 vccd1 vccd1 _16426_/A sky130_fd_sc_hd__nor2_1
XFILLER_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11752_ _17772_/Q _17881_/Q vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__and2b_2
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10703_ _10703_/A vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11683_ _19027_/Q _19026_/Q _19025_/Q _16588_/A vssd1 vssd1 vccd1 vccd1 _16596_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _18778_/Q _18636_/Q _18786_/Q _18620_/Q _16158_/X _16182_/X vssd1 vssd1 vccd1
+ vccd1 _16210_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13422_ _13541_/C _13541_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__or3b_2
X_17190_ _17190_/A vssd1 vssd1 vccd1 vccd1 _19239_/D sky130_fd_sc_hd__clkbuf_1
X_10634_ _18438_/Q _10132_/A _10636_/S vssd1 vssd1 vccd1 vccd1 _10635_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16141_ _18438_/Q _18688_/Q _18696_/Q _18704_/Q _16112_/X _10405_/A vssd1 vssd1 vccd1
+ vccd1 _16142_/B sky130_fd_sc_hd__mux4_1
X_13353_ _13541_/C vssd1 vssd1 vccd1 vccd1 _14069_/B sky130_fd_sc_hd__buf_2
X_10565_ _10580_/S vssd1 vssd1 vccd1 vccd1 _10574_/S sky130_fd_sc_hd__buf_2
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _17560_/Q _17492_/B vssd1 vssd1 vccd1 vccd1 _12306_/C sky130_fd_sc_hd__xnor2_1
XFILLER_154_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14177__454 _14177__454/A vssd1 vssd1 vccd1 vccd1 _18062_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13284_ _17753_/Q _13280_/X _13283_/Y vssd1 vssd1 vccd1 vccd1 _17753_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10496_ _10117_/X _18530_/Q _10502_/S vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15023_ _15034_/A _15023_/B vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__and2_1
X_12235_ _12320_/A vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__buf_1
XFILLER_216_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03400_ clkbuf_0__03400_/X vssd1 vssd1 vccd1 vccd1 _14768__707/A sky130_fd_sc_hd__clkbuf_16
X_12166_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11117_/A vssd1 vssd1 vccd1 vccd1 _18230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12097_ _11898_/X _11903_/X _12012_/X _12096_/X _12037_/S _12029_/A vssd1 vssd1 vccd1
+ vccd1 _12097_/X sky130_fd_sc_hd__mux4_1
X_16974_ _18122_/Q _18114_/Q _18106_/Q _18098_/Q _16893_/X _16894_/X vssd1 vssd1 vccd1
+ vccd1 _16974_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18713_ _18713_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ _18862_/Q _17824_/Q vssd1 vssd1 vccd1 vccd1 _15927_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11048_ _18257_/Q _11047_/X _11057_/S vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 io_in[11] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18644_ _18657_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03193_ clkbuf_0__03193_/X vssd1 vssd1 vccd1 vccd1 _14510__664/A sky130_fd_sc_hd__clkbuf_16
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735__348 _16735__348/A vssd1 vssd1 vccd1 vccd1 _19127_/CLK sky130_fd_sc_hd__inv_2
X_15787_ _15799_/A vssd1 vssd1 vccd1 vccd1 _15787_/X sky130_fd_sc_hd__buf_1
X_18575_ _18922_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_1
X_12999_ _17952_/Q _17685_/Q _12999_/S vssd1 vssd1 vccd1 vccd1 _13000_/B sky130_fd_sc_hd__mux2_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17526_ _17526_/CLK _17526_/D vssd1 vssd1 vccd1 vccd1 _17526_/Q sky130_fd_sc_hd__dfxtp_1
X_14738_ _14640_/X _14737_/X _14604_/A vssd1 vssd1 vccd1 vccd1 _14738_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17457_ _17454_/X _17457_/B vssd1 vssd1 vccd1 vccd1 _17458_/A sky130_fd_sc_hd__and2b_1
X_14669_ _14667_/X _14668_/X _14688_/S vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16408_ _16402_/B _16405_/Y _18970_/Q vssd1 vssd1 vccd1 vccd1 _16411_/C sky130_fd_sc_hd__a21oi_1
XFILLER_242_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17401__93 _17402__94/A vssd1 vssd1 vccd1 vccd1 _19306_/CLK sky130_fd_sc_hd__inv_2
XFILLER_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16339_ _16339_/A vssd1 vssd1 vccd1 vccd1 _16339_/X sky130_fd_sc_hd__buf_1
X_19127_ _19127_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14830__757 _14832__759/A vssd1 vssd1 vccd1 vccd1 _18400_/CLK sky130_fd_sc_hd__inv_2
X_19058_ _19058_/CLK _19058_/D vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18009_ _18010_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04578_ clkbuf_0__04578_/X vssd1 vssd1 vccd1 vccd1 _16680__312/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09713_ _09713_/A vssd1 vssd1 vccd1 vccd1 _18892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09644_ _09644_/A vssd1 vssd1 vccd1 vccd1 _18927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09575_ _09575_/A vssd1 vssd1 vccd1 vccd1 _18945_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03420_ clkbuf_0__03420_/X vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_224_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10350_ _10350_/A vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__clkbuf_1
X_14354__539 _14354__539/A vssd1 vssd1 vccd1 vccd1 _18174_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _09880_/B _09856_/B _09005_/Y _09006_/X _09008_/X vssd1 vssd1 vccd1 vccd1
+ _09009_/X sky130_fd_sc_hd__a2111o_1
X_10281_ _10281_/A vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12020_ _12020_/A _12020_/B vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__or2_1
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17069__55 _17071__57/A vssd1 vssd1 vccd1 vccd1 _19204_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13971_ _13719_/A _13968_/X _13920_/X vssd1 vssd1 vccd1 vccd1 _13971_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15393__895 _15395__897/A vssd1 vssd1 vccd1 vccd1 _18582_/CLK sky130_fd_sc_hd__inv_2
X_12922_ _17661_/Q _12920_/X _12921_/X _17660_/Q vssd1 vssd1 vccd1 vccd1 _12931_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16690_ _16690_/A vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _16061_/A _15641_/B vssd1 vssd1 vccd1 vccd1 _18668_/D sky130_fd_sc_hd__nor2_1
X_12853_ _17644_/Q _12920_/A vssd1 vssd1 vccd1 vccd1 _12853_/Y sky130_fd_sc_hd__nor2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _17934_/Q _11785_/X _11800_/X _11803_/X vssd1 vssd1 vccd1 vccd1 _11804_/X
+ sky130_fd_sc_hd__o211a_4
X_18360_ _18360_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15572_ _18649_/Q _15572_/B _15572_/C vssd1 vssd1 vccd1 vccd1 _15585_/C sky130_fd_sc_hd__and3_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A vssd1 vssd1 vccd1 vccd1 _17637_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17311_ _17304_/X _17311_/B vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__and2b_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _17914_/Q _17564_/Q _17769_/Q vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__mux2_4
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _18291_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A vssd1 vssd1 vccd1 vccd1 _19253_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03980_ _15742_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03980_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ _11666_/A vssd1 vssd1 vccd1 vccd1 _17510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13405_ _13746_/A _13405_/B vssd1 vssd1 vccd1 vccd1 _13405_/Y sky130_fd_sc_hd__nor2_1
X_17173_ _19235_/Q _17173_/B _19233_/Q _17173_/D vssd1 vssd1 vccd1 vccd1 _17186_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_127_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10617_ _10617_/A vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__clkbuf_1
XPeripherals_165 vssd1 vssd1 vccd1 vccd1 Peripherals_165/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_167_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPeripherals_176 vssd1 vssd1 vccd1 vccd1 Peripherals_176/HI io_out[2] sky130_fd_sc_hd__conb_1
X_11597_ _17574_/Q _10710_/A _11599_/S vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__mux2_1
XPeripherals_187 vssd1 vssd1 vccd1 vccd1 Peripherals_187/HI wb_data_o[26] sky130_fd_sc_hd__conb_1
X_16124_ _18711_/Q _18719_/Q _18727_/Q _18492_/Q _16198_/A _16172_/A vssd1 vssd1 vccd1
+ vccd1 _16124_/X sky130_fd_sc_hd__mux4_1
XPeripherals_198 vssd1 vssd1 vccd1 vccd1 io_oeb[5] Peripherals_198/LO sky130_fd_sc_hd__conb_1
X_13336_ _17771_/Q _13329_/X _13335_/Y vssd1 vssd1 vccd1 vccd1 _17771_/D sky130_fd_sc_hd__o21a_1
X_10548_ _18507_/Q _10112_/A _10556_/S vssd1 vssd1 vccd1 vccd1 _10549_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16055_ _16055_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _18881_/D sky130_fd_sc_hd__nor2_1
X_13267_ _17749_/Q _13252_/X _13266_/Y vssd1 vssd1 vccd1 vccd1 _17749_/D sky130_fd_sc_hd__o21a_1
X_14255__459 _14255__459/A vssd1 vssd1 vccd1 vccd1 _18094_/CLK sky130_fd_sc_hd__inv_2
X_10479_ _10479_/A vssd1 vssd1 vccd1 vccd1 _18538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15006_ _15006_/A _15014_/C vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nor2_1
X_12218_ _12218_/A _12218_/B _12218_/C vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__or3_1
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13198_ _17733_/Q _13208_/B vssd1 vssd1 vccd1 vccd1 _13198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12149_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12149_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16702__325 _16704__327/A vssd1 vssd1 vccd1 vccd1 _19100_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__03414_ _14839_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03414_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16957_ _16955_/X _16956_/X _16976_/S vssd1 vssd1 vccd1 vccd1 _16957_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15908_ _17819_/Q _15917_/B _17818_/Q vssd1 vssd1 vccd1 vccd1 _15909_/C sky130_fd_sc_hd__o21ai_1
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16888_ _16819_/X _16878_/Y _16880_/Y _16884_/Y _16887_/Y vssd1 vssd1 vccd1 vccd1
+ _16888_/X sky130_fd_sc_hd__o32a_1
XFILLER_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18627_ _18627_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03176_ clkbuf_0__03176_/X vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _09375_/S vssd1 vssd1 vccd1 vccd1 _09369_/S sky130_fd_sc_hd__clkbuf_2
X_18558_ _18655_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17509_ _17509_/CLK _17509_/D vssd1 vssd1 vccd1 vccd1 _17509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09291_ _19116_/Q _08955_/X _09293_/S vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18489_ _18489_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17386__81 _17386__81/A vssd1 vssd1 vccd1 vccd1 _19294_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18013_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_242_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15800__120 _15801__121/A vssd1 vssd1 vccd1 vccd1 _18792_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput120 _11722_/X vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_2
Xoutput131 _19396_/X vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__buf_2
Xoutput142 _18064_/Q vssd1 vssd1 vccd1 vccd1 wb_ack_o sky130_fd_sc_hd__buf_2
XFILLER_217_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput153 _11804_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[1] sky130_fd_sc_hd__buf_2
XFILLER_161_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09627_ _09625_/X _09630_/A _09616_/X vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__o21ai_1
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ _08937_/X _18952_/Q _09560_/S vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14360__543 _14361__544/A vssd1 vssd1 vccd1 vccd1 _18178_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03403_ clkbuf_0__03403_/X vssd1 vssd1 vccd1 vccd1 _14782__718/A sky130_fd_sc_hd__clkbuf_16
X_09489_ _18885_/Q vssd1 vssd1 vccd1 vccd1 _09489_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_197_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__07171_ clkbuf_0__07171_/X vssd1 vssd1 vccd1 vccd1 _12229_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11520_ _11520_/A vssd1 vssd1 vccd1 vccd1 _18036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _11451_/A vssd1 vssd1 vccd1 vccd1 _18093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ _10402_/A vssd1 vssd1 vccd1 vccd1 _10403_/C sky130_fd_sc_hd__inv_2
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11382_ _11382_/A vssd1 vssd1 vccd1 vccd1 _18123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03196_ clkbuf_0__03196_/X vssd1 vssd1 vccd1 vccd1 _14520__671/A sky130_fd_sc_hd__clkbuf_16
X_13121_ _13892_/A vssd1 vssd1 vccd1 vccd1 _17454_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10333_ _18479_/Q vssd1 vssd1 vccd1 vccd1 _10333_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _13052_/A vssd1 vssd1 vccd1 vccd1 _17694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10264_ _18629_/Q _10186_/X _10266_/S vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12003_ _11994_/X _11996_/X _11997_/X _12001_/X _12087_/S _12029_/A vssd1 vssd1 vccd1
+ vccd1 _12003_/X sky130_fd_sc_hd__mux4_1
X_17860_ _18031_/CLK _17860_/D vssd1 vssd1 vccd1 vccd1 _17860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10195_ _18474_/Q vssd1 vssd1 vccd1 vccd1 _10195_/X sky130_fd_sc_hd__buf_2
XFILLER_132_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16811_ _18056_/Q _18048_/Q _18040_/Q _18032_/Q _16809_/X _16810_/X vssd1 vssd1 vccd1
+ vccd1 _16811_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17791_ _17923_/CLK _17791_/D vssd1 vssd1 vccd1 vccd1 _17791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _17962_/Q _13962_/B vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__nor2_1
X_16742_ _17786_/Q _19130_/Q vssd1 vssd1 vccd1 vccd1 _16742_/X sky130_fd_sc_hd__and2b_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15139__851 _15142__854/A vssd1 vssd1 vccd1 vccd1 _18527_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12905_ _17971_/Q _17665_/Q _12908_/S vssd1 vssd1 vccd1 vccd1 _12906_/B sky130_fd_sc_hd__mux2_1
XFILLER_246_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _13885_/A vssd1 vssd1 vccd1 vccd1 _13885_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18412_ _18465_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
X_12836_ _17637_/Q _12834_/X _12835_/X _17647_/Q vssd1 vssd1 vccd1 vccd1 _12836_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_15624_ _15624_/A _15624_/B vssd1 vssd1 vccd1 vccd1 _18658_/D sky130_fd_sc_hd__nor2_1
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ input26/X vssd1 vssd1 vccd1 vccd1 _19392_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15555_ _15583_/A vssd1 vssd1 vccd1 vccd1 _15579_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18343_ _18343_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _17589_/Q _17590_/Q _17591_/Q _17592_/Q _12443_/X _12556_/A vssd1 vssd1 vccd1
+ vccd1 _12767_/X sky130_fd_sc_hd__mux4_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11718_ _11717_/X _17929_/Q vssd1 vssd1 vccd1 vccd1 _11719_/A sky130_fd_sc_hd__and2b_4
X_18274_ _18274_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_15486_ _17831_/Q _15486_/B vssd1 vssd1 vccd1 vccd1 _15488_/C sky130_fd_sc_hd__nand2_1
XFILLER_148_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12698_ _12707_/B _12707_/C vssd1 vssd1 vccd1 vccd1 _12700_/A sky130_fd_sc_hd__and2_1
X_17225_ _19250_/Q _17225_/B _17225_/C _17225_/D vssd1 vssd1 vccd1 vccd1 _17237_/D
+ sky130_fd_sc_hd__and4_1
Xclkbuf_0__03963_ _15655_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03963_/X sky130_fd_sc_hd__clkbuf_16
X_14437_ _14443_/A vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__buf_1
Xinput11 io_in[21] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
XFILLER_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ _08798_/X _17534_/Q _11653_/S vssd1 vssd1 vccd1 vccd1 _11650_/A sky130_fd_sc_hd__mux2_1
Xinput22 io_in[4] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_6
XFILLER_35_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15443__936 _15444__937/A vssd1 vssd1 vccd1 vccd1 _18623_/CLK sky130_fd_sc_hd__inv_2
XFILLER_174_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput33 wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
X_17156_ _17159_/B _17189_/B _17156_/C vssd1 vssd1 vccd1 vccd1 _17157_/A sky130_fd_sc_hd__and3b_1
Xinput44 wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
XFILLER_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput55 wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_8
X_14368_ _14380_/A vssd1 vssd1 vccd1 vccd1 _14368_/X sky130_fd_sc_hd__buf_1
XFILLER_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput66 wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_6
Xclkbuf_1_1__f__03794_ clkbuf_0__03794_/X vssd1 vssd1 vccd1 vccd1 _15389__892/A sky130_fd_sc_hd__clkbuf_16
XFILLER_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput77 wb_sel_i[2] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _16182_/A vssd1 vssd1 vccd1 vccd1 _16138_/A sky130_fd_sc_hd__buf_2
X_13319_ _17766_/Q _13304_/X _13318_/Y vssd1 vssd1 vccd1 vccd1 _17766_/D sky130_fd_sc_hd__o21a_1
XFILLER_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17087_ _17384_/A vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__buf_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16038_ _18877_/Q vssd1 vssd1 vccd1 vccd1 _16044_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08860_ _08860_/A _16559_/B vssd1 vssd1 vccd1 vccd1 _09148_/C sky130_fd_sc_hd__nand2_1
XFILLER_233_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08791_ _08791_/A vssd1 vssd1 vccd1 vccd1 _19346_/D sky130_fd_sc_hd__clkbuf_1
X_17989_ _19247_/CLK _17989_/D vssd1 vssd1 vccd1 vccd1 _17989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__04377_ _16353_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04377_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09412_ _08941_/X _19059_/Q _09412_/S vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03159_ clkbuf_0__03159_/X vssd1 vssd1 vccd1 vccd1 _14336__524/A sky130_fd_sc_hd__clkbuf_16
XFILLER_164_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09343_ _09343_/A vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09274_ _18475_/Q vssd1 vssd1 vccd1 vccd1 _09274_/X sky130_fd_sc_hd__buf_2
XFILLER_244_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14843__767 _14843__767/A vssd1 vssd1 vccd1 vccd1 _18410_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _08989_/A vssd1 vssd1 vccd1 vccd1 _19212_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _08830_/X _18298_/Q _10959_/S vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13670_ _13669_/X _13666_/X _13661_/X vssd1 vssd1 vccd1 vccd1 _13670_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10882_ _10882_/A vssd1 vssd1 vccd1 vccd1 _18333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15807__126 _15807__126/A vssd1 vssd1 vccd1 vccd1 _18798_/CLK sky130_fd_sc_hd__inv_2
XFILLER_232_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12621_ _12622_/B _12622_/C _12620_/Y vssd1 vssd1 vccd1 vccd1 _17595_/D sky130_fd_sc_hd__a21oi_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ _18676_/Q _18582_/Q _17537_/Q _17512_/Q _15262_/X _15301_/X vssd1 vssd1 vccd1
+ vccd1 _15341_/A sky130_fd_sc_hd__mux4_1
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ _12574_/B _12511_/X _14065_/B vssd1 vssd1 vccd1 vccd1 _12552_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11503_ _18043_/Q _11335_/A _11503_/S vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15271_ _19114_/Q _18945_/Q _18603_/Q _19343_/Q _15245_/X _09626_/A vssd1 vssd1 vccd1
+ vccd1 _15271_/X sky130_fd_sc_hd__mux4_1
X_12483_ _12476_/Y _12478_/Y _12480_/Y _12482_/Y _12408_/X _12560_/S vssd1 vssd1 vccd1
+ vccd1 _12762_/A sky130_fd_sc_hd__mux4_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14222_ _14222_/A vssd1 vssd1 vccd1 vccd1 _18081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11434_ _18100_/Q _11279_/X _11436_/S vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11365_ _11365_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11381_/S sky130_fd_sc_hd__or2_2
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18889_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03179_ clkbuf_0__03179_/X vssd1 vssd1 vccd1 vccd1 _14434__602/A sky130_fd_sc_hd__clkbuf_16
X_10316_ _09682_/X _18606_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _10317_/A sky130_fd_sc_hd__mux2_1
X_14084_ _12556_/X _14070_/X _14083_/Y _13343_/X vssd1 vssd1 vccd1 vccd1 _18011_/D
+ sky130_fd_sc_hd__a211o_1
X_18961_ _18961_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_1
X_11296_ _11296_/A vssd1 vssd1 vccd1 vccd1 _18158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13035_ _13035_/A vssd1 vssd1 vccd1 vccd1 _17689_/D sky130_fd_sc_hd__clkbuf_1
X_17912_ _19128_/CLK _17912_/D vssd1 vssd1 vccd1 vccd1 _17912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10247_ _10247_/A vssd1 vssd1 vccd1 vccd1 _18637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18892_ _18892_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17843_ _17935_/CLK _17843_/D vssd1 vssd1 vccd1 vccd1 _17843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10178_ _18694_/Q _10175_/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14367__549 _14367__549/A vssd1 vssd1 vccd1 vccd1 _18184_/CLK sky130_fd_sc_hd__inv_2
X_17774_ _17776_/CLK _17774_/D vssd1 vssd1 vccd1 vccd1 _17774_/Q sky130_fd_sc_hd__dfxtp_1
X_14986_ _18457_/Q _14986_/B vssd1 vssd1 vccd1 vccd1 _14998_/C sky130_fd_sc_hd__and2_1
Xclkbuf_0__04162_ _16067_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04162_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_235_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16725_ _17006_/A vssd1 vssd1 vccd1 vccd1 _16725_/X sky130_fd_sc_hd__buf_1
X_13937_ _13951_/A vssd1 vssd1 vccd1 vccd1 _13937_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _16584_/A vssd1 vssd1 vccd1 vccd1 _13868_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ _17648_/Q _17987_/Q _12822_/S vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__mux2_1
X_15607_ _18655_/Q _15612_/B vssd1 vssd1 vccd1 vccd1 _15607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16587_ _16613_/A _16587_/B _16587_/C vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__nor3_1
X_13799_ _17909_/Q _13796_/X _13798_/Y vssd1 vssd1 vccd1 vccd1 _17909_/D sky130_fd_sc_hd__o21a_1
XFILLER_76_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18326_ _19013_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
X_15538_ _15624_/A _15538_/B vssd1 vssd1 vccd1 vccd1 _18642_/D sky130_fd_sc_hd__nor2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420__109 _17420__109/A vssd1 vssd1 vccd1 vccd1 _19322_/CLK sky130_fd_sc_hd__inv_2
XFILLER_187_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15469_ _18670_/Q _18669_/Q vssd1 vssd1 vccd1 vccd1 _15643_/B sky130_fd_sc_hd__nor2_1
X_18257_ _18257_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ _17209_/B _17210_/A _17207_/Y vssd1 vssd1 vccd1 vccd1 _19244_/D sky130_fd_sc_hd__a21oi_1
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18188_ _18188_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17139_ _17142_/B _17142_/C vssd1 vssd1 vccd1 vccd1 _17140_/C sky130_fd_sc_hd__nand2_1
XFILLER_144_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _09961_/A vssd1 vssd1 vccd1 vccd1 _18777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08912_ _08945_/B _10372_/A vssd1 vssd1 vccd1 vccd1 _08942_/S sky130_fd_sc_hd__or2_2
X_14311__504 _14311__504/A vssd1 vssd1 vccd1 vccd1 _18139_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09895_/C _09892_/B _09892_/C vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__and3_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120__836 _15122__838/A vssd1 vssd1 vccd1 vccd1 _18512_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08843_ _08844_/A _09441_/A _08842_/Y vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__a21oi_1
XFILLER_112_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08774_ _08773_/X _18923_/Q vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__and2b_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14268__469 _14268__469/A vssd1 vssd1 vccd1 vccd1 _18104_/CLK sky130_fd_sc_hd__inv_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_74_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18465_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09326_ _19097_/Q _08952_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09257_ _10546_/A vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__buf_4
XFILLER_182_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09188_ _19163_/Q _09119_/X _09196_/S vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__mux2_1
X_14472__633 _14472__633/A vssd1 vssd1 vccd1 vccd1 _18268_/CLK sky130_fd_sc_hd__inv_2
XFILLER_182_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11150_ _11329_/A vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10101_ _10101_/A vssd1 vssd1 vccd1 vccd1 _18724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14171__449 _14171__449/A vssd1 vssd1 vccd1 vccd1 _18057_/CLK sky130_fd_sc_hd__inv_2
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11081_ _09047_/X _18245_/Q _11085_/S vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__mux2_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10032_ _18750_/Q _09935_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _14852_/A vssd1 vssd1 vccd1 vccd1 _14840_/X sky130_fd_sc_hd__buf_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16360__250 _16542__254/A vssd1 vssd1 vccd1 vccd1 _18966_/CLK sky130_fd_sc_hd__inv_2
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _14771_/A vssd1 vssd1 vccd1 vccd1 _14771_/X sky130_fd_sc_hd__buf_1
X_11983_ _19233_/Q vssd1 vssd1 vccd1 vccd1 _17169_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13722_ _13777_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13722_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__03797_ clkbuf_0__03797_/X vssd1 vssd1 vccd1 vccd1 _15407__907/A sky130_fd_sc_hd__clkbuf_16
X_16510_ _16511_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16514_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10934_ _10934_/A vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__clkbuf_1
X_17490_ _19326_/Q _17490_/B vssd1 vssd1 vccd1 vccd1 _17493_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13653_ _17860_/Q _13649_/X _13652_/Y vssd1 vssd1 vccd1 vccd1 _17860_/D sky130_fd_sc_hd__o21a_1
XFILLER_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16441_ _18970_/Q _16468_/B vssd1 vssd1 vccd1 vccd1 _16441_/Y sky130_fd_sc_hd__nand2_1
X_10865_ _18340_/Q _10809_/X _10867_/S vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12709_/B sky130_fd_sc_hd__buf_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ _19160_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_1
X_16372_ _17797_/Q _16382_/B vssd1 vssd1 vccd1 vccd1 _16383_/A sky130_fd_sc_hd__or2_1
X_13584_ _17840_/Q _13584_/B vssd1 vssd1 vccd1 vccd1 _13584_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10796_/A vssd1 vssd1 vccd1 vccd1 _18369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _18111_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_1
X_15323_ _18675_/Q _18581_/Q _17536_/Q _17511_/Q _15262_/X _15301_/X vssd1 vssd1 vccd1
+ vccd1 _15324_/A sky130_fd_sc_hd__mux4_1
X_12535_ _17628_/Q _12737_/A _17630_/Q _17631_/Q _12396_/X _12397_/X vssd1 vssd1 vccd1
+ vccd1 _12535_/X sky130_fd_sc_hd__mux4_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19091_ _19108_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03800_ _15417_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03800_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18042_ _18042_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15254_ _15246_/X _15247_/X _15250_/X _15253_/X _09600_/A _09625_/X vssd1 vssd1 vccd1
+ vccd1 _15254_/X sky130_fd_sc_hd__mux4_1
X_12466_ _17602_/Q _12647_/A _17604_/Q _12387_/X _12436_/S _12359_/A vssd1 vssd1 vccd1
+ vccd1 _12466_/X sky130_fd_sc_hd__mux4_2
XFILLER_184_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ _18074_/Q input32/X _14207_/S vssd1 vssd1 vccd1 vccd1 _14206_/A sky130_fd_sc_hd__mux2_1
X_11417_ _11417_/A vssd1 vssd1 vccd1 vccd1 _18108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15185_ _19137_/Q _19138_/Q _19139_/Q _19140_/Q _15626_/B _15626_/A vssd1 vssd1 vccd1
+ vccd1 _15185_/X sky130_fd_sc_hd__mux4_1
X_12397_ _12487_/S vssd1 vssd1 vccd1 vccd1 _12397_/X sky130_fd_sc_hd__buf_2
XFILLER_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14136_ _18031_/Q _14136_/B vssd1 vssd1 vccd1 vccd1 _14136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11348_ _11363_/S vssd1 vssd1 vccd1 vccd1 _11357_/S sky130_fd_sc_hd__buf_2
XFILLER_235_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14067_ _14055_/A _14067_/B vssd1 vssd1 vccd1 vccd1 _14067_/X sky130_fd_sc_hd__and2b_1
X_18944_ _18944_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03593_ _15124_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03593_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_234_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11279_ _18662_/Q vssd1 vssd1 vccd1 vccd1 _11279_/X sky130_fd_sc_hd__clkbuf_2
X_13018_ _17684_/Q _13092_/B vssd1 vssd1 vccd1 vccd1 _13019_/D sky130_fd_sc_hd__xor2_1
XFILLER_230_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18875_ _18888_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17826_ _17935_/CLK _17826_/D vssd1 vssd1 vccd1 vccd1 _17826_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17757_ _19290_/CLK _17757_/D vssd1 vssd1 vccd1 vccd1 _17757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14969_ _15026_/A _14967_/X _14979_/C vssd1 vssd1 vccd1 vccd1 _14970_/B sky130_fd_sc_hd__mux2_1
X_17408__99 _17408__99/A vssd1 vssd1 vccd1 vccd1 _19312_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17688_ _17945_/CLK _17688_/D vssd1 vssd1 vccd1 vccd1 _17688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16639_ _16639_/A vssd1 vssd1 vccd1 vccd1 _16639_/X sky130_fd_sc_hd__buf_1
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09111_ _18988_/Q vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__buf_4
X_18309_ _18309_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
X_19289_ _19290_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ _18664_/Q vssd1 vssd1 vccd1 vccd1 _11335_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _18781_/Q _09943_/X _09956_/S vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _16868_/A vssd1 vssd1 vccd1 vccd1 _09875_/X sky130_fd_sc_hd__buf_2
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_13 _10328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_24 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _19317_/Q _08801_/X _08828_/S vssd1 vssd1 vccd1 vccd1 _08827_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_35 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_46 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_57 _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_79 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _18933_/Q _09789_/B _08756_/X vssd1 vssd1 vccd1 vccd1 _08757_/X sky130_fd_sc_hd__a21o_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10650_ _09274_/X _18431_/Q _10654_/S vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _09309_/A vssd1 vssd1 vccd1 vccd1 _19105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10581_ _10581_/A vssd1 vssd1 vccd1 vccd1 _18492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12320_ _12320_/A vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__buf_1
XFILLER_182_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12251_ _12251_/A vssd1 vssd1 vccd1 vccd1 _17550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11202_ _18195_/Q _11065_/X _11202_/S vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__mux2_1
X_12182_ _12182_/A vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__clkbuf_2
X_15400__901 _15400__901/A vssd1 vssd1 vccd1 vccd1 _18588_/CLK sky130_fd_sc_hd__inv_2
XFILLER_218_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11133_ _11133_/A vssd1 vssd1 vccd1 vccd1 _18223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ _16892_/A _16989_/X _16860_/A vssd1 vssd1 vccd1 vccd1 _16990_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ _17816_/Q _15938_/A _17815_/Q vssd1 vssd1 vccd1 vccd1 _15943_/C sky130_fd_sc_hd__o21ai_1
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11064_ _11064_/A vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ _10015_/A vssd1 vssd1 vccd1 vccd1 _18758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _19144_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _17611_/CLK _17611_/D vssd1 vssd1 vccd1 vccd1 _17611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _18591_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _17542_/CLK _17542_/D vssd1 vssd1 vccd1 vccd1 _17542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11966_ _17250_/B _17252_/A _19257_/Q _17262_/B _11961_/X _11977_/S vssd1 vssd1 vccd1
+ vccd1 _11966_/X sky130_fd_sc_hd__mux4_2
XFILLER_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13705_ _13705_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__or2_2
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10917_ _18313_/Q _10892_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__mux2_1
X_17473_ _17473_/A vssd1 vssd1 vccd1 vccd1 _19338_/D sky130_fd_sc_hd__clkbuf_1
X_14685_ _18327_/Q _14543_/X _14623_/X _14684_/X vssd1 vssd1 vccd1 vccd1 _18327_/D
+ sky130_fd_sc_hd__o211a_1
X_11897_ _12008_/S vssd1 vssd1 vccd1 vccd1 _12032_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_232_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14479__639 _14479__639/A vssd1 vssd1 vccd1 vccd1 _18274_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19212_ _19212_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ _13636_/A vssd1 vssd1 vccd1 vccd1 _13636_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16424_ _16375_/Y _16376_/X _16379_/X _16421_/X _16423_/Y vssd1 vssd1 vccd1 vccd1
+ _16428_/C sky130_fd_sc_hd__a2111oi_4
X_10848_ _10848_/A vssd1 vssd1 vccd1 vccd1 _18348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19143_ _19143_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13567_ _13161_/X _13557_/B _13566_/Y _13555_/X vssd1 vssd1 vccd1 vccd1 _17834_/D
+ sky130_fd_sc_hd__a211oi_1
X_10779_ _18375_/Q _10701_/X _10781_/S vssd1 vssd1 vccd1 vccd1 _10780_/A sky130_fd_sc_hd__mux2_1
X_12518_ _18006_/Q vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15306_ _15298_/X _15300_/X _15304_/X _15305_/X vssd1 vssd1 vccd1 vccd1 _15306_/X
+ sky130_fd_sc_hd__o211a_1
X_16286_ _16284_/X _16285_/X _16286_/S vssd1 vssd1 vccd1 vccd1 _16286_/X sky130_fd_sc_hd__mux2_1
X_19074_ _19074_/CLK _19074_/D vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13498_ _13507_/S vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ _18029_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
X_12449_ _12446_/X _12447_/X _12449_/S vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ _09625_/X _15231_/X _15236_/Y vssd1 vssd1 vccd1 vccd1 _15237_/X sky130_fd_sc_hd__o21a_1
XFILLER_236_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _15168_/X sky130_fd_sc_hd__buf_1
XFILLER_158_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ _18023_/Q _14114_/X _14118_/Y vssd1 vssd1 vccd1 vccd1 _18023_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18927_ _18927_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09660_ _18912_/Q _09262_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09661_/A sky130_fd_sc_hd__mux2_1
X_18858_ _18858_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17809_ _19146_/CLK _17809_/D vssd1 vssd1 vccd1 vccd1 _17809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09591_ _18938_/Q _09495_/X _09591_/S vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__mux2_1
X_18789_ _18789_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__05077_ clkbuf_0__05077_/X vssd1 vssd1 vccd1 vccd1 _17409_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_150 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_161 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_172 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_183 _18882_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_194 _10175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15462__950 _15464__952/A vssd1 vssd1 vccd1 vccd1 _18637_/CLK sky130_fd_sc_hd__inv_2
XFILLER_148_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09025_ _09025_/A _11383_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _11024_/A sky130_fd_sc_hd__nand3_4
XFILLER_191_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16311__211 _16313__213/A vssd1 vssd1 vccd1 vccd1 _18927_/CLK sky130_fd_sc_hd__inv_2
XFILLER_163_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17003__352 _17005__354/A vssd1 vssd1 vccd1 vccd1 _19151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _09927_/A vssd1 vssd1 vccd1 vccd1 _18786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09858_ _09858_/A _18799_/Q _15808_/C vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__and3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ _10220_/A vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__buf_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09789_ _09789_/A _09789_/B _09377_/A vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__or3b_2
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _17929_/Q _11815_/X _11816_/X _11819_/X vssd1 vssd1 vccd1 vccd1 _11820_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11751_ _11751_/A vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15133__846 _15134__847/A vssd1 vssd1 vccd1 vccd1 _18522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10702_ _18407_/Q _10701_/X _10705_/S vssd1 vssd1 vccd1 vccd1 _10703_/A sky130_fd_sc_hd__mux2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _19024_/Q _19023_/Q _19022_/Q _16579_/A vssd1 vssd1 vccd1 vccd1 _16588_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_241_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ _13705_/A vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__clkbuf_4
X_10633_ _10633_/A vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _16171_/A _16140_/B vssd1 vssd1 vccd1 vccd1 _16140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13352_ _13645_/A _13352_/B vssd1 vssd1 vccd1 vccd1 _13541_/C sky130_fd_sc_hd__or2_1
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10564_ _10638_/B _10564_/B vssd1 vssd1 vccd1 vccd1 _10580_/S sky130_fd_sc_hd__or2_2
X_12303_ _17550_/Q _17490_/B vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__xnor2_1
XFILLER_155_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ _13281_/X _13282_/X _13275_/X vssd1 vssd1 vccd1 vccd1 _13283_/Y sky130_fd_sc_hd__a21oi_1
X_10495_ _10495_/A vssd1 vssd1 vccd1 vccd1 _18531_/D sky130_fd_sc_hd__clkbuf_1
X_15022_ _18463_/Q _14991_/X _15021_/Y _14993_/X vssd1 vssd1 vccd1 vccd1 _15023_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _12165_/A vssd1 vssd1 vccd1 vccd1 _17526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11116_ _18230_/Q _11056_/X _11116_/S vssd1 vssd1 vccd1 vccd1 _11117_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12096_ _19258_/Q _17264_/A _19260_/Q _19261_/Q _11995_/X _11938_/A vssd1 vssd1 vccd1
+ vccd1 _12096_/X sky130_fd_sc_hd__mux4_1
X_16973_ _19143_/Q _16797_/A _16972_/X _16915_/X vssd1 vssd1 vccd1 vccd1 _19143_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18712_ _18712_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_1
X_14485__643 _14486__644/A vssd1 vssd1 vccd1 vccd1 _18278_/CLK sky130_fd_sc_hd__inv_2
XFILLER_209_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _18667_/Q vssd1 vssd1 vccd1 vccd1 _11047_/X sky130_fd_sc_hd__buf_2
X_15924_ _18861_/Q vssd1 vssd1 vccd1 vccd1 _15967_/C sky130_fd_sc_hd__clkbuf_2
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16694__319 _16694__319/A vssd1 vssd1 vccd1 vccd1 _19094_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 io_in[19] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_4
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18643_ _18657_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03192_ clkbuf_0__03192_/X vssd1 vssd1 vccd1 vccd1 _14503__658/A sky130_fd_sc_hd__clkbuf_16
X_15855_ _15855_/A vssd1 vssd1 vccd1 vccd1 _15855_/X sky130_fd_sc_hd__buf_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18574_ _18922_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _15861_/A vssd1 vssd1 vccd1 vccd1 _15786_/X sky130_fd_sc_hd__buf_1
X_12998_ _12998_/A vssd1 vssd1 vccd1 vccd1 _17684_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17525_ _17878_/CLK _17525_/D vssd1 vssd1 vccd1 vccd1 _17525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14737_ _18592_/Q _18306_/Q _17572_/Q _18843_/Q _14579_/X _14641_/X vssd1 vssd1 vccd1
+ vccd1 _14737_/X sky130_fd_sc_hd__mux4_1
X_11949_ _19243_/Q _19244_/Q _12007_/S vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17398__90 _17399__91/A vssd1 vssd1 vccd1 vccd1 _19303_/CLK sky130_fd_sc_hd__inv_2
X_17456_ _17743_/Q _19333_/Q _17468_/S vssd1 vssd1 vccd1 vccd1 _17457_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14668_ _18407_/Q _18399_/Q _19312_/Q _17716_/Q _14594_/X _14595_/X vssd1 vssd1 vccd1
+ vccd1 _14668_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ _18970_/Q _16402_/B _16405_/Y _16437_/C _17808_/Q vssd1 vssd1 vccd1 vccd1
+ _16411_/B sky130_fd_sc_hd__a32o_1
XFILLER_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13619_ _13636_/A vssd1 vssd1 vccd1 vccd1 _13619_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_242_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14599_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__clkbuf_4
X_15407__907 _15407__907/A vssd1 vssd1 vccd1 vccd1 _18594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_158_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ _19126_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19057_ _19057_/CLK _19057_/D vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfxtp_1
X_16269_ _18781_/Q _18639_/Q _18789_/Q _18623_/Q _16158_/X _16182_/X vssd1 vssd1 vccd1
+ vccd1 _16269_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15792__114 _15792__114/A vssd1 vssd1 vccd1 vccd1 _18786_/CLK sky130_fd_sc_hd__inv_2
X_18008_ _18010_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04577_ clkbuf_0__04577_/X vssd1 vssd1 vccd1 vccd1 _16683_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09712_ _09691_/X _18892_/Q _09716_/S vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _09649_/C _09643_/B _09643_/C vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__and3_1
XFILLER_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798__731 _14799__732/A vssd1 vssd1 vccd1 vccd1 _18374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _18945_/Q _09498_/X _09578_/S vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ hold26/A _18802_/Q _09856_/C vssd1 vssd1 vccd1 vccd1 _09008_/X sky130_fd_sc_hd__and3_1
X_10280_ _18622_/Q _10183_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10281_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15690__988 _15691__989/A vssd1 vssd1 vccd1 vccd1 _18705_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13970_ _17968_/Q _13967_/X _13969_/Y vssd1 vssd1 vccd1 vccd1 _17968_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12921_ _12921_/A vssd1 vssd1 vccd1 vccd1 _12921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15640_ _16060_/A _15641_/B vssd1 vssd1 vccd1 vccd1 _18667_/D sky130_fd_sc_hd__nor2_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _17640_/Q _13094_/B vssd1 vssd1 vccd1 vccd1 _12859_/A sky130_fd_sc_hd__xor2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ input10/X _11790_/Y _11793_/X _17915_/Q _11802_/X vssd1 vssd1 vccd1 vccd1
+ _11803_/X sky130_fd_sc_hd__a221o_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12761_/X _12783_/B vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__and2b_1
X_15571_ _18649_/Q _15571_/B vssd1 vssd1 vccd1 vccd1 _15573_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17767_/Q _19276_/Q _17381_/B vssd1 vssd1 vccd1 vccd1 _17311_/B sky130_fd_sc_hd__mux2_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11734_/A vssd1 vssd1 vccd1 vccd1 _11734_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _18290_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16318__217 _16318__217/A vssd1 vssd1 vccd1 vccd1 _18933_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17246_/C _17265_/B _17241_/C vssd1 vssd1 vccd1 vccd1 _17242_/A sky130_fd_sc_hd__and3b_1
XFILLER_203_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11665_ _17510_/Q _09688_/A _11665_/S vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13404_ _13404_/A vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__buf_4
X_10616_ _10132_/X _18446_/Q _10618_/S vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__mux2_1
X_17172_ _17172_/A vssd1 vssd1 vccd1 vccd1 _19234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11596_ _11596_/A vssd1 vssd1 vccd1 vccd1 _17575_/D sky130_fd_sc_hd__clkbuf_1
XPeripherals_166 vssd1 vssd1 vccd1 vccd1 Peripherals_166/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_70_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPeripherals_177 vssd1 vssd1 vccd1 vccd1 Peripherals_177/HI io_out[3] sky130_fd_sc_hd__conb_1
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPeripherals_188 vssd1 vssd1 vccd1 vccd1 Peripherals_188/HI wb_data_o[27] sky130_fd_sc_hd__conb_1
X_13335_ _13237_/X _13330_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13335_/Y sky130_fd_sc_hd__a21oi_1
X_16123_ _18743_/Q _18751_/Q _18759_/Q _18767_/Q _16198_/A _16172_/A vssd1 vssd1 vccd1
+ vccd1 _16123_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10547_ _10562_/S vssd1 vssd1 vccd1 vccd1 _10556_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15856__155 _15860__159/A vssd1 vssd1 vccd1 vccd1 _18830_/CLK sky130_fd_sc_hd__inv_2
X_13266_ _13265_/X _13259_/X _13260_/X vssd1 vssd1 vccd1 vccd1 _13266_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _16054_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _18880_/D sky130_fd_sc_hd__nor2_1
X_10478_ _18538_/Q _10333_/X _10484_/S vssd1 vssd1 vccd1 vccd1 _10479_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12217_ _12217_/A _12217_/B _12217_/C _12217_/D vssd1 vssd1 vccd1 vccd1 _12218_/C
+ sky130_fd_sc_hd__or4_1
X_15005_ _15005_/A _15005_/B vssd1 vssd1 vccd1 vccd1 _15014_/C sky130_fd_sc_hd__and2_1
XFILLER_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13197_ _14081_/A vssd1 vssd1 vccd1 vccd1 _16057_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ _12148_/A vssd1 vssd1 vccd1 vccd1 _17521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03413_ _14833_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03413_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ _12214_/A _12186_/A _12180_/A _12181_/A vssd1 vssd1 vccd1 vccd1 _12079_/X
+ sky130_fd_sc_hd__and4b_1
X_16956_ _18153_/Q _18145_/Q _18137_/Q _18281_/Q _16809_/X _16810_/X vssd1 vssd1 vccd1
+ vccd1 _16956_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15907_ _18874_/Q _15907_/B vssd1 vssd1 vccd1 vccd1 _15945_/B sky130_fd_sc_hd__xor2_1
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16887_ _09868_/X _16885_/X _16886_/X vssd1 vssd1 vccd1 vccd1 _16887_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_225_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18626_ _18626_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03175_ clkbuf_0__03175_/X vssd1 vssd1 vccd1 vccd1 _14417__589/A sky130_fd_sc_hd__clkbuf_16
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18557_ _18993_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _17508_/CLK _17508_/D vssd1 vssd1 vccd1 vccd1 _17508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09290_ _09290_/A vssd1 vssd1 vccd1 vccd1 _19117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18488_ _18488_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17439_ _17748_/Q _19328_/Q _17451_/S vssd1 vssd1 vccd1 vccd1 _17440_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19109_ _19109_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_99_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18987_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput110 _11755_/X vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_2
XFILLER_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput121 _11715_/X vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_2
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput132 _19397_/X vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__buf_2
XFILLER_217_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19337_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput143 _11801_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[0] sky130_fd_sc_hd__buf_2
Xoutput154 _11808_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_114_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09626_ _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__and2_1
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09557_ _09557_/A vssd1 vssd1 vccd1 vccd1 _18953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15772__1054 _15772__1054/A vssd1 vssd1 vccd1 vccd1 _18771_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09488_ _09488_/A vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__03402_ clkbuf_0__03402_/X vssd1 vssd1 vccd1 vccd1 _14802_/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f__07170_ clkbuf_0__07170_/X vssd1 vssd1 vccd1 vccd1 _11881__364/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11450_ _18093_/Q _11276_/X _11454_/S vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14436__604 _14436__604/A vssd1 vssd1 vccd1 vccd1 _18239_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ _16198_/A vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__clkbuf_4
X_17392__85 _17396__89/A vssd1 vssd1 vccd1 vccd1 _19298_/CLK sky130_fd_sc_hd__inv_2
X_11381_ _11344_/X _18123_/Q _11381_/S vssd1 vssd1 vccd1 vccd1 _11382_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03195_ clkbuf_0__03195_/X vssd1 vssd1 vccd1 vccd1 _14517__669/A sky130_fd_sc_hd__clkbuf_16
XFILLER_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ _10332_/A vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13051_ _13049_/X _13051_/B vssd1 vssd1 vccd1 vccd1 _13052_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _10263_/A vssd1 vssd1 vccd1 vccd1 _18630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12002_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12087_/S sky130_fd_sc_hd__buf_2
XFILLER_106_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10194_ _10194_/A vssd1 vssd1 vccd1 vccd1 _18689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16810_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16810_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17790_ _17923_/CLK _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16741_ _19129_/Q _19136_/Q _16741_/S vssd1 vssd1 vccd1 vccd1 _16741_/X sky130_fd_sc_hd__mux2_1
X_13953_ _13964_/B vssd1 vssd1 vccd1 vccd1 _13962_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _12904_/A vssd1 vssd1 vccd1 vccd1 _17664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _17937_/Q _13878_/X _13883_/Y vssd1 vssd1 vccd1 vccd1 _17937_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _19040_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15623_ _15621_/X _15622_/Y _15626_/B vssd1 vssd1 vccd1 vccd1 _15624_/B sky130_fd_sc_hd__mux2_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ input30/X vssd1 vssd1 vccd1 vccd1 _19391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_234_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12835_ _12835_/A vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__buf_2
XFILLER_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18342_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15554_ _15551_/X _15552_/Y _15553_/X vssd1 vssd1 vccd1 vccd1 _18645_/D sky130_fd_sc_hd__a21oi_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A vssd1 vssd1 vccd1 vccd1 _12766_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261__464 _14261__464/A vssd1 vssd1 vccd1 vccd1 _18099_/CLK sky130_fd_sc_hd__inv_2
XFILLER_187_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _14505_/A vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__buf_1
X_11717_ _11869_/B vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__clkbuf_2
X_18273_ _18273_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12707_/C _12697_/B vssd1 vssd1 vccd1 vccd1 _17616_/D sky130_fd_sc_hd__nor2_1
X_15485_ _18655_/Q _15485_/B vssd1 vssd1 vccd1 vccd1 _15485_/X sky130_fd_sc_hd__xor2_1
XFILLER_203_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17224_ _17225_/B _17222_/A _17223_/Y vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ _11648_/A vssd1 vssd1 vccd1 vccd1 _17535_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03962_ _15649_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03962_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 io_in[22] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_4
XFILLER_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput23 jtag_tdo vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_2
XFILLER_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput34 wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
X_17155_ _17158_/B _17162_/D vssd1 vssd1 vccd1 vccd1 _17156_/C sky130_fd_sc_hd__or2_1
Xinput45 wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_2
XFILLER_155_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11579_ _17582_/Q _10907_/X _11581_/S vssd1 vssd1 vccd1 vccd1 _11580_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03793_ clkbuf_0__03793_/X vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__clkbuf_16
Xinput56 wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput67 wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_6
XFILLER_156_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput78 wb_stb_i vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_4
X_16106_ _16195_/A vssd1 vssd1 vccd1 vccd1 _16106_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13318_ _13268_/X _13311_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _13318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16037_ _16037_/A vssd1 vssd1 vccd1 vccd1 _18876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13249_ _17744_/Q _13219_/X _13248_/Y vssd1 vssd1 vccd1 vccd1 _17744_/D sky130_fd_sc_hd__o21a_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08790_ _19346_/Q _08789_/X _08796_/S vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__mux2_1
X_17988_ _19247_/CLK _17988_/D vssd1 vssd1 vccd1 vccd1 _17988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04376_ _16347_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04376_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16939_ _19209_/Q _19161_/Q _18272_/Q _18264_/Q _16882_/A _16868_/X vssd1 vssd1 vccd1
+ vccd1 _16939_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _09411_/A vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _18609_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03158_ clkbuf_0__03158_/X vssd1 vssd1 vccd1 vccd1 _14330__519/A sky130_fd_sc_hd__clkbuf_16
XFILLER_213_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09342_ _19090_/Q _09223_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03189_ _14481_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03189_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03089_ clkbuf_0__03089_/X vssd1 vssd1 vccd1 vccd1 _14141__426/A sky130_fd_sc_hd__clkbuf_16
X_12344__404 _12344__404/A vssd1 vssd1 vccd1 vccd1 _17585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_221_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09273_ _09273_/A vssd1 vssd1 vccd1 vccd1 _19123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _19212_/Q _08967_/X _08988_/S vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10950_ hold9/A vssd1 vssd1 vccd1 vccd1 _10959_/S sky130_fd_sc_hd__buf_2
XFILLER_84_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09609_ _15301_/A vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10881_ _18333_/Q _10806_/X _10885_/S vssd1 vssd1 vccd1 vccd1 _10882_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12620_ _12622_/B _12622_/C _12607_/X vssd1 vssd1 vccd1 vccd1 _12620_/Y sky130_fd_sc_hd__o21ai_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12551_ _12511_/X _18004_/Q _12351_/X _12838_/A vssd1 vssd1 vccd1 vccd1 _12563_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _11502_/A vssd1 vssd1 vccd1 vccd1 _18044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ _12482_/A vssd1 vssd1 vccd1 vccd1 _12482_/Y sky130_fd_sc_hd__clkinv_2
X_15270_ _16064_/A vssd1 vssd1 vccd1 vccd1 _15270_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14221_ _18081_/Q input39/X _14229_/S vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__mux2_1
X_11433_ _11433_/A vssd1 vssd1 vccd1 vccd1 _18101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11364_ _11364_/A vssd1 vssd1 vccd1 vccd1 _18131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03178_ clkbuf_0__03178_/X vssd1 vssd1 vccd1 vccd1 _14430__599/A sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13103_ _13103_/A vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__buf_1
X_10315_ _10315_/A vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__clkbuf_1
X_14083_ _14083_/A _14083_/B vssd1 vssd1 vccd1 vccd1 _14083_/Y sky130_fd_sc_hd__nor2_2
X_18960_ _18960_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ _18158_/Q _11273_/X _11295_/S vssd1 vssd1 vccd1 vccd1 _11296_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13034_ _13032_/X _13034_/B vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__and2b_1
X_17911_ _19128_/CLK _17911_/D vssd1 vssd1 vccd1 vccd1 _17911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10246_ _18637_/Q _10186_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _10247_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18891_ _18891_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17842_ _17935_/CLK _17842_/D vssd1 vssd1 vccd1 vccd1 _17842_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10177_ _10199_/S vssd1 vssd1 vccd1 vccd1 _10190_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17773_ _17776_/CLK _17773_/D vssd1 vssd1 vccd1 vccd1 _17773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14985_ _18457_/Q _14986_/B vssd1 vssd1 vccd1 vccd1 _14987_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13936_ _17956_/Q _13941_/B vssd1 vssd1 vccd1 vccd1 _13936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13867_ input65/X _13867_/B vssd1 vssd1 vccd1 vccd1 _13867_/X sky130_fd_sc_hd__and2_1
XFILLER_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15606_ _15611_/A _15606_/B _15610_/B vssd1 vssd1 vccd1 vccd1 _15606_/X sky130_fd_sc_hd__or3_1
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12818_ _12818_/A vssd1 vssd1 vccd1 vccd1 _17647_/D sky130_fd_sc_hd__clkbuf_1
X_16586_ _19022_/Q _16585_/C _19023_/Q vssd1 vssd1 vccd1 vccd1 _16587_/C sky130_fd_sc_hd__a21oi_1
X_13798_ _13394_/X _13797_/X _13789_/X vssd1 vssd1 vccd1 vccd1 _13798_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18325_ _19013_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
X_15537_ _15551_/A _15615_/B _15543_/C vssd1 vssd1 vccd1 vccd1 _15538_/B sky130_fd_sc_hd__mux2_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ _12758_/D _12749_/B vssd1 vssd1 vccd1 vccd1 _17632_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18256_ _18256_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15468_ _15581_/A vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__buf_2
XFILLER_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16667__302 _16669__304/A vssd1 vssd1 vccd1 vccd1 _19076_/CLK sky130_fd_sc_hd__inv_2
X_17207_ _17209_/B _17210_/A _17191_/X vssd1 vssd1 vccd1 vccd1 _17207_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14419_ _14425_/A vssd1 vssd1 vccd1 vccd1 _14419_/X sky130_fd_sc_hd__buf_1
XFILLER_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18187_ _18187_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _17142_/B _17142_/C vssd1 vssd1 vccd1 vccd1 _17140_/B sky130_fd_sc_hd__or2_1
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _18777_/Q _09959_/X _09968_/S vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08911_ _09648_/A _08911_/B _08889_/B vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__or3b_4
X_15771__1053 _15771__1053/A vssd1 vssd1 vccd1 vccd1 _18770_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _10583_/B _09891_/B vssd1 vssd1 vccd1 vccd1 _09892_/C sky130_fd_sc_hd__or2_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _19050_/Q hold15/A vssd1 vssd1 vccd1 vccd1 _08842_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_246_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08773_ _08773_/A _08773_/B _08773_/C vssd1 vssd1 vccd1 vccd1 _08773_/X sky130_fd_sc_hd__and3_1
XFILLER_111_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15869__165 _15872__168/A vssd1 vssd1 vccd1 vccd1 _18840_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17036__29 _17036__29/A vssd1 vssd1 vccd1 vccd1 _19178_/CLK sky130_fd_sc_hd__inv_2
XFILLER_211_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14506__660 _14510__664/A vssd1 vssd1 vccd1 vccd1 _18295_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09325_ _09325_/A vssd1 vssd1 vccd1 vccd1 _19098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _10432_/A _09256_/B _09936_/C vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__or3_4
XFILLER_22_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_opt_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19252_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ _09202_/S vssd1 vssd1 vccd1 vccd1 _09196_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_193_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _18724_/Q _10057_/X _10104_/S vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__mux2_1
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11080_ _11080_/A vssd1 vssd1 vccd1 vccd1 _18246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _10046_/S vssd1 vssd1 vccd1 vccd1 _10040_/S sky130_fd_sc_hd__buf_2
XFILLER_248_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11982_ _17142_/A _11978_/X _19229_/Q _17158_/B _11980_/X _11981_/X vssd1 vssd1 vccd1
+ vccd1 _11982_/X sky130_fd_sc_hd__mux4_2
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03796_ clkbuf_0__03796_/X vssd1 vssd1 vccd1 vccd1 _15403__904/A sky130_fd_sc_hd__clkbuf_16
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13721_ _13735_/B vssd1 vssd1 vccd1 vccd1 _13733_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10933_ _18306_/Q _10887_/X _10941_/S vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14891__806 _14892__807/A vssd1 vssd1 vccd1 vccd1 _18451_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16440_ _16440_/A vssd1 vssd1 vccd1 vccd1 _16468_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_231_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13652_ _13649_/X _13707_/A _13532_/X vssd1 vssd1 vccd1 vccd1 _13652_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10864_ _10864_/A vssd1 vssd1 vccd1 vccd1 _18341_/D sky130_fd_sc_hd__clkbuf_1
X_14407__580 _14411__584/A vssd1 vssd1 vccd1 vccd1 _18215_/CLK sky130_fd_sc_hd__inv_2
XFILLER_231_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12603_ _17591_/Q _12603_/B vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__or2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _17798_/Q _16389_/B vssd1 vssd1 vccd1 vccd1 _16382_/B sky130_fd_sc_hd__or2_1
X_13583_ _16058_/A _13574_/B _13582_/Y _13569_/X vssd1 vssd1 vccd1 vccd1 _17839_/D
+ sky130_fd_sc_hd__a211oi_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10795_ _18369_/Q _10794_/X _10804_/S vssd1 vssd1 vccd1 vccd1 _10796_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ _18110_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15322_ _18832_/Q _18824_/Q _18816_/Q _18683_/Q _15299_/X _15225_/X vssd1 vssd1 vccd1
+ vccd1 _15322_/X sky130_fd_sc_hd__mux4_2
XFILLER_223_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12534_ _12528_/Y _12529_/Y _12532_/Y _12533_/Y _12586_/S _12504_/A vssd1 vssd1 vccd1
+ vccd1 _12845_/A sky130_fd_sc_hd__mux4_2
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _19090_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18041_ _18041_/CLK _18041_/D vssd1 vssd1 vccd1 vccd1 _18041_/Q sky130_fd_sc_hd__dfxtp_1
X_15253_ _18936_/Q _18899_/Q _18891_/Q _18845_/Q _15251_/X _15252_/X vssd1 vssd1 vccd1
+ vccd1 _15253_/X sky130_fd_sc_hd__mux4_1
X_12465_ _12631_/A _17599_/Q _17600_/Q _12383_/X _12436_/S _12359_/A vssd1 vssd1 vccd1
+ vccd1 _12465_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204_ _14204_/A vssd1 vssd1 vccd1 vccd1 _18073_/D sky130_fd_sc_hd__clkbuf_1
X_11416_ _11341_/X _18108_/Q _11418_/S vssd1 vssd1 vccd1 vccd1 _11417_/A sky130_fd_sc_hd__mux2_1
X_12396_ _12432_/S vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_193_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15184_ _18659_/Q vssd1 vssd1 vccd1 vccd1 _15626_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14373__554 _14373__554/A vssd1 vssd1 vccd1 vccd1 _18189_/CLK sky130_fd_sc_hd__inv_2
X_14750__692 _14752__694/A vssd1 vssd1 vccd1 vccd1 _18335_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _13147_/B _13434_/X _14134_/Y _11697_/X vssd1 vssd1 vccd1 vccd1 _18030_/D
+ sky130_fd_sc_hd__a211oi_1
X_11347_ _11493_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11363_/S sky130_fd_sc_hd__nor2_2
XFILLER_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03592_ _15118_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03592_/X sky130_fd_sc_hd__clkbuf_16
X_14066_ input73/X _16518_/B _14054_/X _14065_/X _13343_/X vssd1 vssd1 vccd1 vccd1
+ _18004_/D sky130_fd_sc_hd__a311o_1
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18943_ _18943_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_1
X_11278_ _11278_/A vssd1 vssd1 vccd1 vccd1 _18165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16662__298 _16663__299/A vssd1 vssd1 vccd1 vccd1 _19072_/CLK sky130_fd_sc_hd__inv_2
X_13017_ _17675_/Q _13095_/B vssd1 vssd1 vccd1 vccd1 _13019_/C sky130_fd_sc_hd__xnor2_1
X_10229_ _10229_/A vssd1 vssd1 vccd1 vccd1 _18675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18874_ _18879_/CLK _18874_/D vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17825_ _19146_/CLK _17825_/D vssd1 vssd1 vccd1 vccd1 _17825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17756_ _19290_/CLK _17756_/D vssd1 vssd1 vccd1 vccd1 _17756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14968_ _18454_/Q vssd1 vssd1 vccd1 vccd1 _14979_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16707_ _16707_/A vssd1 vssd1 vccd1 vccd1 _16707_/X sky130_fd_sc_hd__buf_1
XFILLER_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13919_ _17950_/Q _13903_/X _13918_/Y vssd1 vssd1 vccd1 vccd1 _17950_/D sky130_fd_sc_hd__o21a_1
X_17687_ _17703_/CLK _17687_/D vssd1 vssd1 vccd1 vccd1 _17687_/Q sky130_fd_sc_hd__dfxtp_1
X_14899_ _17855_/Q _17854_/Q _14942_/B vssd1 vssd1 vccd1 vccd1 _14930_/A sky130_fd_sc_hd__or3_2
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14792__726 _14793__727/A vssd1 vssd1 vccd1 vccd1 _18369_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16569_ _16578_/A _16569_/B _16569_/C vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__nor3_1
XFILLER_149_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09110_ _09110_/A vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18308_ _18308_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19288_ _19288_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12228__374 _12228__374/A vssd1 vssd1 vccd1 vccd1 _17538_/CLK sky130_fd_sc_hd__inv_2
X_09041_ _09041_/A vssd1 vssd1 vccd1 vccd1 _19208_/D sky130_fd_sc_hd__clkbuf_1
X_18239_ _18239_/CLK _18239_/D vssd1 vssd1 vccd1 vccd1 _18239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14274__474 _14274__474/A vssd1 vssd1 vccd1 vccd1 _18109_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09943_ _10117_/A vssd1 vssd1 vccd1 vccd1 _09943_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _09874_/A _09874_/B vssd1 vssd1 vccd1 vccd1 _18808_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08825_ _08825_/A vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_14 _10333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_25 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_36 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_47 _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_58 _17908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_69 _19388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ _18934_/Q hold10/A vssd1 vssd1 vccd1 vccd1 _08756_/X sky130_fd_sc_hd__xor2_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ _08921_/X _19105_/Q _09312_/S vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__mux2_1
X_10580_ _10135_/X _18492_/Q _10580_/S vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09239_ _09972_/A _18559_/Q _10403_/B _09238_/Y vssd1 vssd1 vccd1 vccd1 _09247_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_194_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12250_ _12245_/X _12250_/B vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__and2b_1
XFILLER_154_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ _11201_/A vssd1 vssd1 vccd1 vccd1 _18196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12181_ _12181_/A vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__buf_2
XFILLER_123_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11132_ _18223_/Q _11053_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _11133_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15654__959 _15654__959/A vssd1 vssd1 vccd1 vccd1 _18676_/CLK sky130_fd_sc_hd__inv_2
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11063_ _18252_/Q _11062_/X _11066_/S vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__mux2_1
X_15940_ _18869_/Q _15940_/B vssd1 vssd1 vccd1 vccd1 _15940_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _18758_/Q _09935_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__mux2_1
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _17618_/CLK _17610_/D vssd1 vssd1 vccd1 vccd1 _17610_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _18590_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17541_ _17541_/CLK _17541_/D vssd1 vssd1 vccd1 vccd1 _17541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14759_/A vssd1 vssd1 vccd1 vccd1 _14753_/X sky130_fd_sc_hd__buf_1
XFILLER_229_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11965_ _19258_/Q vssd1 vssd1 vccd1 vccd1 _17262_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13704_ _14053_/B _13704_/B vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__nand2_1
XFILLER_233_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17472_ _16736_/A _17472_/B vssd1 vssd1 vccd1 vccd1 _17473_/A sky130_fd_sc_hd__and2b_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10916_ _10916_/A vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14684_ _14544_/X _14673_/X _14683_/Y vssd1 vssd1 vccd1 vccd1 _14684_/X sky130_fd_sc_hd__a21o_1
XFILLER_225_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ _17780_/Q vssd1 vssd1 vccd1 vccd1 _12008_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19211_ _19211_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16423_ _18983_/Q _16423_/B vssd1 vssd1 vccd1 vccd1 _16423_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_204_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13635_ _17857_/Q _13635_/B vssd1 vssd1 vccd1 vccd1 _13635_/Y sky130_fd_sc_hd__nor2_1
X_14856__778 _14857__779/A vssd1 vssd1 vccd1 vccd1 _18423_/CLK sky130_fd_sc_hd__inv_2
X_15770__1052 _15771__1053/A vssd1 vssd1 vccd1 vccd1 _18769_/CLK sky130_fd_sc_hd__inv_2
X_10847_ _18348_/Q _10809_/X _10849_/S vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19142_ _19143_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
X_13566_ _17834_/Q _13568_/B vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10778_ _10778_/A vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12517_ _12517_/A vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__buf_2
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19073_ _19073_/CLK _19073_/D vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16285_ _18718_/Q _18726_/Q _18734_/Q _18499_/Q _16205_/X _16206_/X vssd1 vssd1 vccd1
+ vccd1 _16285_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13599_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13507_/S sky130_fd_sc_hd__nor2_2
XFILLER_185_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18024_ _18024_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ _09614_/A _15235_/Y _09600_/A vssd1 vssd1 vccd1 vccd1 _15236_/Y sky130_fd_sc_hd__a21oi_1
X_12448_ _12448_/A vssd1 vssd1 vccd1 vccd1 _12449_/S sky130_fd_sc_hd__buf_2
XFILLER_161_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _12377_/X _12378_/X _12390_/S vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14118_ _13400_/A _14115_/X _14108_/X vssd1 vssd1 vccd1 vccd1 _14118_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_236_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _13812_/X _14039_/X _14046_/X vssd1 vssd1 vccd1 vccd1 _14049_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18926_ _18926_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18857_ _18857_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09590_ _09590_/A vssd1 vssd1 vccd1 vccd1 _18939_/D sky130_fd_sc_hd__clkbuf_1
X_17808_ _19108_/CLK _17808_/D vssd1 vssd1 vccd1 vccd1 _17808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18788_ _18788_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17739_ _19337_/CLK _17739_/D vssd1 vssd1 vccd1 vccd1 _17739_/Q sky130_fd_sc_hd__dfxtp_1
X_14800__733 _14801__734/A vssd1 vssd1 vccd1 vccd1 _18376_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__05076_ clkbuf_0__05076_/X vssd1 vssd1 vccd1 vccd1 _17386__81/A sky130_fd_sc_hd__clkbuf_16
XFILLER_211_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17014__10 _17016__12/A vssd1 vssd1 vccd1 vccd1 _19159_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_140 _11804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_151 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_162 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_173 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_184 _18884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_195 _10336_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14757__698 _14757__698/A vssd1 vssd1 vccd1 vccd1 _18341_/CLK sky130_fd_sc_hd__inv_2
XFILLER_149_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09024_ hold22/X vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09926_ _18786_/Q _09271_/X _09926_/S vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09857_/A _09857_/B _09857_/C _09004_/Y vssd1 vssd1 vccd1 vccd1 _15808_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08808_ _08889_/B _09648_/A _08911_/B vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__or3_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _09788_/A vssd1 vssd1 vccd1 vccd1 _18836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _08746_/B vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11750_ _17861_/Q _19340_/Q _17771_/Q vssd1 vssd1 vccd1 vccd1 _11751_/A sky130_fd_sc_hd__mux2_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10701_ _10701_/A vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11681_ _19021_/Q _19020_/Q _19019_/Q _16571_/A vssd1 vssd1 vccd1 vccd1 _16579_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ _19147_/Q _13420_/B vssd1 vssd1 vccd1 vccd1 _13705_/A sky130_fd_sc_hd__nand2_2
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10632_ _18439_/Q _10129_/A _10636_/S vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13351_ _13623_/A vssd1 vssd1 vccd1 vccd1 _14069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10563_ _10563_/A vssd1 vssd1 vccd1 vccd1 _18500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _17558_/Q _17491_/B vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__xnor2_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14519__670 _14520__671/A vssd1 vssd1 vccd1 vccd1 _18305_/CLK sky130_fd_sc_hd__inv_2
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13282_ _13288_/A vssd1 vssd1 vccd1 vccd1 _13282_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10494_ _10112_/X _18531_/Q _10502_/S vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15021_ _15021_/A _15031_/C vssd1 vssd1 vccd1 vccd1 _15021_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ _12149_/X _12164_/B vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__and2b_1
XFILLER_68_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11115_ _11115_/A vssd1 vssd1 vccd1 vccd1 _18231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12095_ _12095_/A vssd1 vssd1 vccd1 vccd1 _12199_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16972_ _16892_/X _16961_/X _16971_/Y vssd1 vssd1 vccd1 vccd1 _16972_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18711_ _18711_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_1
X_15923_ _15970_/A _15929_/B _15923_/C vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__and3_1
X_11046_ _11046_/A vssd1 vssd1 vccd1 vccd1 _18258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15889__179 _15889__179/A vssd1 vssd1 vccd1 vccd1 _18855_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18642_ _18657_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03191_ clkbuf_0__03191_/X vssd1 vssd1 vccd1 vccd1 _14496__652/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _18922_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15785_ _15785_/A vssd1 vssd1 vccd1 vccd1 _15785_/X sky130_fd_sc_hd__buf_1
X_12997_ _12992_/X _12997_/B vssd1 vssd1 vccd1 vccd1 _12998_/A sky130_fd_sc_hd__and2b_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _19329_/CLK _17524_/D vssd1 vssd1 vccd1 vccd1 _17524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _14736_/A _14736_/B vssd1 vssd1 vccd1 vccd1 _14736_/Y sky130_fd_sc_hd__nor2_1
XFILLER_229_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11948_ _17781_/Q vssd1 vssd1 vccd1 vccd1 _12007_/S sky130_fd_sc_hd__buf_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17455_ _17474_/S vssd1 vssd1 vccd1 vccd1 _17468_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _19176_/Q _19168_/Q _19200_/Q _18335_/Q _14591_/X _14592_/X vssd1 vssd1 vccd1
+ vccd1 _14667_/X sky130_fd_sc_hd__mux4_2
XFILLER_177_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16406_ _18968_/Q vssd1 vssd1 vccd1 vccd1 _16437_/C sky130_fd_sc_hd__clkbuf_2
X_13618_ _17851_/Q _13621_/B vssd1 vssd1 vccd1 vccd1 _13618_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _18364_/Q _18316_/Q _18372_/Q _17705_/Q _14637_/A _14569_/X vssd1 vssd1 vccd1
+ vccd1 _14598_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19125_ _19125_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _13568_/B vssd1 vssd1 vccd1 vccd1 _13549_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_203_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19056_ _19056_/CLK _19056_/D vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfxtp_1
X_16076__191 _16077__192/A vssd1 vssd1 vccd1 vccd1 _18896_/CLK sky130_fd_sc_hd__inv_2
XFILLER_145_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16268_ _18631_/Q _18506_/Q _18912_/Q _18514_/Q _16155_/X _16156_/X vssd1 vssd1 vccd1
+ vccd1 _16268_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18007_ _18007_/CLK _18007_/D vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_2
X_15219_ _18935_/Q _18898_/Q _18890_/Q _18844_/Q _15209_/X _15218_/X vssd1 vssd1 vccd1
+ vccd1 _15219_/X sky130_fd_sc_hd__mux4_1
X_16199_ _18440_/Q _18690_/Q _18698_/Q _18706_/Q _16198_/X _16172_/X vssd1 vssd1 vccd1
+ vccd1 _16200_/B sky130_fd_sc_hd__mux4_1
XFILLER_142_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04576_ clkbuf_0__04576_/X vssd1 vssd1 vccd1 vccd1 _16675__309/A sky130_fd_sc_hd__clkbuf_16
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09711_ _09711_/A vssd1 vssd1 vccd1 vccd1 _18893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18909_ _18909_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09642_ _10219_/C _09647_/A vssd1 vssd1 vccd1 vccd1 _09643_/C sky130_fd_sc_hd__or2_1
XFILLER_56_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09573_ _09573_/A vssd1 vssd1 vccd1 vccd1 _18946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ _18809_/Q hold22/A vssd1 vssd1 vccd1 vccd1 _09856_/C sky130_fd_sc_hd__xnor2_1
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14807__739 _14807__739/A vssd1 vssd1 vccd1 vccd1 _18382_/CLK sky130_fd_sc_hd__inv_2
XFILLER_247_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09909_ _18793_/Q _09735_/X _09913_/S vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12920_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _17650_/Q _13092_/B _12850_/X _17636_/Q vssd1 vssd1 vccd1 vccd1 _12860_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11802_/A vssd1 vssd1 vccd1 vccd1 _11802_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15568_/X _15569_/Y _15553_/X vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__a21oi_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12782_ _17637_/Q _17998_/Q _12862_/B vssd1 vssd1 vccd1 vccd1 _12783_/B sky130_fd_sc_hd__mux2_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _17769_/Q _17933_/Q vssd1 vssd1 vccd1 vccd1 _11734_/A sky130_fd_sc_hd__and2b_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _19253_/Q _17240_/B vssd1 vssd1 vccd1 vccd1 _17241_/C sky130_fd_sc_hd__or2_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11664_ _11664_/A vssd1 vssd1 vccd1 vccd1 _17511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13403_ _16741_/S vssd1 vssd1 vccd1 vccd1 _16767_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17171_ _17169_/X _17171_/B _17191_/A vssd1 vssd1 vccd1 vccd1 _17172_/A sky130_fd_sc_hd__and3b_1
XFILLER_31_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10615_ _10615_/A vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328__390 _12329__391/A vssd1 vssd1 vccd1 vccd1 _17571_/CLK sky130_fd_sc_hd__inv_2
X_11595_ _17575_/Q _10707_/A _11599_/S vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__mux2_1
XPeripherals_167 vssd1 vssd1 vccd1 vccd1 Peripherals_167/HI io_oeb[30] sky130_fd_sc_hd__conb_1
XFILLER_128_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPeripherals_178 vssd1 vssd1 vccd1 vccd1 Peripherals_178/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16122_ _18568_/Q vssd1 vssd1 vccd1 vccd1 _16234_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13334_ _17770_/Q _13329_/X _13333_/Y vssd1 vssd1 vccd1 vccd1 _17770_/D sky130_fd_sc_hd__o21a_1
XFILLER_41_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPeripherals_189 vssd1 vssd1 vccd1 vccd1 Peripherals_189/HI wb_data_o[28] sky130_fd_sc_hd__conb_1
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10546_ _10546_/A _10546_/B vssd1 vssd1 vccd1 vccd1 _10562_/S sky130_fd_sc_hd__nor2_2
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16053_ _16061_/B vssd1 vssd1 vccd1 vccd1 _16058_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13265_ _14081_/A vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__buf_6
XFILLER_124_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10477_ _10477_/A vssd1 vssd1 vccd1 vccd1 _18539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__05079_ clkbuf_0__05079_/X vssd1 vssd1 vccd1 vccd1 _17399__91/A sky130_fd_sc_hd__clkbuf_16
X_15004_ _15005_/A _15005_/B vssd1 vssd1 vccd1 vccd1 _15006_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_0__04530_ _16556_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04530_/X sky130_fd_sc_hd__clkbuf_16
X_12216_ _17515_/Q _12180_/A _12298_/A _17529_/Q _12215_/X vssd1 vssd1 vccd1 vccd1
+ _12217_/D sky130_fd_sc_hd__a221o_1
XFILLER_29_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13196_ _13411_/A vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12147_ _12132_/X _12147_/B vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__and2b_1
XFILLER_229_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03412_ _14827_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03412_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12078_ _12022_/A _12073_/X _12075_/Y _12077_/Y vssd1 vssd1 vccd1 vccd1 _12181_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_16955_ _18121_/Q _18113_/Q _18105_/Q _18097_/Q _16893_/X _16894_/X vssd1 vssd1 vccd1
+ vccd1 _16955_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11029_ _11029_/A vssd1 vssd1 vccd1 vccd1 _18265_/D sky130_fd_sc_hd__clkbuf_1
X_15906_ _15951_/A _15906_/B vssd1 vssd1 vccd1 vccd1 _15907_/B sky130_fd_sc_hd__nand2_1
X_16886_ _16902_/A vssd1 vssd1 vccd1 vccd1 _16886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15413__912 _15413__912/A vssd1 vssd1 vccd1 vccd1 _18599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_225_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15837_ _15843_/A vssd1 vssd1 vccd1 vccd1 _15837_/X sky130_fd_sc_hd__buf_1
X_18625_ _18625_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03174_ clkbuf_0__03174_/X vssd1 vssd1 vccd1 vccd1 _14410__583/A sky130_fd_sc_hd__clkbuf_16
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18556_ _18921_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15667__969 _15667__969/A vssd1 vssd1 vccd1 vccd1 _18686_/CLK sky130_fd_sc_hd__inv_2
XFILLER_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14719_ _14640_/X _14718_/X _14604_/A vssd1 vssd1 vccd1 vccd1 _14719_/Y sky130_fd_sc_hd__o21ai_1
X_17507_ _17507_/CLK _17507_/D vssd1 vssd1 vccd1 vccd1 _17507_/Q sky130_fd_sc_hd__dfxtp_1
X_18487_ _18487_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_1
X_15699_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15699_/X sky130_fd_sc_hd__buf_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17438_ _17474_/S vssd1 vssd1 vccd1 vccd1 _17451_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14500__655 _14504__659/A vssd1 vssd1 vccd1 vccd1 _18290_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17369_ _17364_/Y _17365_/X _17366_/X _17368_/X vssd1 vssd1 vccd1 vccd1 _17369_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_242_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19108_ _19108_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19039_/CLK _19039_/D vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput100 _11711_/X vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_133_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput111 _11751_/X vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_2
Xoutput122 _11713_/X vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_2
Xoutput133 _18801_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput144 _11838_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput155 _11811_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_115_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _17953_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09625_ _15307_/A vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09556_ _08933_/X _18953_/Q _09560_/S vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03401_ clkbuf_0__03401_/X vssd1 vssd1 vccd1 vccd1 _14773__711/A sky130_fd_sc_hd__clkbuf_16
XFILLER_52_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09487_ _19011_/Q _09486_/X _09496_/S vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401__575 _14403__577/A vssd1 vssd1 vccd1 vccd1 _18210_/CLK sky130_fd_sc_hd__inv_2
XFILLER_221_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10400_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16198_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14813__743 _14813__743/A vssd1 vssd1 vccd1 vccd1 _18386_/CLK sky130_fd_sc_hd__inv_2
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11380_ _11380_/A vssd1 vssd1 vccd1 vccd1 _18124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03194_ clkbuf_0__03194_/X vssd1 vssd1 vccd1 vccd1 _14536_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10331_ _18600_/Q _10328_/X _10343_/S vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ _17944_/Q _17694_/Q _13053_/S vssd1 vssd1 vccd1 vccd1 _13051_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10262_ _18630_/Q _10183_/X _10266_/S vssd1 vssd1 vccd1 vccd1 _10263_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12001_ _17274_/B _17276_/A _17279_/A _19264_/Q _11931_/S _12017_/S vssd1 vssd1 vccd1
+ vccd1 _12001_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10193_ _18689_/Q _10192_/X _10199_/S vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16740_ _16740_/A vssd1 vssd1 vccd1 vccd1 _16740_/Y sky130_fd_sc_hd__inv_2
X_16324__222 _16326__224/A vssd1 vssd1 vccd1 vccd1 _18938_/CLK sky130_fd_sc_hd__inv_2
X_13952_ _16060_/A _13946_/X _13950_/Y _13951_/X vssd1 vssd1 vccd1 vccd1 _17961_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12903_ _12894_/X _12903_/B vssd1 vssd1 vccd1 vccd1 _12904_/A sky130_fd_sc_hd__and2b_1
X_13883_ _13285_/X _13879_/X _13880_/X vssd1 vssd1 vccd1 vccd1 _13883_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15622_ _15642_/A _15622_/B vssd1 vssd1 vccd1 vccd1 _15622_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18410_ _18410_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19390_ input29/X vssd1 vssd1 vccd1 vccd1 _19390_/X sky130_fd_sc_hd__clkbuf_1
X_12834_ _12834_/A vssd1 vssd1 vccd1 vccd1 _12834_/X sky130_fd_sc_hd__buf_2
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18341_ _18341_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15553_ _15581_/A vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12433_/X _12418_/X _12765_/S vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04579_ clkbuf_0__04579_/X vssd1 vssd1 vccd1 vccd1 _16694__319/A sky130_fd_sc_hd__clkbuf_16
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11716_ _17783_/Q vssd1 vssd1 vccd1 vccd1 _11869_/B sky130_fd_sc_hd__buf_2
X_18272_ _18272_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15529_/B _15484_/B vssd1 vssd1 vccd1 vccd1 _15485_/B sky130_fd_sc_hd__nand2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _17616_/Q _12693_/A _12695_/X vssd1 vssd1 vccd1 vccd1 _12697_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17223_ _17225_/B _17222_/A _17191_/X vssd1 vssd1 vccd1 vccd1 _17223_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_230_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _08795_/X _17535_/Q _11647_/S vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 io_in[23] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_8
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ _17158_/B _17162_/D vssd1 vssd1 vccd1 vccd1 _17159_/B sky130_fd_sc_hd__and2_1
XFILLER_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput24 vga_b[0] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_8
Xinput35 wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11578_ _11578_/A vssd1 vssd1 vccd1 vccd1 _17583_/D sky130_fd_sc_hd__clkbuf_1
Xinput46 wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_2
XFILLER_155_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput57 wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_4
X_16105_ _16194_/A vssd1 vssd1 vccd1 vccd1 _16171_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ _17765_/Q _13303_/X _13316_/Y vssd1 vssd1 vccd1 vccd1 _17765_/D sky130_fd_sc_hd__o21a_1
Xinput79 wb_we_i vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_4
X_10529_ _10544_/S vssd1 vssd1 vccd1 vccd1 _10538_/S sky130_fd_sc_hd__clkbuf_2
X_15146__857 _15148__859/A vssd1 vssd1 vccd1 vccd1 _18533_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222__369 _12222__369/A vssd1 vssd1 vccd1 vccd1 _17533_/CLK sky130_fd_sc_hd__inv_2
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _16036_/A _16036_/B _16036_/C _16036_/D vssd1 vssd1 vccd1 vccd1 _16037_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13248_ _13247_/X _13232_/A _13241_/X vssd1 vssd1 vccd1 vccd1 _13248_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16626__269 _16626__269/A vssd1 vssd1 vccd1 vccd1 _19043_/CLK sky130_fd_sc_hd__inv_2
X_13179_ _14074_/A vssd1 vssd1 vccd1 vccd1 _16060_/A sky130_fd_sc_hd__buf_12
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _19247_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 _17987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048__38 _17048__38/A vssd1 vssd1 vccd1 vccd1 _19187_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__04375_ _16341_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04375_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16938_ _16936_/X _16937_/X _16976_/S vssd1 vssd1 vccd1 vccd1 _16938_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _19206_/Q _19158_/Q _18269_/Q _18261_/Q _16882_/A _16868_/X vssd1 vssd1 vccd1
+ vccd1 _16869_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09410_ _08937_/X _19060_/Q _09412_/S vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18608_ _18608_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03157_ clkbuf_0__03157_/X vssd1 vssd1 vccd1 vccd1 _14349_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _09356_/S vssd1 vssd1 vccd1 vccd1 _09350_/S sky130_fd_sc_hd__buf_2
XFILLER_206_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03188_ _14480_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03188_/X sky130_fd_sc_hd__clkbuf_16
X_18539_ _18539_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498__654 _14498__654/A vssd1 vssd1 vccd1 vccd1 _18289_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09272_ _19123_/Q _09271_/X _09272_/S vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _08987_/A vssd1 vssd1 vccd1 vccd1 _19213_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09608_ _15208_/A vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_204_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10880_ _10880_/A vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09539_ _09539_/A vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__clkbuf_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _12775_/D vssd1 vssd1 vccd1 vccd1 _12838_/A sky130_fd_sc_hd__buf_2
XFILLER_197_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14399__574 _14399__574/A vssd1 vssd1 vccd1 vccd1 _18209_/CLK sky130_fd_sc_hd__inv_2
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11501_ _18044_/Q _11332_/A _11503_/S vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _12403_/X _12386_/X _12547_/S vssd1 vssd1 vccd1 vccd1 _12482_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14220_ _14231_/A vssd1 vssd1 vccd1 vccd1 _14229_/S sky130_fd_sc_hd__clkbuf_2
X_11432_ _18101_/Q _11276_/X _11436_/S vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _14151_/A vssd1 vssd1 vccd1 vccd1 _14151_/X sky130_fd_sc_hd__buf_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ _18131_/Q _11282_/X _11363_/S vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03177_ clkbuf_0__03177_/X vssd1 vssd1 vccd1 vccd1 _14423__593/A sky130_fd_sc_hd__clkbuf_16
X_10314_ _09679_/X _18607_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__mux2_1
X_14082_ _12449_/S _14070_/X _14081_/Y _13343_/X vssd1 vssd1 vccd1 vccd1 _18010_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11294_ _11294_/A vssd1 vssd1 vccd1 vccd1 _18159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13033_ _17949_/Q _17689_/Q _13099_/B vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__mux2_1
X_17910_ _18007_/CLK _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545__256 _16548__259/A vssd1 vssd1 vccd1 vccd1 _19002_/CLK sky130_fd_sc_hd__inv_2
X_10245_ _10245_/A vssd1 vssd1 vccd1 vccd1 _18638_/D sky130_fd_sc_hd__clkbuf_1
X_18890_ _18890_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17841_ _17935_/CLK _17841_/D vssd1 vssd1 vccd1 vccd1 _17841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10176_ _10546_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10199_/S sky130_fd_sc_hd__nor2_2
XFILLER_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17772_ _17772_/CLK _17772_/D vssd1 vssd1 vccd1 vccd1 _17772_/Q sky130_fd_sc_hd__dfxtp_1
X_14984_ _14984_/A vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14744__689 _14744__689/A vssd1 vssd1 vccd1 vccd1 _18332_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13935_ _13146_/X _13925_/X _13934_/Y _13636_/X vssd1 vssd1 vccd1 vccd1 _17955_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13866_ _17933_/Q _13863_/B _13865_/X _13857_/X vssd1 vssd1 vccd1 vccd1 _17933_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_207_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15605_ _18655_/Q _18654_/Q _15605_/C vssd1 vssd1 vccd1 vccd1 _15610_/B sky130_fd_sc_hd__and3_1
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12817_ _12812_/X _12817_/B vssd1 vssd1 vccd1 vccd1 _12818_/A sky130_fd_sc_hd__and2b_1
X_16585_ _19023_/Q _19022_/Q _16585_/C vssd1 vssd1 vccd1 vccd1 _16587_/B sky130_fd_sc_hd__and3_1
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13797_ _13802_/A vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15536_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15615_/B sky130_fd_sc_hd__inv_2
X_18324_ _19013_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
X_12748_ _12746_/A _12745_/A _12734_/X vssd1 vssd1 vccd1 vccd1 _12749_/B sky130_fd_sc_hd__o21ai_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18255_ _18255_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
X_15467_ _15470_/A vssd1 vssd1 vccd1 vccd1 _15581_/A sky130_fd_sc_hd__clkbuf_2
X_12679_ _12679_/A _12679_/B vssd1 vssd1 vccd1 vccd1 _17611_/D sky130_fd_sc_hd__nor2_1
XFILLER_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17206_ _17210_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _19243_/D sky130_fd_sc_hd__nor2_1
XFILLER_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14418_ _14449_/A vssd1 vssd1 vccd1 vccd1 _14418_/X sky130_fd_sc_hd__buf_1
XFILLER_163_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18186_ _18186_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ _15410_/A vssd1 vssd1 vccd1 vccd1 _15398_/X sky130_fd_sc_hd__buf_1
XFILLER_144_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17137_ _17137_/A vssd1 vssd1 vccd1 vccd1 _19225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14349_ _14349_/A vssd1 vssd1 vccd1 vccd1 _14349_/X sky130_fd_sc_hd__buf_1
XFILLER_116_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17068_ _17068_/A vssd1 vssd1 vccd1 vccd1 _17068_/X sky130_fd_sc_hd__buf_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08910_ _09674_/A vssd1 vssd1 vccd1 vccd1 _08910_/X sky130_fd_sc_hd__clkbuf_4
X_16019_ _16024_/A _16019_/B _16027_/C vssd1 vssd1 vccd1 vccd1 _16019_/X sky130_fd_sc_hd__or3_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09894_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__and2_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08841_ _09446_/A hold12/A vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__and2_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08772_/A _08772_/B _08772_/C vssd1 vssd1 vccd1 vccd1 _08773_/C sky130_fd_sc_hd__nor3_1
XFILLER_100_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09324_ _19098_/Q _08949_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15088__811 _15089__812/A vssd1 vssd1 vccd1 vccd1 _18487_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ _09255_/A _09970_/A vssd1 vssd1 vccd1 vccd1 _09936_/C sky130_fd_sc_hd__nand2_1
XFILLER_193_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15426__922 _15428__924/A vssd1 vssd1 vccd1 vccd1 _18609_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09186_ _11024_/A _11260_/A vssd1 vssd1 vccd1 vccd1 _09202_/S sky130_fd_sc_hd__nor2_4
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_83_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18657_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14513__665 _14514__666/A vssd1 vssd1 vccd1 vccd1 _18300_/CLK sky130_fd_sc_hd__inv_2
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19108_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _10620_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10046_/S sky130_fd_sc_hd__nor2_2
XFILLER_88_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15095__815 _15095__815/A vssd1 vssd1 vccd1 vccd1 _18491_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11981_ _12005_/S vssd1 vssd1 vccd1 vccd1 _11981_/X sky130_fd_sc_hd__buf_2
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _17883_/Q _13715_/X _13719_/Y _13710_/X vssd1 vssd1 vccd1 vccd1 _17883_/D
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__03795_ clkbuf_0__03795_/X vssd1 vssd1 vccd1 vccd1 _15395__897/A sky130_fd_sc_hd__clkbuf_16
X_10932_ hold16/A vssd1 vssd1 vccd1 vccd1 _10941_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13651_ input64/X _16532_/B vssd1 vssd1 vccd1 vccd1 _13707_/A sky130_fd_sc_hd__nand2_2
XFILLER_232_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10863_ _18341_/Q _10806_/X _10867_/S vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ _12614_/D vssd1 vssd1 vccd1 vccd1 _12610_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _17800_/Q _17799_/Q _16393_/B vssd1 vssd1 vccd1 vccd1 _16389_/B sky130_fd_sc_hd__or3_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13582_ _17839_/Q _13584_/B vssd1 vssd1 vccd1 vccd1 _13582_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _10794_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15321_ _15317_/X _15318_/X _15319_/X _15320_/X _15281_/X _09600_/X vssd1 vssd1 vccd1
+ vccd1 _15321_/X sky130_fd_sc_hd__mux4_1
X_12533_ _12533_/A vssd1 vssd1 vccd1 vccd1 _12533_/Y sky130_fd_sc_hd__clkinv_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16551__260 _16552__261/A vssd1 vssd1 vccd1 vccd1 _19006_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _18040_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
X_15252_ _15291_/A vssd1 vssd1 vccd1 vccd1 _15252_/X sky130_fd_sc_hd__clkbuf_2
X_12464_ _12375_/X _12377_/X _12464_/S vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14203_ _18073_/Q input53/X _14207_/S vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _11415_/A vssd1 vssd1 vccd1 vccd1 _18109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15183_ _18658_/Q vssd1 vssd1 vccd1 vccd1 _15626_/B sky130_fd_sc_hd__clkbuf_2
X_12395_ _17595_/Q vssd1 vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _18030_/Q _14134_/B vssd1 vssd1 vccd1 vccd1 _14134_/Y sky130_fd_sc_hd__nor2_1
X_11346_ _11346_/A vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070__186 _16071__187/A vssd1 vssd1 vccd1 vccd1 _18891_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _14055_/A _14065_/B vssd1 vssd1 vccd1 vccd1 _14065_/X sky130_fd_sc_hd__and2b_1
X_18942_ _18942_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03591_ _15112_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03591_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11277_ _18165_/Q _11276_/X _11283_/S vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__mux2_1
X_13016_ _17679_/Q _13093_/B vssd1 vssd1 vccd1 vccd1 _13019_/B sky130_fd_sc_hd__xnor2_1
XFILLER_140_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10228_ _18675_/Q _09755_/X _10230_/S vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__mux2_1
X_18873_ _18879_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17824_ _19146_/CLK _17824_/D vssd1 vssd1 vccd1 vccd1 _17824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _18702_/Q _10048_/X _10167_/S vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17755_ _19290_/CLK _17755_/D vssd1 vssd1 vccd1 vccd1 _17755_/Q sky130_fd_sc_hd__dfxtp_1
X_14967_ _14991_/A vssd1 vssd1 vccd1 vccd1 _14967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13918_ _13812_/X _13908_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13918_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17686_ _17963_/CLK _17686_/D vssd1 vssd1 vccd1 vccd1 _17686_/Q sky130_fd_sc_hd__dfxtp_1
X_14898_ _17859_/Q _17858_/Q _17857_/Q _17856_/Q vssd1 vssd1 vccd1 vccd1 _14942_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _14243_/A _13849_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__nand2_2
XFILLER_223_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17041__33 _17042__34/A vssd1 vssd1 vccd1 vccd1 _19182_/CLK sky130_fd_sc_hd__inv_2
X_16568_ _16567_/A _19016_/Q _19017_/Q vssd1 vssd1 vccd1 vccd1 _16569_/C sky130_fd_sc_hd__a21oi_1
XFILLER_204_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18307_ _18307_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15519_ _15517_/B _15517_/C _15557_/B vssd1 vssd1 vccd1 vccd1 _15523_/B sky130_fd_sc_hd__a21oi_1
X_19287_ _19287_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
X_16499_ _18982_/Q _16499_/B vssd1 vssd1 vccd1 vccd1 _16499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_241_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09040_ _09039_/X _19208_/Q _09044_/S vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__mux2_1
X_18238_ _18238_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18169_ _18169_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15875__170 _15878__173/A vssd1 vssd1 vccd1 vccd1 _18845_/CLK sky130_fd_sc_hd__inv_2
XFILLER_239_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09942_ _18479_/Q vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__buf_4
XFILLER_143_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09873_ _09869_/A _09869_/B _09870_/X vssd1 vssd1 vccd1 vccd1 _09874_/B sky130_fd_sc_hd__o21ai_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _19318_/Q _08798_/X _08828_/S vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_15 _16578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_26 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_37 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15159__867 _15161__869/A vssd1 vssd1 vccd1 vccd1 _18543_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_48 _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_59 _17890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08755_ hold1/X vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__inv_2
XFILLER_39_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ _09307_/A vssd1 vssd1 vccd1 vccd1 _19106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09238_ _09238_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _09238_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09169_ _09184_/S vssd1 vssd1 vccd1 vccd1 _09178_/S sky130_fd_sc_hd__buf_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17502__9 _17502__9/A vssd1 vssd1 vccd1 vccd1 _19344_/CLK sky130_fd_sc_hd__inv_2
X_11200_ _18196_/Q _11062_/X _11202_/S vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12180_ _12180_/A vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ _11131_/A vssd1 vssd1 vccd1 vccd1 _18224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15103__822 _15103__822/A vssd1 vssd1 vccd1 vccd1 _18498_/CLK sky130_fd_sc_hd__inv_2
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _18662_/Q vssd1 vssd1 vccd1 vccd1 _11062_/X sky130_fd_sc_hd__buf_2
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _10028_/S vssd1 vssd1 vccd1 vccd1 _10022_/S sky130_fd_sc_hd__buf_2
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14821_/X sky130_fd_sc_hd__buf_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17540_ _17540_/CLK _17540_/D vssd1 vssd1 vccd1 vccd1 _17540_/Q sky130_fd_sc_hd__dfxtp_1
X_11964_ _19256_/Q vssd1 vssd1 vccd1 vccd1 _17252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _17878_/Q _13683_/X _13702_/Y vssd1 vssd1 vccd1 vccd1 _17878_/D sky130_fd_sc_hd__o21a_1
X_14147__431 _14149__433/A vssd1 vssd1 vccd1 vccd1 _18039_/CLK sky130_fd_sc_hd__inv_2
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _17738_/Q _19338_/Q _17474_/S vssd1 vssd1 vccd1 vccd1 _17472_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10915_ _18314_/Q _10887_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ _14664_/A _14682_/X _14619_/X vssd1 vssd1 vccd1 vccd1 _14683_/Y sky130_fd_sc_hd__o21ai_1
X_11895_ _17225_/C _19249_/Q _11924_/S vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19210_ _19210_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13634_ _13192_/X _13626_/B _13633_/Y _13619_/X vssd1 vssd1 vccd1 vccd1 _17856_/D
+ sky130_fd_sc_hd__a211oi_1
X_16422_ _17794_/Q _16422_/B vssd1 vssd1 vccd1 vccd1 _16423_/B sky130_fd_sc_hd__or2_1
X_10846_ _10846_/A vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16353_ _16359_/A vssd1 vssd1 vccd1 vccd1 _16353_/X sky130_fd_sc_hd__buf_1
X_19141_ _19143_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13565_ _13155_/X _13549_/X _13564_/Y _13555_/X vssd1 vssd1 vccd1 vccd1 _17833_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10777_ _18376_/Q _10698_/X _10781_/S vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15304_ _15304_/A _15303_/X vssd1 vssd1 vccd1 vccd1 _15304_/X sky130_fd_sc_hd__or2b_1
X_12516_ _12580_/A _12512_/X _12515_/X vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__o21ai_1
XFILLER_200_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19072_ _19072_/CLK _19072_/D vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16284_ _18750_/Q _18758_/Q _18766_/Q _18774_/Q _16149_/X _16150_/X vssd1 vssd1 vccd1
+ vccd1 _16284_/X sky130_fd_sc_hd__mux4_1
X_13496_ _17810_/Q _13490_/Y _13495_/Y vssd1 vssd1 vccd1 vccd1 _17810_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18023_ _18027_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _15235_/A vssd1 vssd1 vccd1 vccd1 _15235_/Y sky130_fd_sc_hd__clkinv_2
X_12447_ _12626_/A _12631_/A _17599_/Q _12638_/A _12443_/X _12429_/S vssd1 vssd1 vccd1
+ vccd1 _12447_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12378_ _17614_/Q _17615_/Q _12443_/A vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04592_ clkbuf_0__04592_/X vssd1 vssd1 vccd1 vccd1 _16735__348/A sky130_fd_sc_hd__clkbuf_16
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _18022_/Q _14114_/X _14116_/Y vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__o21a_1
XFILLER_113_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11329_ _11329_/A vssd1 vssd1 vccd1 vccd1 _11329_/X sky130_fd_sc_hd__buf_2
XFILLER_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14048_ _17997_/Q _14033_/X _14047_/Y vssd1 vssd1 vccd1 vccd1 _17997_/D sky130_fd_sc_hd__o21a_1
XFILLER_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18925_ _18925_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18856_ _18856_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17807_ _19108_/CLK _17807_/D vssd1 vssd1 vccd1 vccd1 _17807_/Q sky130_fd_sc_hd__dfxtp_1
X_18787_ _18787_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_1
X_15999_ _16002_/B _16020_/B vssd1 vssd1 vccd1 vccd1 _15999_/Y sky130_fd_sc_hd__nand2_1
X_17738_ _19339_/CLK _17738_/D vssd1 vssd1 vccd1 vccd1 _17738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16558__266 _16558__266/A vssd1 vssd1 vccd1 vccd1 _19012_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_130 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17669_ _18006_/CLK _17669_/D vssd1 vssd1 vccd1 vccd1 _17669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_141 _11804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_152 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_163 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_174 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_185 _18078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_196 _10789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _19339_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09023_ _11068_/B vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _09925_/A vssd1 vssd1 vccd1 vccd1 _18787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _09010_/X _09856_/B _09856_/C vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__nand3b_1
XFILLER_219_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08807_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _08911_/B sky130_fd_sc_hd__nand2_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _08886_/X _18836_/Q _09787_/S vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08738_ _18090_/Q _18089_/Q vssd1 vssd1 vccd1 vccd1 _08746_/B sky130_fd_sc_hd__or2_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10700_/A vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11680_ _19015_/Q _19018_/Q _19017_/Q _19016_/Q vssd1 vssd1 vccd1 vccd1 _16571_/A
+ sky130_fd_sc_hd__and4_1
X_17010__358 _17011__359/A vssd1 vssd1 vccd1 vccd1 _19157_/CLK sky130_fd_sc_hd__inv_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _10631_/A vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13350_ _14243_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__nand2_4
XFILLER_22_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10562_ _18500_/Q _10135_/A _10562_/S vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__mux2_1
X_15660__964 _15660__964/A vssd1 vssd1 vccd1 vccd1 _18681_/CLK sky130_fd_sc_hd__inv_2
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12301_ _12301_/A _12301_/B _12301_/C vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__and3_1
X_13281_ _13434_/A vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__buf_4
X_10493_ _10508_/S vssd1 vssd1 vccd1 vccd1 _10502_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15020_ _18463_/Q _15020_/B vssd1 vssd1 vccd1 vccd1 _15031_/C sky130_fd_sc_hd__and2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12163_ _17526_/Q _17725_/Q _12170_/S vssd1 vssd1 vccd1 vccd1 _12164_/B sky130_fd_sc_hd__mux2_1
XFILLER_155_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11114_ _18231_/Q _11053_/X _11116_/S vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12094_ _11945_/X _12090_/X _12093_/X vssd1 vssd1 vccd1 vccd1 _12095_/A sky130_fd_sc_hd__o21ai_1
X_16971_ _16892_/A _16970_/X _16860_/A vssd1 vssd1 vccd1 vccd1 _16971_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_231_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18710_ _18710_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ _15929_/B _15923_/C _15970_/A vssd1 vssd1 vccd1 vccd1 _15922_/Y sky130_fd_sc_hd__a21oi_1
X_11045_ _18258_/Q _11042_/X _11057_/S vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__mux2_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862__783 _14862__783/A vssd1 vssd1 vccd1 vccd1 _18428_/CLK sky130_fd_sc_hd__inv_2
XFILLER_237_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _19144_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03190_ clkbuf_0__03190_/X vssd1 vssd1 vccd1 vccd1 _14490__647/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _18572_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12996_ _17953_/Q _17684_/Q _12999_/S vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__mux2_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17523_ _17737_/CLK _17523_/D vssd1 vssd1 vccd1 vccd1 _17523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11947_ _11947_/A vssd1 vssd1 vccd1 vccd1 _17490_/B sky130_fd_sc_hd__buf_4
X_14735_ _17588_/Q _18386_/Q _18394_/Q _18428_/Q _14574_/X _14637_/X vssd1 vssd1 vccd1
+ vccd1 _14736_/B sky130_fd_sc_hd__mux4_2
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15826__131 _15826__131/A vssd1 vssd1 vccd1 vccd1 _18806_/CLK sky130_fd_sc_hd__inv_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _17454_/A vssd1 vssd1 vccd1 vccd1 _17454_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14666_ _18326_/Q _14543_/X _14623_/X _14665_/Y vssd1 vssd1 vccd1 vccd1 _18326_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13617_ _13155_/X _13601_/X _13616_/Y _13604_/X vssd1 vssd1 vccd1 vccd1 _17850_/D
+ sky130_fd_sc_hd__a211oi_1
X_16405_ _17808_/Q _17807_/Q _17806_/Q vssd1 vssd1 vccd1 vccd1 _16405_/Y sky130_fd_sc_hd__o21ai_1
X_10829_ _18356_/Q _10809_/X _10831_/S vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14597_ _14593_/X _14596_/X _14688_/S vssd1 vssd1 vccd1 vccd1 _14597_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ _19124_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ _13559_/S vssd1 vssd1 vccd1 vccd1 _13568_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_146_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14492__649 _14492__649/A vssd1 vssd1 vccd1 vccd1 _18284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ _16265_/X _16266_/X _16286_/S vssd1 vssd1 vccd1 vccd1 _16267_/X sky130_fd_sc_hd__mux2_1
X_19055_ _19055_/CLK _19055_/D vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfxtp_1
X_13479_ input66/X _13483_/B vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__and2_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _18006_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15218_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15218_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16198_ _16198_/A vssd1 vssd1 vccd1 vccd1 _16198_/X sky130_fd_sc_hd__buf_2
XFILLER_142_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15149_ _15149_/A vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__buf_1
XFILLER_236_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04575_ clkbuf_0__04575_/X vssd1 vssd1 vccd1 vccd1 _16669__304/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09710_ _09688_/X _18893_/Q _09710_/S vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__mux2_1
X_18908_ _18908_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09641_ _09641_/A vssd1 vssd1 vccd1 vccd1 _18928_/D sky130_fd_sc_hd__clkbuf_1
X_18839_ _18839_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09572_ _18946_/Q _09495_/X _09572_/S vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04009_ clkbuf_0__04009_/X vssd1 vssd1 vccd1 vccd1 _15851__151/A sky130_fd_sc_hd__clkbuf_16
XFILLER_196_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14393__569 _14393__569/A vssd1 vssd1 vccd1 vccd1 _18204_/CLK sky130_fd_sc_hd__inv_2
X_09006_ _09001_/Y hold25/A _09011_/A _09004_/Y vssd1 vssd1 vccd1 vccd1 _09006_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09908_ _09908_/A vssd1 vssd1 vccd1 vccd1 _18794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09839_ _09839_/A vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12850_ _12850_/A vssd1 vssd1 vccd1 vccd1 _12850_/X sky130_fd_sc_hd__buf_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _17935_/Q _11785_/X _11797_/X _11800_/X vssd1 vssd1 vccd1 vccd1 _11801_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_215_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12781_/A vssd1 vssd1 vccd1 vccd1 _17636_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17819_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_215_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11663_ _17511_/Q _09685_/A _11665_/S vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__mux2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13402_ _17786_/Q vssd1 vssd1 vccd1 vccd1 _16741_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_17170_ _17169_/B _17169_/C _17173_/B vssd1 vssd1 vccd1 vccd1 _17171_/B sky130_fd_sc_hd__a21o_1
X_10614_ _10129_/X _18447_/Q _10618_/S vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11594_ _11594_/A vssd1 vssd1 vccd1 vccd1 _17576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16121_ _10406_/A _16104_/Y _16110_/Y _16114_/Y _16120_/Y vssd1 vssd1 vccd1 vccd1
+ _16121_/X sky130_fd_sc_hd__o32a_2
XPeripherals_168 vssd1 vssd1 vccd1 vccd1 Peripherals_168/HI io_oeb[31] sky130_fd_sc_hd__conb_1
X_13333_ _13146_/X _13330_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13333_/Y sky130_fd_sc_hd__a21oi_1
XPeripherals_179 vssd1 vssd1 vccd1 vccd1 Peripherals_179/HI io_out[5] sky130_fd_sc_hd__conb_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10545_ _10545_/A vssd1 vssd1 vccd1 vccd1 _18508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15895__184 _15895__184/A vssd1 vssd1 vccd1 vccd1 _18860_/CLK sky130_fd_sc_hd__inv_2
X_16052_ _16052_/A _16294_/B _16052_/C vssd1 vssd1 vccd1 vccd1 _16061_/B sky130_fd_sc_hd__nand3_4
X_13264_ _17748_/Q _13252_/X _13263_/Y vssd1 vssd1 vccd1 vccd1 _17748_/D sky130_fd_sc_hd__o21a_1
XFILLER_155_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10476_ _18539_/Q _10328_/X _10484_/S vssd1 vssd1 vccd1 vccd1 _10477_/A sky130_fd_sc_hd__mux2_1
X_15003_ _15080_/B vssd1 vssd1 vccd1 vccd1 _15034_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__05078_ clkbuf_0__05078_/X vssd1 vssd1 vccd1 vccd1 _17396__89/A sky130_fd_sc_hd__clkbuf_16
X_12215_ _17520_/Q _17478_/B vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__xor2_1
X_17416__105 _17420__109/A vssd1 vssd1 vccd1 vccd1 _19318_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ input67/X _13483_/B vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12146_ _17521_/Q _17730_/Q _12153_/S vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03411_ _14821_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03411_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_238_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12077_ _12098_/S _12076_/X _12069_/A vssd1 vssd1 vccd1 vccd1 _12077_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16954_ _19142_/Q _16797_/A _16953_/X _16915_/X vssd1 vssd1 vccd1 vccd1 _19142_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11028_ _18265_/Q _09127_/X _11034_/S vssd1 vssd1 vccd1 vccd1 _11029_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15905_ _17812_/Q _15947_/A vssd1 vssd1 vccd1 vccd1 _15906_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ _18213_/Q _18197_/Q _18486_/Q _18189_/Q _16834_/X _09875_/X vssd1 vssd1 vccd1
+ vccd1 _16885_/X sky130_fd_sc_hd__mux4_1
X_18624_ _18624_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03173_ clkbuf_0__03173_/X vssd1 vssd1 vccd1 vccd1 _14405__579/A sky130_fd_sc_hd__clkbuf_16
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__05012_ _17298_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05012_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14307__500 _14311__504/A vssd1 vssd1 vccd1 vccd1 _18135_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18555_ _18555_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
X_12979_ _12999_/S vssd1 vssd1 vccd1 vccd1 _12993_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15767_/A vssd1 vssd1 vccd1 vccd1 _15767_/X sky130_fd_sc_hd__buf_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14718_ _18591_/Q _18305_/Q _17571_/Q _18842_/Q _14579_/X _14641_/X vssd1 vssd1 vccd1
+ vccd1 _14718_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18486_ _18486_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17437_ _17437_/A vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _14679_/A _14649_/B vssd1 vssd1 vccd1 vccd1 _14649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17368_ _19275_/Q _12180_/X _12298_/A _19289_/Q _17367_/X vssd1 vssd1 vccd1 vccd1
+ _17368_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19107_ _19107_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19038_ _19039_/CLK _19038_/D vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput101 _11706_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__buf_2
X_15420__917 _15422__919/A vssd1 vssd1 vccd1 vccd1 _18604_/CLK sky130_fd_sc_hd__inv_2
Xoutput112 _11747_/X vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_2
X_14869__789 _14869__789/A vssd1 vssd1 vccd1 vccd1 _18434_/CLK sky130_fd_sc_hd__inv_2
Xoutput123 _11708_/X vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_2
Xoutput134 _17871_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_2
XFILLER_142_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput145 _11843_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput156 _11814_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__04589_ _16718_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04589_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_214_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09624_ _15303_/A vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__buf_2
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14167__445 _14168__446/A vssd1 vssd1 vccd1 vccd1 _18053_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _09555_/A vssd1 vssd1 vccd1 vccd1 _18954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _17776_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03400_ clkbuf_0__03400_/X vssd1 vssd1 vccd1 vccd1 _14770__709/A sky130_fd_sc_hd__clkbuf_16
X_09486_ _18886_/Q vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__buf_4
XFILLER_196_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03193_ clkbuf_0__03193_/X vssd1 vssd1 vccd1 vccd1 _14509__663/A sky130_fd_sc_hd__clkbuf_16
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ _10352_/S vssd1 vssd1 vccd1 vccd1 _10343_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ _10261_/A vssd1 vssd1 vccd1 vccd1 _18631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12000_ _19263_/Q vssd1 vssd1 vccd1 vccd1 _17279_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10192_ _18475_/Q vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13951_/A vssd1 vssd1 vccd1 vccd1 _13951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12902_ _17972_/Q _17664_/Q _12908_/S vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__mux2_1
XFILLER_143_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13882_ _17936_/Q _13878_/X _13881_/Y vssd1 vssd1 vccd1 vccd1 _17936_/D sky130_fd_sc_hd__o21a_1
X_16670_ _16670_/A vssd1 vssd1 vccd1 vccd1 _16670_/X sky130_fd_sc_hd__buf_1
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12833_ _12833_/A vssd1 vssd1 vccd1 vccd1 _17651_/D sky130_fd_sc_hd__clkbuf_1
X_15621_ _15630_/A _15622_/B vssd1 vssd1 vccd1 vccd1 _15621_/X sky130_fd_sc_hd__or2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18340_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12764_/A vssd1 vssd1 vccd1 vccd1 _12764_/Y sky130_fd_sc_hd__inv_2
X_15552_ _15557_/B _15569_/B vssd1 vssd1 vccd1 vccd1 _15552_/Y sky130_fd_sc_hd__nand2_1
X_17080__64 _17080__64/A vssd1 vssd1 vccd1 vccd1 _19213_/CLK sky130_fd_sc_hd__inv_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04578_ clkbuf_0__04578_/X vssd1 vssd1 vccd1 vccd1 _16682__314/A sky130_fd_sc_hd__clkbuf_16
XFILLER_70_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ _11715_/A vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15483_ _17830_/Q _15489_/B _17829_/Q vssd1 vssd1 vccd1 vccd1 _15484_/B sky130_fd_sc_hd__o21ai_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _18271_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
X_12695_ _12695_/A vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17222_ _17222_/A _17222_/B vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__nor2_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11646_ _11646_/A vssd1 vssd1 vccd1 vccd1 _17536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 io_in[24] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_6
XFILLER_122_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17153_ _17153_/A vssd1 vssd1 vccd1 vccd1 _19229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput25 vga_b[1] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_8
X_14302__496 _14302__496/A vssd1 vssd1 vccd1 vccd1 _18131_/CLK sky130_fd_sc_hd__inv_2
Xinput36 wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
X_11577_ _17583_/Q _10904_/X _11581_/S vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput47 wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
X_13316_ _13265_/X _13311_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _13316_/Y sky130_fd_sc_hd__a21oi_1
Xinput58 wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16104_ _16280_/A _16104_/B vssd1 vssd1 vccd1 vccd1 _16104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput69 wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_4
X_10528_ _10546_/B _10528_/B vssd1 vssd1 vccd1 vccd1 _10544_/S sky130_fd_sc_hd__nor2_2
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13247_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13247_/X sky130_fd_sc_hd__buf_4
X_16035_ _18876_/Q _16035_/B _16035_/C vssd1 vssd1 vccd1 vccd1 _16036_/D sky130_fd_sc_hd__nand3_1
X_10459_ _10459_/A vssd1 vssd1 vccd1 vccd1 _18547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _13362_/A vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12129_ _17516_/Q _17735_/Q _12136_/S vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__mux2_1
X_15673__974 _15673__974/A vssd1 vssd1 vccd1 vccd1 _18691_/CLK sky130_fd_sc_hd__inv_2
X_17986_ _19247_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 _17986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__04374_ _16340_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04374_/X sky130_fd_sc_hd__clkbuf_16
X_16937_ _18152_/Q _18144_/Q _18136_/Q _18280_/Q _16809_/X _16810_/X vssd1 vssd1 vccd1
+ vccd1 _16937_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16868_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16868_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_225_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18607_ _18607_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03156_ clkbuf_0__03156_/X vssd1 vssd1 vccd1 vccd1 _14323__514/A sky130_fd_sc_hd__clkbuf_16
X_15819_ _15813_/Y _15815_/X _15818_/X vssd1 vssd1 vccd1 vccd1 _15819_/X sky130_fd_sc_hd__a21o_1
X_16799_ _16881_/A vssd1 vssd1 vccd1 vccd1 _16799_/X sky130_fd_sc_hd__buf_4
XFILLER_241_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ _10638_/A _10157_/A vssd1 vssd1 vccd1 vccd1 _09356_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_0__03187_ _14474_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03187_/X sky130_fd_sc_hd__clkbuf_16
X_18538_ _18538_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09271_ _18476_/Q vssd1 vssd1 vccd1 vccd1 _09271_/X sky130_fd_sc_hd__clkbuf_4
X_14875__793 _14876__794/A vssd1 vssd1 vccd1 vccd1 _18438_/CLK sky130_fd_sc_hd__inv_2
X_18469_ _18482_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03989_ clkbuf_0__03989_/X vssd1 vssd1 vccd1 vccd1 _15824_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_146_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15839__141 _15840__142/A vssd1 vssd1 vccd1 vccd1 _18816_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ _19213_/Q _08964_/X _08988_/S vssd1 vssd1 vccd1 vccd1 _08987_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17295__72 _17296__73/A vssd1 vssd1 vccd1 vccd1 _19268_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09607_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__buf_2
XFILLER_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09538_ _18961_/Q _09498_/X _09542_/S vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__mux2_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09469_ hold13/A _11547_/A vssd1 vssd1 vccd1 vccd1 _10670_/S sky130_fd_sc_hd__nor2_2
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14141__426 _14141__426/A vssd1 vssd1 vccd1 vccd1 _18034_/CLK sky130_fd_sc_hd__inv_2
X_11500_ _11500_/A vssd1 vssd1 vccd1 vccd1 _18045_/D sky130_fd_sc_hd__clkbuf_1
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12480_ _12480_/A vssd1 vssd1 vccd1 vccd1 _12480_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11431_ _11431_/A vssd1 vssd1 vccd1 vccd1 _18102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11362_ _11362_/A vssd1 vssd1 vccd1 vccd1 _18132_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__03176_ clkbuf_0__03176_/X vssd1 vssd1 vccd1 vccd1 _14425_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10313_ _10313_/A vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ _14081_/A _14083_/B vssd1 vssd1 vccd1 vccd1 _14081_/Y sky130_fd_sc_hd__nor2_2
X_11293_ _18159_/Q _11270_/X _11295_/S vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _13066_/A vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10244_ _18638_/Q _10183_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17840_ _17840_/CLK _17840_/D vssd1 vssd1 vccd1 vccd1 _17840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10175_ _18480_/Q vssd1 vssd1 vccd1 vccd1 _10175_/X sky130_fd_sc_hd__buf_4
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17771_ _17772_/CLK _17771_/D vssd1 vssd1 vccd1 vccd1 _17771_/Q sky130_fd_sc_hd__dfxtp_2
X_14983_ _15001_/A _14983_/B vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__and2_1
XFILLER_247_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13934_ _17955_/Q _13941_/B vssd1 vssd1 vccd1 vccd1 _13934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_234_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13865_ input66/X _13867_/B vssd1 vssd1 vccd1 vccd1 _13865_/X sky130_fd_sc_hd__and2_1
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053__42 _17053__42/A vssd1 vssd1 vccd1 vccd1 _19191_/CLK sky130_fd_sc_hd__inv_2
X_15604_ _18655_/Q _15604_/B vssd1 vssd1 vccd1 vccd1 _15606_/B sky130_fd_sc_hd__nor2_1
X_12816_ _17647_/Q _17988_/Q _12822_/S vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__mux2_1
X_16584_ _16584_/A vssd1 vssd1 vccd1 vccd1 _16613_/A sky130_fd_sc_hd__buf_2
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13796_ _13802_/A vssd1 vssd1 vccd1 vccd1 _13796_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152__862 _15153__863/A vssd1 vssd1 vccd1 vccd1 _18538_/CLK sky130_fd_sc_hd__inv_2
XFILLER_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18323_ _19013_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15535_ _15535_/A _18669_/Q _15535_/C vssd1 vssd1 vccd1 vccd1 _15574_/A sky130_fd_sc_hd__and3_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A vssd1 vssd1 vccd1 vccd1 _12758_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18254_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
X_12678_ _17611_/Q _12673_/X _12663_/X vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__o21ai_1
X_15466_ _08998_/Y _14244_/A _13892_/A vssd1 vssd1 vccd1 vccd1 _15470_/A sky130_fd_sc_hd__a21o_4
XFILLER_176_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16632__274 _16632__274/A vssd1 vssd1 vccd1 vccd1 _19048_/CLK sky130_fd_sc_hd__inv_2
XFILLER_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17205_ _19243_/Q _17202_/A _17164_/X vssd1 vssd1 vccd1 vccd1 _17206_/B sky130_fd_sc_hd__o21ai_1
XFILLER_128_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11629_ _17543_/Q _09688_/A _11629_/S vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18185_ _18185_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17136_ _17142_/C _17136_/B _17277_/B vssd1 vssd1 vccd1 vccd1 _17137_/A sky130_fd_sc_hd__and3b_1
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16018_ _18872_/Q _16018_/B _16018_/C vssd1 vssd1 vccd1 vccd1 _16027_/C sky130_fd_sc_hd__and3_1
XFILLER_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762__702 _14763__703/A vssd1 vssd1 vccd1 vccd1 _18345_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08840_ _19049_/Q vssd1 vssd1 vccd1 vccd1 _09446_/A sky130_fd_sc_hd__inv_2
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08756_/X _08761_/B _09611_/B _08769_/B vssd1 vssd1 vccd1 vccd1 _08772_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17969_ _17969_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200__885 _15203__888/A vssd1 vssd1 vccd1 vccd1 _18564_/CLK sky130_fd_sc_hd__inv_2
X_16674__308 _16674__308/A vssd1 vssd1 vccd1 vccd1 _19082_/CLK sky130_fd_sc_hd__inv_2
XFILLER_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09323_ _09323_/A vssd1 vssd1 vccd1 vccd1 _19099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09254_ _08728_/X _09253_/X _11675_/A vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__a21oi_4
X_15716__1009 _15716__1009/A vssd1 vssd1 vccd1 vccd1 _18726_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ _09185_/A vssd1 vssd1 vccd1 vccd1 _19164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19240_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ _08969_/A vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11980_ _11980_/A vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03794_ clkbuf_0__03794_/X vssd1 vssd1 vccd1 vccd1 _15391__894/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _10931_/A _11601_/B vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__nor2_2
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13650_ _13650_/A vssd1 vssd1 vccd1 vccd1 _16532_/B sky130_fd_sc_hd__clkbuf_4
X_10862_ _10862_/A vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _18013_/Q _17591_/Q _17590_/Q _17589_/Q vssd1 vssd1 vccd1 vccd1 _12614_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ _16059_/A _13574_/B _13580_/Y _13569_/X vssd1 vssd1 vccd1 vccd1 _17838_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _10793_/A vssd1 vssd1 vccd1 vccd1 _18370_/D sky130_fd_sc_hd__clkbuf_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12532_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15320_ _18939_/Q _18902_/Q _18894_/Q _18848_/Q _15248_/X _15252_/X vssd1 vssd1 vccd1
+ vccd1 _15320_/X sky130_fd_sc_hd__mux4_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ _12389_/X _12374_/X _12464_/S vssd1 vssd1 vccd1 vccd1 _12463_/X sky130_fd_sc_hd__mux2_1
X_15251_ _15273_/A vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__buf_2
XFILLER_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _11338_/X _18109_/Q _11418_/S vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__mux2_1
X_14202_ _14202_/A vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15182_ _18660_/Q vssd1 vssd1 vccd1 vccd1 _15182_/Y sky130_fd_sc_hd__inv_2
X_12394_ _17594_/Q vssd1 vssd1 vccd1 vccd1 _12394_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14133_ _18029_/Q _14115_/X _14132_/Y vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__o21a_1
X_11345_ _11344_/X _18139_/Q _11345_/S vssd1 vssd1 vccd1 vccd1 _11346_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03159_ clkbuf_0__03159_/X vssd1 vssd1 vccd1 vccd1 _14334__522/A sky130_fd_sc_hd__clkbuf_16
X_14064_ _18003_/Q _14054_/X _14063_/Y vssd1 vssd1 vccd1 vccd1 _18003_/D sky130_fd_sc_hd__o21a_1
XFILLER_180_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18941_ _18941_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03590_ _15106_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03590_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11276_ _18663_/Q vssd1 vssd1 vccd1 vccd1 _11276_/X sky130_fd_sc_hd__buf_2
XFILLER_180_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ _17674_/Q _13094_/B vssd1 vssd1 vccd1 vccd1 _13019_/A sky130_fd_sc_hd__xnor2_1
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14414__586 _14414__586/A vssd1 vssd1 vccd1 vccd1 _18221_/CLK sky130_fd_sc_hd__inv_2
X_10227_ _10227_/A vssd1 vssd1 vccd1 vccd1 _18676_/D sky130_fd_sc_hd__clkbuf_1
X_18872_ _18879_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_1
X_14826__754 _14826__754/A vssd1 vssd1 vccd1 vccd1 _18397_/CLK sky130_fd_sc_hd__inv_2
X_17823_ _19147_/CLK _17823_/D vssd1 vssd1 vccd1 vccd1 _17823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _10173_/S vssd1 vssd1 vccd1 vccd1 _10167_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15788__110 _15788__110/A vssd1 vssd1 vccd1 vccd1 _18782_/CLK sky130_fd_sc_hd__inv_2
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17754_ _19290_/CLK _17754_/D vssd1 vssd1 vccd1 vccd1 _17754_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14966_ _18481_/Q _15074_/C vssd1 vssd1 vccd1 vccd1 _14991_/A sky130_fd_sc_hd__and2_1
X_10089_ _10089_/A vssd1 vssd1 vccd1 vccd1 _18729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13917_ _17949_/Q _13903_/X _13916_/Y vssd1 vssd1 vccd1 vccd1 _17949_/D sky130_fd_sc_hd__o21a_1
X_17026__20 _17028__22/A vssd1 vssd1 vccd1 vccd1 _19169_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17685_ _17703_/CLK _17685_/D vssd1 vssd1 vccd1 vccd1 _17685_/Q sky130_fd_sc_hd__dfxtp_1
X_14897_ _18469_/Q vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__inv_2
XFILLER_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13848_ _17927_/Q _13829_/A _13847_/X _13841_/X vssd1 vssd1 vccd1 vccd1 _17927_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16567_ _16567_/A _19017_/Q _19016_/Q vssd1 vssd1 vccd1 vccd1 _16569_/B sky130_fd_sc_hd__and3_1
XFILLER_210_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13779_ _13777_/X _13778_/X _13774_/X vssd1 vssd1 vccd1 vccd1 _13779_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16337__233 _16337__233/A vssd1 vssd1 vccd1 vccd1 _18949_/CLK sky130_fd_sc_hd__inv_2
X_18306_ _18306_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15518_ _18645_/Q vssd1 vssd1 vccd1 vccd1 _15557_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _19287_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16498_ _16498_/A _16498_/B _16498_/C vssd1 vssd1 vccd1 vccd1 _16498_/X sky130_fd_sc_hd__or3_1
XFILLER_200_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _18237_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15449_ _15455_/A vssd1 vssd1 vccd1 vccd1 _15449_/X sky130_fd_sc_hd__buf_1
XFILLER_102_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ _18168_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17119_ _17119_/A vssd1 vssd1 vccd1 vccd1 _19221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18099_ _18099_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16680__312 _16680__312/A vssd1 vssd1 vccd1 vccd1 _19086_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _09941_/A vssd1 vssd1 vccd1 vccd1 _18782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _18809_/D sky130_fd_sc_hd__nor2_1
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__clkbuf_1
X_16344__237 _16344__237/A vssd1 vssd1 vccd1 vccd1 _18953_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15198__884 _15198__884/A vssd1 vssd1 vccd1 vccd1 _18563_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_16 _11707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_27 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_38 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08754_ _08769_/B vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_49 _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09306_ _08917_/X _19106_/Q _09312_/S vssd1 vssd1 vccd1 vccd1 _09307_/A sky130_fd_sc_hd__mux2_1
X_15389__892 _15389__892/A vssd1 vssd1 vccd1 vccd1 _18579_/CLK sky130_fd_sc_hd__inv_2
XFILLER_179_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09237_ _18566_/Q _10075_/B vssd1 vssd1 vccd1 vccd1 _10403_/B sky130_fd_sc_hd__xnor2_2
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09168_ _10869_/A _10752_/A vssd1 vssd1 vccd1 vccd1 _09184_/S sky130_fd_sc_hd__nor2_2
XFILLER_182_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14769__708 _14770__709/A vssd1 vssd1 vccd1 vccd1 _18351_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09099_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322__386 _12322__386/A vssd1 vssd1 vccd1 vccd1 _17567_/CLK sky130_fd_sc_hd__inv_2
XFILLER_218_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11130_ _18224_/Q _11050_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11061_ _11061_/A vssd1 vssd1 vccd1 vccd1 _18253_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10012_ _10094_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10028_/S sky130_fd_sc_hd__nor2_2
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11963_ _19255_/Q vssd1 vssd1 vccd1 vccd1 _17250_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13274_/X _13688_/A _13701_/X vssd1 vssd1 vccd1 vccd1 _13702_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_233_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17470_ _17470_/A vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__clkbuf_1
X_10914_ _10929_/S vssd1 vssd1 vccd1 vccd1 _10923_/S sky130_fd_sc_hd__clkbuf_2
X_11894_ _11975_/S vssd1 vssd1 vccd1 vccd1 _11924_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_232_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14607_/X _14675_/Y _14677_/Y _14679_/Y _14681_/Y vssd1 vssd1 vccd1 vccd1
+ _14682_/X sky130_fd_sc_hd__o32a_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _16421_/A _16421_/B _16421_/C _16421_/D vssd1 vssd1 vccd1 vccd1 _16421_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_232_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13633_ _17856_/Q _13635_/B vssd1 vssd1 vccd1 vccd1 _13633_/Y sky130_fd_sc_hd__nor2_1
X_10845_ _18349_/Q _10806_/X _10849_/S vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19140_ _19144_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13564_ _17833_/Q _13568_/B vssd1 vssd1 vccd1 vccd1 _13564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10776_ _10776_/A vssd1 vssd1 vccd1 vccd1 _18377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ _15303_/A vssd1 vssd1 vccd1 vccd1 _15303_/X sky130_fd_sc_hd__clkbuf_1
X_12515_ _12515_/A _12515_/B vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__or2_1
X_19071_ _19071_/CLK _19071_/D vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfxtp_1
X_14420__590 _14424__594/A vssd1 vssd1 vccd1 vccd1 _18225_/CLK sky130_fd_sc_hd__inv_2
X_13495_ _13712_/A _13490_/Y _13494_/X vssd1 vssd1 vccd1 vccd1 _13495_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16283_ _16191_/X _16276_/Y _16278_/Y _16280_/Y _16282_/Y vssd1 vssd1 vccd1 vccd1
+ _16283_/X sky130_fd_sc_hd__o32a_2
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18022_ _18029_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ _17593_/Q _12394_/X _17595_/Q _12622_/A _12443_/X _12556_/A vssd1 vssd1 vccd1
+ vccd1 _12446_/X sky130_fd_sc_hd__mux4_1
X_15234_ _19067_/Q _19059_/Q _19051_/Q _19005_/Q _15232_/X _15233_/X vssd1 vssd1 vccd1
+ vccd1 _15235_/A sky130_fd_sc_hd__mux4_1
XFILLER_154_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12377_ _17612_/Q _17613_/Q _12443_/A vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04591_ clkbuf_0__04591_/X vssd1 vssd1 vccd1 vccd1 _16730__344/A sky130_fd_sc_hd__clkbuf_16
XFILLER_236_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14116_ _13740_/A _14115_/X _14108_/X vssd1 vssd1 vccd1 vccd1 _14116_/Y sky130_fd_sc_hd__a21oi_1
X_11328_ _11328_/A vssd1 vssd1 vccd1 vccd1 _18145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18924_ _18924_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_1
X_14047_ _13414_/A _14039_/X _14046_/X vssd1 vssd1 vccd1 vccd1 _14047_/Y sky130_fd_sc_hd__a21oi_1
X_11259_ _18668_/Q vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18855_ _18855_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_1
X_15715__1008 _15716__1009/A vssd1 vssd1 vccd1 vccd1 _18725_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17806_ _19133_/CLK _17806_/D vssd1 vssd1 vccd1 vccd1 _17806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ _18786_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15998_ _16025_/B vssd1 vssd1 vccd1 vccd1 _16020_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_243_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17737_ _17737_/CLK _17737_/D vssd1 vssd1 vccd1 vccd1 _17737_/Q sky130_fd_sc_hd__dfxtp_1
X_14949_ _18456_/Q _14949_/B vssd1 vssd1 vccd1 vccd1 _14950_/D sky130_fd_sc_hd__xor2_1
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17668_ _19027_/CLK _17668_/D vssd1 vssd1 vccd1 vccd1 _17668_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_120 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_131 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_142 _11811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16619_ _16619_/A _16619_/B _16619_/C vssd1 vssd1 vccd1 vccd1 _19038_/D sky130_fd_sc_hd__nor3_1
XINSDIODE2_153 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_164 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ _17602_/CLK _17599_/D vssd1 vssd1 vccd1 vccd1 _17599_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_175 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_186 _16228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19338_ _19339_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_197 _10797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19269_ _19269_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
X_09022_ _11222_/A vssd1 vssd1 vccd1 vccd1 _09025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03809_ clkbuf_0__03809_/X vssd1 vssd1 vccd1 vccd1 _15464__952/A sky130_fd_sc_hd__clkbuf_16
X_15165__872 _15165__872/A vssd1 vssd1 vccd1 vccd1 _18548_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16088__201 _16090__203/A vssd1 vssd1 vccd1 vccd1 _18906_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09924_ _18787_/Q _09268_/X _09926_/S vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _16868_/A vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__buf_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ _08806_/A vssd1 vssd1 vccd1 vccd1 _19341_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09786_ _09786_/A vssd1 vssd1 vccd1 vccd1 _18837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _18077_/Q vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _18440_/Q _10126_/A _10630_/S vssd1 vssd1 vccd1 vccd1 _10631_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17020__15 _17022__17/A vssd1 vssd1 vccd1 vccd1 _19164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10561_ _10561_/A vssd1 vssd1 vccd1 vccd1 _18501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12300_ _17562_/Q _12298_/X _12182_/X _17551_/Q _12299_/Y vssd1 vssd1 vccd1 vccd1
+ _12301_/C sky130_fd_sc_hd__o221a_1
XFILLER_167_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13280_ _13288_/A vssd1 vssd1 vccd1 vccd1 _13280_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10492_ _10602_/B _10492_/B vssd1 vssd1 vccd1 vccd1 _10508_/S sky130_fd_sc_hd__or2_2
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14257__460 _14261__464/A vssd1 vssd1 vccd1 vccd1 _18095_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12162_ _12162_/A vssd1 vssd1 vccd1 vccd1 _17525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11113_ _11113_/A vssd1 vssd1 vccd1 vccd1 _18232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _12034_/A _12075_/B _12092_/X _12020_/A vssd1 vssd1 vccd1 vccd1 _12093_/X
+ sky130_fd_sc_hd__a211o_1
X_16970_ _16836_/X _16963_/Y _16965_/Y _16967_/Y _16969_/Y vssd1 vssd1 vccd1 vccd1
+ _16970_/X sky130_fd_sc_hd__o32a_1
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15439__933 _15439__933/A vssd1 vssd1 vccd1 vccd1 _18620_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _11066_/S vssd1 vssd1 vccd1 vccd1 _11057_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15921_ _18863_/Q vssd1 vssd1 vccd1 vccd1 _15970_/A sky130_fd_sc_hd__inv_2
XFILLER_237_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _18640_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18571_ _18572_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12995_ _12995_/A vssd1 vssd1 vccd1 vccd1 _17683_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14526__676 _14527__677/A vssd1 vssd1 vccd1 vccd1 _18311_/CLK sky130_fd_sc_hd__inv_2
XFILLER_229_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17522_ _17737_/CLK _17522_/D vssd1 vssd1 vccd1 vccd1 _17522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14734_/A _14734_/B vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11946_ _11907_/X _11918_/X _11927_/X _11939_/X _12016_/S _11945_/X vssd1 vssd1 vccd1
+ vccd1 _11947_/A sky130_fd_sc_hd__mux4_2
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _17453_/A vssd1 vssd1 vccd1 vccd1 _19332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14665_ _09433_/X _14656_/X _14664_/Y _14543_/A vssd1 vssd1 vccd1 vccd1 _14665_/Y
+ sky130_fd_sc_hd__o211ai_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16404_ _18971_/Q _16404_/B vssd1 vssd1 vccd1 vccd1 _16411_/A sky130_fd_sc_hd__xor2_1
X_13616_ _17850_/Q _13621_/B vssd1 vssd1 vccd1 vccd1 _13616_/Y sky130_fd_sc_hd__nor2_1
X_10828_ _10828_/A vssd1 vssd1 vccd1 vccd1 _18357_/D sky130_fd_sc_hd__clkbuf_1
X_17384_ _17384_/A vssd1 vssd1 vccd1 vccd1 _17384_/X sky130_fd_sc_hd__buf_1
X_14596_ _18404_/Q _18396_/Q _19309_/Q _17713_/Q _14594_/X _14595_/X vssd1 vssd1 vccd1
+ vccd1 _14596_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19123_ _19123_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_13547_ _13599_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _13559_/S sky130_fd_sc_hd__nor2_4
X_10759_ _10759_/A vssd1 vssd1 vccd1 vccd1 _18384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19054_ _19054_/CLK _19054_/D vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfxtp_1
X_16266_ _18717_/Q _18725_/Q _18733_/Q _18498_/Q _16205_/X _16206_/X vssd1 vssd1 vccd1
+ vccd1 _16266_/X sky130_fd_sc_hd__mux4_2
XFILLER_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13478_ _16057_/A _13463_/B _13477_/Y _13472_/X vssd1 vssd1 vccd1 vccd1 _17806_/D
+ sky130_fd_sc_hd__a211oi_1
X_18005_ _18014_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
X_15217_ _18997_/Q _18959_/Q _18951_/Q _17540_/Q _15214_/X _15215_/X vssd1 vssd1 vccd1
+ vccd1 _15217_/X sky130_fd_sc_hd__mux4_1
X_12429_ _12426_/X _12428_/X _12429_/S vssd1 vssd1 vccd1 vccd1 _12429_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16197_ _16278_/A _16197_/B vssd1 vssd1 vccd1 vccd1 _16197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__04574_ clkbuf_0__04574_/X vssd1 vssd1 vccd1 vccd1 _16659__295/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_9_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15833__136 _15833__136/A vssd1 vssd1 vccd1 vccd1 _18811_/CLK sky130_fd_sc_hd__inv_2
X_15079_ _18482_/Q _15079_/B vssd1 vssd1 vccd1 vccd1 _15079_/Y sky130_fd_sc_hd__nor2_1
X_18907_ _18907_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09640_ _09636_/Y _09640_/B _09649_/C vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__and3b_1
X_18838_ _18838_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09571_ _09571_/A vssd1 vssd1 vccd1 vccd1 _18947_/D sky130_fd_sc_hd__clkbuf_1
X_18769_ _18769_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16083__197 _16085__199/A vssd1 vssd1 vccd1 vccd1 _18902_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14427__596 _14427__596/A vssd1 vssd1 vccd1 vccd1 _18231_/CLK sky130_fd_sc_hd__inv_2
XFILLER_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04008_ clkbuf_0__04008_/X vssd1 vssd1 vccd1 vccd1 _15848__149/A sky130_fd_sc_hd__clkbuf_16
XFILLER_212_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _09001_/Y _11068_/B _09011_/A _09004_/Y vssd1 vssd1 vccd1 vccd1 _09005_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09907_ _18794_/Q _09732_/X _09907_/S vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09838_ _09691_/X _18814_/Q _09842_/S vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09769_ _09769_/A vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _16689_/A vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784__1064 _15784__1064/A vssd1 vssd1 vccd1 vccd1 _18781_/CLK sky130_fd_sc_hd__inv_2
X_12780_ _12761_/X _12780_/B vssd1 vssd1 vccd1 vccd1 _12781_/A sky130_fd_sc_hd__and2b_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11731_ _17913_/Q _17787_/Q _11869_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__mux2_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14456_/A vssd1 vssd1 vccd1 vccd1 _14450_/X sky130_fd_sc_hd__buf_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _11662_/A vssd1 vssd1 vccd1 vccd1 _17512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13401_ _17785_/Q _13405_/B _13400_/Y _13376_/X vssd1 vssd1 vccd1 vccd1 _17785_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ _10613_/A vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11593_ _17576_/Q _10704_/A _11593_/S vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__mux2_1
X_15714__1007 _15714__1007/A vssd1 vssd1 vccd1 vccd1 _18724_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _10406_/B _16118_/X _16119_/X vssd1 vssd1 vccd1 vccd1 _16120_/Y sky130_fd_sc_hd__o21ai_1
XPeripherals_169 vssd1 vssd1 vccd1 vccd1 Peripherals_169/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XFILLER_183_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13332_ _17769_/Q _13329_/X _13331_/Y vssd1 vssd1 vccd1 vccd1 _17769_/D sky130_fd_sc_hd__o21a_1
X_10544_ _18508_/Q _10351_/X _10544_/S vssd1 vssd1 vccd1 vccd1 _10545_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16051_ _18879_/Q _16050_/A _16050_/Y _15242_/X vssd1 vssd1 vccd1 vccd1 _18879_/D
+ sky130_fd_sc_hd__o211a_1
X_13263_ _13192_/X _13259_/X _13260_/X vssd1 vssd1 vccd1 vccd1 _13263_/Y sky130_fd_sc_hd__a21oi_1
X_10475_ _10490_/S vssd1 vssd1 vccd1 vccd1 _10484_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_124_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__05077_ clkbuf_0__05077_/X vssd1 vssd1 vccd1 vccd1 _17415_/A sky130_fd_sc_hd__clkbuf_16
X_15002_ _15002_/A vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _12214_/A vssd1 vssd1 vccd1 vccd1 _17478_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13194_ _13170_/X _13192_/X _13193_/Y _13187_/X vssd1 vssd1 vccd1 vccd1 _17732_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12145_ _12145_/A vssd1 vssd1 vccd1 vccd1 _17520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03410_ _14815_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03410_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12076_ _11957_/X _11962_/X _12076_/S vssd1 vssd1 vccd1 vccd1 _12076_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16953_ _16892_/X _16942_/X _16952_/Y vssd1 vssd1 vccd1 vccd1 _16953_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11027_ _11027_/A vssd1 vssd1 vccd1 vccd1 _18266_/D sky130_fd_sc_hd__clkbuf_1
X_15904_ _17812_/Q _15947_/A vssd1 vssd1 vccd1 vccd1 _15951_/A sky130_fd_sc_hd__or2_1
XFILLER_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16884_ _16929_/A _16884_/B vssd1 vssd1 vccd1 vccd1 _16884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12335__396 _12335__396/A vssd1 vssd1 vccd1 vccd1 _17577_/CLK sky130_fd_sc_hd__inv_2
X_18623_ _18623_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03172_ clkbuf_0__03172_/X vssd1 vssd1 vccd1 vccd1 _14396__571/A sky130_fd_sc_hd__clkbuf_16
XFILLER_237_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18554_ _18554_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _12978_/A vssd1 vssd1 vccd1 vccd1 _17678_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15116__833 _15117__834/A vssd1 vssd1 vccd1 vccd1 _18509_/CLK sky130_fd_sc_hd__inv_2
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14717_ _14736_/A _14717_/B vssd1 vssd1 vccd1 vccd1 _14717_/Y sky130_fd_sc_hd__nor2_1
X_11929_ _17781_/Q vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__buf_2
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18485_ _18485_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17436_ _17436_/A vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14648_ _19151_/Q _18416_/Q _18310_/Q _18294_/Q _14580_/X _09444_/A vssd1 vssd1 vccd1
+ vccd1 _14649_/B sky130_fd_sc_hd__mux4_1
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17367_ _19276_/Q _12187_/A _12199_/A _19286_/Q vssd1 vssd1 vccd1 vccd1 _17367_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_242_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14579_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14579_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19106_ _19106_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17298_ _17384_/A vssd1 vssd1 vccd1 vccd1 _17298_/X sky130_fd_sc_hd__buf_1
X_19037_ _19037_/CLK _19037_/D vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfxtp_1
X_16249_ _18630_/Q _18505_/Q _18911_/Q _18513_/Q _16155_/X _16156_/X vssd1 vssd1 vccd1
+ vccd1 _16249_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput102 _11702_/X vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput113 _11743_/X vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_2
Xoutput124 _11704_/X vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_2
XFILLER_173_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput135 _19386_/X vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_2
Xoutput146 _11846_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[12] sky130_fd_sc_hd__buf_2
XFILLER_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput157 _11818_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _09623_/A vssd1 vssd1 vccd1 vccd1 _18933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09554_ _08929_/X _18954_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09485_ _09485_/A vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_77_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17602_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_168_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03192_ clkbuf_0__03192_/X vssd1 vssd1 vccd1 vccd1 _14504__659/A sky130_fd_sc_hd__clkbuf_16
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _18631_/Q _10180_/X _10266_/S vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10191_ _10191_/A vssd1 vssd1 vccd1 vccd1 _18690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _17961_/Q _13950_/B vssd1 vssd1 vccd1 vccd1 _13950_/Y sky130_fd_sc_hd__nor2_1
X_14369__550 _14370__551/A vssd1 vssd1 vccd1 vccd1 _18185_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12901_ _12901_/A vssd1 vssd1 vccd1 vccd1 _17663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13881_ _13281_/X _13879_/X _13880_/X vssd1 vssd1 vccd1 vccd1 _13881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14820__749 _14820__749/A vssd1 vssd1 vccd1 vccd1 _18392_/CLK sky130_fd_sc_hd__inv_2
XFILLER_207_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15620_ _15618_/Y _15642_/B _15619_/X vssd1 vssd1 vccd1 vccd1 _15622_/B sky130_fd_sc_hd__o21bai_1
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _12830_/X _12832_/B vssd1 vssd1 vccd1 vccd1 _12833_/A sky130_fd_sc_hd__and2b_1
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15551_ _15551_/A _15551_/B _15562_/C vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__or3_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12763_/A vssd1 vssd1 vccd1 vccd1 _13081_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04577_ clkbuf_0__04577_/X vssd1 vssd1 vccd1 vccd1 _16707_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _17909_/Q _11714_/B vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__and2_4
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _18270_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15482_ _18656_/Q _15482_/B vssd1 vssd1 vccd1 vccd1 _15482_/X sky130_fd_sc_hd__or2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _17616_/Q _17615_/Q _12694_/C _12694_/D vssd1 vssd1 vccd1 vccd1 _12707_/C
+ sky130_fd_sc_hd__and4_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17225_/C _17225_/D _17126_/X vssd1 vssd1 vccd1 vccd1 _17222_/B sky130_fd_sc_hd__o21ai_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11645_ _08792_/X _17536_/Q _11647_/S vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17152_ _17162_/D _17189_/B _17152_/C vssd1 vssd1 vccd1 vccd1 _17153_/A sky130_fd_sc_hd__and3b_1
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput15 io_in[25] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_6
XFILLER_156_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 vga_g[0] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_16
X_11576_ _11576_/A vssd1 vssd1 vccd1 vccd1 _17584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput48 wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
X_16331__228 _16332__229/A vssd1 vssd1 vccd1 vccd1 _18944_/CLK sky130_fd_sc_hd__inv_2
X_16103_ _18524_/Q _18532_/Q _18540_/Q _18548_/Q _10404_/A _16102_/X vssd1 vssd1 vccd1
+ vccd1 _16104_/B sky130_fd_sc_hd__mux4_1
X_13315_ _17764_/Q _13303_/X _13314_/Y vssd1 vssd1 vccd1 vccd1 _17764_/D sky130_fd_sc_hd__o21a_1
Xinput59 wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_2
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10527_ _10527_/A vssd1 vssd1 vccd1 vccd1 _18516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16034_ _16035_/B _16035_/C _18876_/Q vssd1 vssd1 vccd1 vccd1 _16036_/C sky130_fd_sc_hd__a21o_1
X_13246_ _17743_/Q _13219_/X _13245_/Y vssd1 vssd1 vccd1 vccd1 _17743_/D sky130_fd_sc_hd__o21a_1
X_10458_ _18547_/Q _10328_/X _10466_/S vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ input70/X _13446_/B vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__nand2_1
X_10389_ _10389_/A vssd1 vssd1 vccd1 vccd1 _18577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ _12128_/A vssd1 vssd1 vccd1 vccd1 _17515_/D sky130_fd_sc_hd__clkbuf_1
X_17985_ _19247_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 _17985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12059_ _17117_/B _19222_/Q _19223_/Q _17129_/A _11980_/A _12005_/S vssd1 vssd1 vccd1
+ vccd1 _12060_/B sky130_fd_sc_hd__mux4_1
X_16936_ _18120_/Q _18112_/Q _18104_/Q _18096_/Q _16893_/X _16894_/X vssd1 vssd1 vccd1
+ vccd1 _16936_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_0__04373_ _16339_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04373_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16867_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16882_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18606_ _18606_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_1
X_15818_ _18879_/Q _15816_/X _16049_/A _16063_/A vssd1 vssd1 vccd1 vccd1 _15818_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__03155_ clkbuf_0__03155_/X vssd1 vssd1 vccd1 vccd1 _14314__506/A sky130_fd_sc_hd__clkbuf_16
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16798_ _18807_/Q vssd1 vssd1 vccd1 vccd1 _16881_/A sky130_fd_sc_hd__buf_2
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03186_ _14468_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03186_/X sky130_fd_sc_hd__clkbuf_16
X_18537_ _18537_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09270_ _09270_/A vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _18482_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18399_ _18399_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03988_ clkbuf_0__03988_/X vssd1 vssd1 vccd1 vccd1 _15861_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_147_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15783__1063 _15784__1064/A vssd1 vssd1 vccd1 vccd1 _18780_/CLK sky130_fd_sc_hd__inv_2
X_14173__450 _14173__450/A vssd1 vssd1 vccd1 vccd1 _18058_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _08985_/A vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15713__1006 _15714__1007/A vssd1 vssd1 vccd1 vccd1 _18723_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09606_ _15291_/A vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09537_ _09537_/A vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _11529_/B vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09399_ _09399_/A vssd1 vssd1 vccd1 vccd1 _19066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _18102_/Q _11273_/X _11430_/S vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _18132_/Q _11279_/X _11363_/S vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03175_ clkbuf_0__03175_/X vssd1 vssd1 vccd1 vccd1 _14414__586/A sky130_fd_sc_hd__clkbuf_16
X_13100_ _13100_/A vssd1 vssd1 vccd1 vccd1 _17703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ _09674_/X _18608_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14080_ _12504_/A _14070_/X _14079_/Y _13868_/X vssd1 vssd1 vccd1 vccd1 _18009_/D
+ sky130_fd_sc_hd__a211o_1
X_11292_ _11292_/A vssd1 vssd1 vccd1 vccd1 _18160_/D sky130_fd_sc_hd__clkbuf_1
X_13031_ _13031_/A vssd1 vssd1 vccd1 vccd1 _17688_/D sky130_fd_sc_hd__clkbuf_1
X_10243_ _10243_/A vssd1 vssd1 vccd1 vccd1 _18639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10174_ _10174_/A vssd1 vssd1 vccd1 vccd1 _18695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17770_ _17772_/CLK _17770_/D vssd1 vssd1 vccd1 vccd1 _17770_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_232_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14982_ _18456_/Q _14978_/X _14981_/Y _15057_/A vssd1 vssd1 vccd1 vccd1 _14983_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13933_ _13140_/X _13925_/X _13932_/Y _13636_/X vssd1 vssd1 vccd1 vccd1 _17954_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16652_ _16658_/A vssd1 vssd1 vccd1 vccd1 _16652_/X sky130_fd_sc_hd__buf_1
X_13864_ _17932_/Q _13850_/X _13863_/Y _13857_/X vssd1 vssd1 vccd1 vccd1 _17932_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15603_ _15601_/X _15602_/Y _15581_/X vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__a21oi_1
XFILLER_62_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ _12815_/A vssd1 vssd1 vccd1 vccd1 _17646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16583_ _19022_/Q _16585_/C _16582_/Y vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__o21a_1
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ _14069_/A _13795_/B vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18322_ _18322_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15534_ _15583_/A vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12746_ _12746_/A _12746_/B _12746_/C _12746_/D vssd1 vssd1 vccd1 vccd1 _12747_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_163_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _18253_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12677_ _17611_/Q _12680_/C _12680_/D vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__and3_1
X_17204_ _17216_/C vssd1 vssd1 vccd1 vccd1 _17210_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11628_ _11628_/A vssd1 vssd1 vccd1 vccd1 _17544_/D sky130_fd_sc_hd__clkbuf_1
X_18184_ _18184_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17135_ _19225_/Q _17135_/B vssd1 vssd1 vccd1 vccd1 _17136_/B sky130_fd_sc_hd__or2_1
XFILLER_155_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11559_ _17706_/Q _10904_/X _11563_/S vssd1 vssd1 vccd1 vccd1 _11560_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16017_ _16018_/B _16018_/C _18872_/Q vssd1 vssd1 vccd1 vccd1 _16019_/B sky130_fd_sc_hd__a21oi_1
X_13229_ _13219_/X _13719_/A _13224_/X vssd1 vssd1 vccd1 vccd1 _13229_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14350__535 _14352__537/A vssd1 vssd1 vccd1 vccd1 _18170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08770_ hold14/A _08769_/B _09611_/A vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__a21oi_1
X_17968_ _19016_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16919_ _16917_/X _16918_/X _16976_/S vssd1 vssd1 vccd1 vccd1 _16919_/X sky130_fd_sc_hd__mux2_1
X_17899_ _17923_/CLK _17899_/D vssd1 vssd1 vccd1 vccd1 _17899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09322_ _19099_/Q _08944_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03169_ _14386_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03169_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_209_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09253_ _09253_/A _15064_/A vssd1 vssd1 vccd1 vccd1 _09253_/X sky130_fd_sc_hd__and2_2
XFILLER_194_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09184_ _19164_/Q _09116_/X _09184_/S vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15129__843 _15130__844/A vssd1 vssd1 vccd1 vccd1 _18519_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08968_ _19267_/Q _08967_/X _08968_/S vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15433__928 _15433__928/A vssd1 vssd1 vccd1 vccd1 _18615_/CLK sky130_fd_sc_hd__inv_2
XFILLER_216_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08899_ _19304_/Q _08792_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03793_ clkbuf_0__03793_/X vssd1 vssd1 vccd1 vccd1 _15410_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10930_ _10930_/A vssd1 vssd1 vccd1 vccd1 _18307_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_92_wb_clk_i clkbuf_opt_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19144_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _18029_/CLK sky130_fd_sc_hd__clkbuf_16
X_10861_ _18342_/Q _10803_/X _10861_/S vssd1 vssd1 vccd1 vccd1 _10862_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ _12600_/A vssd1 vssd1 vccd1 vccd1 _17590_/D sky130_fd_sc_hd__clkbuf_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _17838_/Q _13584_/B vssd1 vssd1 vccd1 vccd1 _13580_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _18370_/Q _10789_/X _10804_/S vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12500_/X _12530_/X _12765_/S vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _19317_/Q _19301_/Q _19293_/Q _19268_/Q _15248_/X _15249_/X vssd1 vssd1 vccd1
+ vccd1 _15250_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _12453_/X _12457_/X _12458_/X _12459_/X _12567_/S _12408_/A vssd1 vssd1 vccd1
+ vccd1 _12462_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14201_ _18072_/Q input52/X _14207_/S vssd1 vssd1 vccd1 vccd1 _14202_/A sky130_fd_sc_hd__mux2_1
X_11413_ _11413_/A vssd1 vssd1 vccd1 vccd1 _18110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15181_ _08998_/Y _14244_/X _13428_/A vssd1 vssd1 vccd1 vccd1 _16915_/A sky130_fd_sc_hd__a21oi_4
X_12393_ _17593_/Q vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _13815_/A _14120_/A _14123_/X vssd1 vssd1 vccd1 vccd1 _14132_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11344_ _11344_/A vssd1 vssd1 vccd1 vccd1 _11344_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__03158_ clkbuf_0__03158_/X vssd1 vssd1 vccd1 vccd1 _14329__518/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _13786_/X _14055_/X _14060_/X vssd1 vssd1 vccd1 vccd1 _14063_/Y sky130_fd_sc_hd__a21oi_1
X_18940_ _18940_/CLK _18940_/D vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11275_/A vssd1 vssd1 vccd1 vccd1 _18166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03089_ clkbuf_0__03089_/X vssd1 vssd1 vccd1 vccd1 _14144__429/A sky130_fd_sc_hd__clkbuf_16
X_13014_ _17673_/Q _12932_/A _12850_/A _17670_/Q vssd1 vssd1 vccd1 vccd1 _13020_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10226_ _18676_/Q _09752_/X _10230_/S vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18871_ _18879_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17822_ _19147_/CLK _17822_/D vssd1 vssd1 vccd1 vccd1 _17822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _10157_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10173_/S sky130_fd_sc_hd__nor2_2
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17753_ _19290_/CLK _17753_/D vssd1 vssd1 vccd1 vccd1 _17753_/Q sky130_fd_sc_hd__dfxtp_1
X_14965_ _14965_/A _14965_/B vssd1 vssd1 vccd1 vccd1 _15074_/C sky130_fd_sc_hd__nor2_1
X_10088_ _18729_/Q _10066_/X _10092_/S vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__mux2_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13916_ _13268_/X _13908_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13916_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17684_ _17963_/CLK _17684_/D vssd1 vssd1 vccd1 vccd1 _17684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14896_ _15080_/B vssd1 vssd1 vccd1 vccd1 _15001_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13847_ input72/X _13847_/B vssd1 vssd1 vccd1 vccd1 _13847_/X sky130_fd_sc_hd__and2_1
XFILLER_235_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15782__1062 _15782__1062/A vssd1 vssd1 vccd1 vccd1 _18779_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16566_ _16567_/A _19016_/Q _16565_/Y vssd1 vssd1 vccd1 vccd1 _19016_/D sky130_fd_sc_hd__o21a_1
X_13778_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13778_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_245_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15517_ _18645_/Q _15517_/B _15517_/C vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__and3_1
X_18305_ _18305_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _12737_/D _12729_/B vssd1 vssd1 vccd1 vccd1 _17626_/D sky130_fd_sc_hd__nor2_1
X_19285_ _19287_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16497_ _18982_/Q _16497_/B vssd1 vssd1 vccd1 vccd1 _16498_/C sky130_fd_sc_hd__and2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _18236_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15448_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15448_/X sky130_fd_sc_hd__buf_1
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15712__1005 _15714__1007/A vssd1 vssd1 vccd1 vccd1 _18722_/CLK sky130_fd_sc_hd__inv_2
X_18167_ _18167_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15379_ _15379_/A vssd1 vssd1 vccd1 vccd1 _15379_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _17289_/A _17118_/B _17118_/C vssd1 vssd1 vccd1 vccd1 _17119_/A sky130_fd_sc_hd__and3_1
XFILLER_128_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18098_ _18098_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09940_ _18782_/Q _09935_/X _09956_/S vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _09868_/X _09874_/A _09870_/X vssd1 vssd1 vccd1 vccd1 _09872_/B sky130_fd_sc_hd__o21ai_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _19319_/Q _08795_/X _08822_/S vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_17 _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_28 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_39 _11775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08753_ _18925_/Q vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_227_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15882__176 _15882__176/A vssd1 vssd1 vccd1 vccd1 _18851_/CLK sky130_fd_sc_hd__inv_2
XFILLER_242_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09305_ _09305_/A vssd1 vssd1 vccd1 vccd1 _19107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09236_ _09244_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__nor2_2
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09167_ _09167_/A vssd1 vssd1 vccd1 vccd1 _19172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09098_ _09098_/A vssd1 vssd1 vccd1 vccd1 _19193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _18253_/Q _11059_/X _11066_/S vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _10011_/A vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16696__320 _16697__321/A vssd1 vssd1 vccd1 vccd1 _19095_/CLK sky130_fd_sc_hd__inv_2
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _19251_/Q _17237_/B _19253_/Q _19254_/Q _11961_/X _11957_/S vssd1 vssd1 vccd1
+ vccd1 _11962_/X sky130_fd_sc_hd__mux4_2
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13880_/A vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _10931_/A hold8/X vssd1 vssd1 vccd1 vccd1 _10929_/S sky130_fd_sc_hd__nor2_2
XFILLER_217_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14640_/X _14680_/X _14561_/X vssd1 vssd1 vccd1 vccd1 _14681_/Y sky130_fd_sc_hd__o21ai_1
X_11893_ _19248_/Q vssd1 vssd1 vccd1 vccd1 _17225_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_204_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16420_ _16420_/A _16420_/B _16420_/C vssd1 vssd1 vccd1 vccd1 _16421_/D sky130_fd_sc_hd__or3_1
X_13632_ _13184_/X _13626_/B _13631_/Y _13619_/X vssd1 vssd1 vccd1 vccd1 _17855_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10844_ _10844_/A vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13563_ _13150_/X _13549_/X _13562_/Y _13555_/X vssd1 vssd1 vccd1 vccd1 _17832_/D
+ sky130_fd_sc_hd__a211oi_1
X_10775_ _18377_/Q _10695_/X _10781_/S vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15302_ _18674_/Q _18580_/Q _17535_/Q _17510_/Q _15262_/X _15301_/X vssd1 vssd1 vccd1
+ vccd1 _15304_/A sky130_fd_sc_hd__mux4_1
X_15110__828 _15111__829/A vssd1 vssd1 vccd1 vccd1 _18504_/CLK sky130_fd_sc_hd__inv_2
X_12514_ _12486_/X _12487_/X _12489_/X _12513_/X _12536_/A _12538_/A vssd1 vssd1 vccd1
+ vccd1 _12515_/B sky130_fd_sc_hd__mux4_1
XFILLER_201_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19070_ _19070_/CLK _19070_/D vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16282_ _16171_/A _16281_/X _16162_/S vssd1 vssd1 vccd1 vccd1 _16282_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13494_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13494_/X sky130_fd_sc_hd__buf_2
X_18021_ _18021_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15233_ _15308_/A vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__clkbuf_2
X_12445_ _12464_/S vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__buf_2
XFILLER_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12376_ _12374_/X _12375_/X _12390_/S vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04590_ clkbuf_0__04590_/X vssd1 vssd1 vccd1 vccd1 _16723__338/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14115_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11327_ _11326_/X _18145_/Q _11336_/S vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14154__437 _14155__438/A vssd1 vssd1 vccd1 vccd1 _18045_/CLK sky130_fd_sc_hd__inv_2
X_14046_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18923_ _19146_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_1
X_11258_ _11258_/A vssd1 vssd1 vccd1 vccd1 _18171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10209_ _18683_/Q _09755_/X _10211_/S vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__mux2_1
X_18854_ _18854_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ _11189_/A vssd1 vssd1 vccd1 vccd1 _18202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17805_ _19133_/CLK _17805_/D vssd1 vssd1 vccd1 vccd1 _17805_/Q sky130_fd_sc_hd__dfxtp_1
X_15997_ _16002_/B _16002_/C _15996_/Y vssd1 vssd1 vccd1 vccd1 _15997_/Y sky130_fd_sc_hd__o21ai_1
X_18785_ _18785_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14948_ _14948_/A _14948_/B vssd1 vssd1 vccd1 vccd1 _14949_/B sky130_fd_sc_hd__nand2_1
X_17736_ _19147_/CLK _17736_/D vssd1 vssd1 vccd1 vccd1 _17736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17667_ _19016_/CLK _17667_/D vssd1 vssd1 vccd1 vccd1 _17667_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_110 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_121 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_132 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16618_ _19037_/Q _16614_/B _19038_/Q vssd1 vssd1 vccd1 vccd1 _16619_/C sky130_fd_sc_hd__a21oi_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_143 _11814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17598_ _17602_/CLK _17598_/D vssd1 vssd1 vccd1 vccd1 _17598_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_154 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_165 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17404__95 _17405__96/A vssd1 vssd1 vccd1 vccd1 _19308_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_176 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19337_ _19337_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
X_16549_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16549_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_187 _08877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_198 _11843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19268_ _19268_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09021_ hold17/X vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18219_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19199_ _19199_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
X_16350__242 _16352__244/A vssd1 vssd1 vccd1 vccd1 _18958_/CLK sky130_fd_sc_hd__inv_2
XFILLER_145_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03808_ clkbuf_0__03808_/X vssd1 vssd1 vccd1 vccd1 _15460__949/A sky130_fd_sc_hd__clkbuf_16
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09923_ _09923_/A vssd1 vssd1 vccd1 vccd1 _18788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _16893_/A vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _19341_/Q _08804_/X _08805_/S vssd1 vssd1 vccd1 vccd1 _08806_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _08883_/X _18837_/Q _09787_/S vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _18076_/Q vssd1 vssd1 vccd1 vccd1 _13488_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_39_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14363__545 _14364__546/A vssd1 vssd1 vccd1 vccd1 _18180_/CLK sky130_fd_sc_hd__inv_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14775__713 _14776__714/A vssd1 vssd1 vccd1 vccd1 _18356_/CLK sky130_fd_sc_hd__inv_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _18501_/Q _10132_/A _10562_/S vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _19149_/Q _09112_/X _09221_/S vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _10491_/A vssd1 vssd1 vccd1 vccd1 _18532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15701__996 _15701__996/A vssd1 vssd1 vccd1 vccd1 _18713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _12149_/X _12161_/B vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__and2b_1
XFILLER_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _18232_/Q _11050_/X _11116_/S vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__mux2_1
X_15781__1061 _15782__1062/A vssd1 vssd1 vccd1 vccd1 _18778_/CLK sky130_fd_sc_hd__inv_2
XFILLER_190_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12092_ _12018_/X _11974_/X _12091_/X _12016_/S vssd1 vssd1 vccd1 vccd1 _12092_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _15927_/A _17824_/Q _17823_/Q vssd1 vssd1 vccd1 vccd1 _15923_/C sky130_fd_sc_hd__o21ai_1
X_11043_ _11365_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11066_/S sky130_fd_sc_hd__nor2_2
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14802_/A vssd1 vssd1 vccd1 vccd1 _14802_/X sky130_fd_sc_hd__buf_1
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18570_ _18572_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _12992_/X _12994_/B vssd1 vssd1 vccd1 vccd1 _12995_/A sky130_fd_sc_hd__and2b_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17521_ _17737_/CLK _17521_/D vssd1 vssd1 vccd1 vccd1 _17521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14733_ _19082_/Q _18346_/Q _17580_/Q _18798_/Q _14568_/X _14569_/X vssd1 vssd1 vccd1
+ vccd1 _14734_/B sky130_fd_sc_hd__mux4_2
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11945_ _12022_/A vssd1 vssd1 vccd1 vccd1 _11945_/X sky130_fd_sc_hd__buf_2
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17452_ _17437_/X _17452_/B vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__and2b_1
X_14264__465 _14265__466/A vssd1 vssd1 vccd1 vccd1 _18100_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14664_ _14664_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14664_/Y sky130_fd_sc_hd__nand2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11876_ _11876_/A vssd1 vssd1 vccd1 vccd1 _11876_/X sky130_fd_sc_hd__buf_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _16412_/B _16403_/B vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__nand2_1
X_13615_ _13150_/X _13601_/X _13614_/Y _13604_/X vssd1 vssd1 vccd1 vccd1 _17849_/D
+ sky130_fd_sc_hd__a211oi_1
X_10827_ _18357_/Q _10806_/X _10831_/S vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__mux2_1
X_14595_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14595_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19122_ _19122_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
X_13546_ _13712_/A _13545_/B _13545_/Y _13472_/X vssd1 vssd1 vccd1 vccd1 _17827_/D
+ sky130_fd_sc_hd__a211oi_1
X_10758_ _18384_/Q _10698_/X _10762_/S vssd1 vssd1 vccd1 vccd1 _10759_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19053_ _19053_/CLK _19053_/D vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ _18749_/Q _18757_/Q _18765_/Q _18773_/Q _16149_/X _16150_/X vssd1 vssd1 vccd1
+ vccd1 _16265_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13477_ _17806_/Q _13477_/B vssd1 vssd1 vccd1 vccd1 _13477_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10689_ _10689_/A vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18004_ _18013_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
X_15216_ _19316_/Q _19300_/Q _19292_/Q _19267_/Q _15214_/X _15215_/X vssd1 vssd1 vccd1
+ vccd1 _15216_/X sky130_fd_sc_hd__mux4_1
X_12428_ _17611_/Q _17612_/Q _12440_/S vssd1 vssd1 vccd1 vccd1 _12428_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16196_ _18596_/Q _18612_/Q _18738_/Q _18519_/Q _16195_/X _16138_/X vssd1 vssd1 vccd1
+ vccd1 _16197_/B sky130_fd_sc_hd__mux4_1
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12359_ _12359_/A vssd1 vssd1 vccd1 vccd1 _12390_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1__f__04573_ clkbuf_0__04573_/X vssd1 vssd1 vccd1 vccd1 _16657__294/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15078_ _15076_/A _15075_/X _15077_/Y _14247_/X vssd1 vssd1 vccd1 vccd1 _18481_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ _13792_/X _14017_/A _14020_/X vssd1 vssd1 vccd1 vccd1 _14029_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18906_ _18906_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18837_ _18837_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11878__361 _11879__362/A vssd1 vssd1 vccd1 vccd1 _17508_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _18947_/Q _09492_/X _09572_/S vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__mux2_1
X_18768_ _18768_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ _17719_/CLK _17719_/D vssd1 vssd1 vccd1 vccd1 _17719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18699_ _18699_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04007_ clkbuf_0__04007_/X vssd1 vssd1 vccd1 vccd1 _15840__142/A sky130_fd_sc_hd__clkbuf_16
XFILLER_208_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ _18811_/Q hold17/A vssd1 vssd1 vccd1 vccd1 _09004_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__07559_ clkbuf_0__07559_/X vssd1 vssd1 vccd1 vccd1 _12344__404/A sky130_fd_sc_hd__clkbuf_16
XFILLER_219_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09906_ _09906_/A vssd1 vssd1 vccd1 vccd1 _18795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _18815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09768_ _18844_/Q _09767_/X _09768_/S vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09699_/A vssd1 vssd1 vccd1 vccd1 _18898_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11730_/A vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_215_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16357__248 _16358__249/A vssd1 vssd1 vccd1 vccd1 _18964_/CLK sky130_fd_sc_hd__inv_2
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _17512_/Q _09682_/A _11665_/S vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _13400_/A _13405_/B vssd1 vssd1 vccd1 vccd1 _13400_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ _10126_/X _18448_/Q _10612_/S vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14380_ _14380_/A vssd1 vssd1 vccd1 vccd1 _14380_/X sky130_fd_sc_hd__buf_1
X_11592_ _11592_/A vssd1 vssd1 vccd1 vccd1 _17577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ _13231_/X _13330_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13331_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ _10543_/A vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _16050_/A _16050_/B vssd1 vssd1 vccd1 vccd1 _16050_/Y sky130_fd_sc_hd__nand2_1
X_13262_ _17747_/Q _13252_/X _13261_/Y vssd1 vssd1 vccd1 vccd1 _17747_/D sky130_fd_sc_hd__o21a_1
XFILLER_157_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _10546_/A _10492_/B vssd1 vssd1 vccd1 vccd1 _10490_/S sky130_fd_sc_hd__nor2_2
XFILLER_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ _15001_/A _15001_/B vssd1 vssd1 vccd1 vccd1 _15002_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_0__f__05076_ clkbuf_0__05076_/X vssd1 vssd1 vccd1 vccd1 _17389__84/A sky130_fd_sc_hd__clkbuf_16
X_12213_ _17523_/Q _12212_/X _12202_/A _17521_/Q vssd1 vssd1 vccd1 vccd1 _12217_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_13193_ _17732_/Q _13208_/B vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15729__1019 _15729__1019/A vssd1 vssd1 vccd1 vccd1 _18736_/CLK sky130_fd_sc_hd__inv_2
XFILLER_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _12132_/X _12144_/B vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__and2b_1
XFILLER_124_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14532__681 _14532__681/A vssd1 vssd1 vccd1 vccd1 _18316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _12075_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12075_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16952_ _16892_/A _16951_/X _16860_/X vssd1 vssd1 vccd1 vccd1 _16952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_238_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11026_ _18266_/Q _09119_/X _11034_/S vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15903_ _17814_/Q _17813_/Q _15943_/B vssd1 vssd1 vccd1 vccd1 _15947_/A sky130_fd_sc_hd__or3_1
XFILLER_103_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16883_ _18181_/Q _18173_/Q _18165_/Q _18157_/Q _16881_/X _16882_/X vssd1 vssd1 vccd1
+ vccd1 _16884_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18622_ _18622_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452__942 _15454__944/A vssd1 vssd1 vccd1 vccd1 _18629_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03171_ clkbuf_0__03171_/X vssd1 vssd1 vccd1 vccd1 _14391__567/A sky130_fd_sc_hd__clkbuf_16
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18553_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
X_12977_ _12975_/X _12977_/B vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__and2b_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11928_ _19223_/Q vssd1 vssd1 vccd1 vccd1 _17129_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14716_ _17587_/Q _18385_/Q _18393_/Q _18427_/Q _14574_/X _14637_/X vssd1 vssd1 vccd1
+ vccd1 _14717_/B sky130_fd_sc_hd__mux4_2
X_18484_ _18484_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _17356_/X _17435_/B vssd1 vssd1 vccd1 vccd1 _17436_/A sky130_fd_sc_hd__and2b_1
X_14647_ _18325_/Q _14543_/X _14623_/X _14646_/X vssd1 vssd1 vccd1 vccd1 _18325_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11859_ _13820_/A _11865_/B _11859_/C vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__and3_1
XFILLER_61_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17366_ _19283_/Q _12212_/X _12202_/X _19281_/Q vssd1 vssd1 vccd1 vccd1 _17366_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14578_ _19048_/Q vssd1 vssd1 vccd1 vccd1 _14696_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19105_ _19105_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_1
X_13529_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13529_/X sky130_fd_sc_hd__buf_4
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19036_ _19037_/CLK _19036_/D vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfxtp_1
X_16248_ _16246_/X _16247_/X _16248_/S vssd1 vssd1 vccd1 vccd1 _16248_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 _17890_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput114 _19385_/X vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_2
XFILLER_173_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _18713_/Q _18721_/Q _18729_/Q _18494_/Q _16149_/X _16150_/X vssd1 vssd1 vccd1
+ vccd1 _16179_/X sky130_fd_sc_hd__mux4_1
Xoutput125 _19390_/X vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_2
XFILLER_154_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput136 _19387_/X vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_2
X_14314__506 _14314__506/A vssd1 vssd1 vccd1 vccd1 _18141_/CLK sky130_fd_sc_hd__inv_2
XFILLER_217_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput147 _11849_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput158 _11820_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_88_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__04587_ _16707_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04587_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_247_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09622_ _09615_/X _09622_/B _09649_/C vssd1 vssd1 vccd1 vccd1 _09623_/A sky130_fd_sc_hd__and3b_1
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09553_ _09553_/A vssd1 vssd1 vccd1 vccd1 _18955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09484_ _19012_/Q _09481_/X _09496_/S vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15780__1060 _15782__1062/A vssd1 vssd1 vccd1 vccd1 _18777_/CLK sky130_fd_sc_hd__inv_2
XFILLER_212_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14475__635 _14476__636/A vssd1 vssd1 vccd1 vccd1 _18270_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03191_ clkbuf_0__03191_/X vssd1 vssd1 vccd1 vccd1 _14498__654/A sky130_fd_sc_hd__clkbuf_16
X_14887__803 _14888__804/A vssd1 vssd1 vccd1 vccd1 _18448_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19246_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10190_ _18690_/Q _10189_/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _12894_/X _12900_/B vssd1 vssd1 vccd1 vccd1 _12901_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13880_ _13880_/A vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17065__52 _17066__53/A vssd1 vssd1 vccd1 vccd1 _19201_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ _17651_/Q _17984_/Q _12831_/S vssd1 vssd1 vccd1 vccd1 _12832_/B sky130_fd_sc_hd__mux2_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15557_/B _15557_/C vssd1 vssd1 vccd1 vccd1 _15562_/C sky130_fd_sc_hd__and2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12762_/A vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__buf_2
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04576_ clkbuf_0__04576_/X vssd1 vssd1 vccd1 vccd1 _16674__308/A sky130_fd_sc_hd__clkbuf_16
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15481_ _18656_/Q _15482_/B vssd1 vssd1 vccd1 vccd1 _15481_/Y sky130_fd_sc_hd__nand2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _17615_/D sky130_fd_sc_hd__nor2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17225_/C _17225_/D vssd1 vssd1 vccd1 vccd1 _17222_/A sky130_fd_sc_hd__and2_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11644_/A vssd1 vssd1 vccd1 vccd1 _17537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17151_ _11978_/X _17142_/X _19229_/Q vssd1 vssd1 vccd1 vccd1 _17152_/C sky130_fd_sc_hd__a21o_1
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 io_in[26] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_6
X_11575_ _17584_/Q _10901_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__mux2_1
Xinput27 vga_g[1] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_8
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16102_ _16172_/A vssd1 vssd1 vccd1 vccd1 _16102_/X sky130_fd_sc_hd__clkbuf_4
X_13314_ _13192_/X _13311_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _13314_/Y sky130_fd_sc_hd__a21oi_1
Xinput38 wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_2
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
X_10526_ _18516_/Q _10351_/X _10526_/S vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _14300_/A vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__buf_1
X_14788__723 _14789__724/A vssd1 vssd1 vccd1 vccd1 _18366_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _16033_/A _16033_/B vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__nor2_1
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13245_ _13244_/X _13232_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _13245_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10457_ _10472_/S vssd1 vssd1 vccd1 vccd1 _10466_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_237_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13176_ _13170_/X _13173_/X _13175_/Y _13158_/X vssd1 vssd1 vccd1 vccd1 _17729_/D
+ sky130_fd_sc_hd__a211oi_1
X_10388_ _08804_/X _18577_/Q _10388_/S vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _11888_/X _12127_/B vssd1 vssd1 vccd1 vccd1 _12128_/A sky130_fd_sc_hd__and2b_1
X_17984_ _17991_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 _17984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04372_ _16333_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04372_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12058_ _19221_/Q vssd1 vssd1 vccd1 vccd1 _17117_/B sky130_fd_sc_hd__clkbuf_2
X_16935_ _19141_/Q _16797_/X _16934_/X _16915_/X vssd1 vssd1 vccd1 vccd1 _19141_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105__411 _13106__412/A vssd1 vssd1 vccd1 vccd1 _17707_/CLK sky130_fd_sc_hd__inv_2
XFILLER_226_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ _11009_/A vssd1 vssd1 vccd1 vccd1 _18274_/D sky130_fd_sc_hd__clkbuf_1
X_16866_ _16864_/X _16865_/X _16982_/A vssd1 vssd1 vccd1 vccd1 _16866_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18605_ _18605_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03154_ clkbuf_0__03154_/X vssd1 vssd1 vccd1 vccd1 _14311__504/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15817_ _18889_/Q vssd1 vssd1 vccd1 vccd1 _16049_/A sky130_fd_sc_hd__inv_2
XFILLER_19_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16797_ _16797_/A vssd1 vssd1 vccd1 vccd1 _16797_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03185_ _14462_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03185_/X sky130_fd_sc_hd__clkbuf_16
X_18536_ _18536_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
X_15748_ _15748_/A vssd1 vssd1 vccd1 vccd1 _15748_/X sky130_fd_sc_hd__buf_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18467_ _18482_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18398_ _18398_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349_ _17349_/A vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14539__687 _14539__687/A vssd1 vssd1 vccd1 vccd1 _18322_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03987_ clkbuf_0__03987_/X vssd1 vssd1 vccd1 vccd1 _15782__1062/A sky130_fd_sc_hd__clkbuf_16
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19019_ _19027_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15459__948 _15460__949/A vssd1 vssd1 vccd1 vccd1 _18635_/CLK sky130_fd_sc_hd__inv_2
XFILLER_170_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08984_ _19214_/Q _08961_/X _08988_/S vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14882__799 _14882__799/A vssd1 vssd1 vccd1 vccd1 _18444_/CLK sky130_fd_sc_hd__inv_2
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09605_ _09605_/A vssd1 vssd1 vccd1 vccd1 _15291_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15846__147 _15846__147/A vssd1 vssd1 vccd1 vccd1 _18822_/CLK sky130_fd_sc_hd__inv_2
X_09536_ _18962_/Q _09495_/X _09536_/S vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _16559_/B _09467_/B vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__nand2_8
X_15728__1018 _15729__1019/A vssd1 vssd1 vccd1 vccd1 _18735_/CLK sky130_fd_sc_hd__inv_2
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09398_ _08910_/X _19066_/Q _09406_/S vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11360_/A vssd1 vssd1 vccd1 vccd1 _18133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03174_ clkbuf_0__03174_/X vssd1 vssd1 vccd1 vccd1 _14411__584/A sky130_fd_sc_hd__clkbuf_16
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10326_/S vssd1 vssd1 vccd1 vccd1 _10320_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11291_ _18160_/Q _11267_/X _11295_/S vssd1 vssd1 vccd1 vccd1 _11292_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13030_ _12992_/X _13030_/B vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10242_ _18639_/Q _10180_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _18695_/Q _10072_/X _10173_/S vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14981_ _14986_/B _14981_/B vssd1 vssd1 vccd1 vccd1 _14981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_248_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _17954_/Q _13941_/B vssd1 vssd1 vccd1 vccd1 _13932_/Y sky130_fd_sc_hd__nor2_1
X_17038__30 _17039__31/A vssd1 vssd1 vccd1 vccd1 _19179_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13863_ _14081_/A _13863_/B vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12814_ _12812_/X _12814_/B vssd1 vssd1 vccd1 vccd1 _12815_/A sky130_fd_sc_hd__and2b_1
X_15602_ _18654_/Q _15612_/B vssd1 vssd1 vccd1 vccd1 _15602_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16582_ _19022_/Q _16585_/C _16564_/X vssd1 vssd1 vccd1 vccd1 _16582_/Y sky130_fd_sc_hd__a21oi_1
X_13794_ _17908_/Q _13771_/X _13793_/Y vssd1 vssd1 vccd1 vccd1 _17908_/D sky130_fd_sc_hd__o21a_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18321_ _18321_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
X_12745_ _12745_/A _12745_/B vssd1 vssd1 vccd1 vccd1 _17631_/D sky130_fd_sc_hd__nor2_1
XFILLER_231_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15533_ _15643_/B _15642_/B vssd1 vssd1 vccd1 vccd1 _15583_/A sky130_fd_sc_hd__or2_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _18252_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
X_12676_ _12676_/A vssd1 vssd1 vccd1 vccd1 _17610_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17203_ _19243_/Q _19242_/Q _17203_/C _17203_/D vssd1 vssd1 vccd1 vccd1 _17216_/C
+ sky130_fd_sc_hd__and4_1
X_11627_ _17544_/Q _09685_/A _11629_/S vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18183_ _18183_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17134_ _17149_/C vssd1 vssd1 vccd1 vccd1 _17142_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _11558_/A vssd1 vssd1 vccd1 vccd1 _17707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _10509_/A vssd1 vssd1 vccd1 vccd1 _18524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11489_ _09142_/X _18049_/Q _11491_/S vssd1 vssd1 vccd1 vccd1 _11490_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16016_ _16014_/Y _16015_/Y _16010_/X vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__a21oi_1
X_13228_ _13441_/A vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__buf_4
XFILLER_98_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13159_ _13135_/X _13155_/X _13156_/Y _13158_/X vssd1 vssd1 vccd1 vccd1 _17726_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_135_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _19039_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16918_ _18151_/Q _18143_/Q _18135_/Q _18279_/Q _16803_/X _16804_/X vssd1 vssd1 vccd1
+ vccd1 _16918_/X sky130_fd_sc_hd__mux4_1
X_17898_ _17923_/CLK _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_226_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16849_ _16881_/A vssd1 vssd1 vccd1 vccd1 _16849_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_225_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09321_ _09336_/S vssd1 vssd1 vccd1 vccd1 _09330_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18519_ _18519_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03168_ _14380_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03168_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_206_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09252_ _09252_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__nor2_4
XFILLER_221_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _09183_/A vssd1 vssd1 vccd1 vccd1 _19165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15656__960 _15657__961/A vssd1 vssd1 vccd1 vccd1 _18677_/CLK sky130_fd_sc_hd__inv_2
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08967_ _09697_/A vssd1 vssd1 vccd1 vccd1 _08967_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ _08898_/A vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14327__516 _14329__518/A vssd1 vssd1 vccd1 vccd1 _18151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10860_ _10860_/A vssd1 vssd1 vccd1 vccd1 _18343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09519_ _09519_/A vssd1 vssd1 vccd1 vccd1 _19000_/D sky130_fd_sc_hd__clkbuf_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10791_ _10813_/S vssd1 vssd1 vccd1 vccd1 _10804_/S sky130_fd_sc_hd__buf_2
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12530_ _17629_/Q _17630_/Q _17631_/Q _17632_/Q _12443_/X _12429_/S vssd1 vssd1 vccd1
+ vccd1 _12530_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_61_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _18024_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12768_/S vssd1 vssd1 vccd1 vccd1 _12567_/S sky130_fd_sc_hd__buf_2
XFILLER_200_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _14200_/A vssd1 vssd1 vccd1 vccd1 _18071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11412_ _11335_/X _18110_/Q _11412_/S vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__mux2_1
X_15180_ _15642_/A vssd1 vssd1 vccd1 vccd1 _15190_/B sky130_fd_sc_hd__inv_2
X_12392_ _12392_/A vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_166_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ _18028_/Q _14115_/X _14130_/Y vssd1 vssd1 vccd1 vccd1 _18028_/D sky130_fd_sc_hd__o21a_1
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11343_ _11343_/A vssd1 vssd1 vccd1 vccd1 _18140_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03157_ clkbuf_0__03157_/X vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__clkbuf_16
X_14062_ _18002_/Q _14054_/X _14061_/Y vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__o21a_1
X_11274_ _18166_/Q _11273_/X _11274_/S vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__mux2_1
X_13013_ _17676_/Q _12924_/X _12920_/X _17678_/Q vssd1 vssd1 vccd1 vccd1 _13020_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_10225_ _10225_/A vssd1 vssd1 vccd1 vccd1 _18677_/D sky130_fd_sc_hd__clkbuf_1
X_18870_ _18870_/CLK _18870_/D vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_1
X_14488__645 _14490__647/A vssd1 vssd1 vccd1 vccd1 _18280_/CLK sky130_fd_sc_hd__inv_2
X_17821_ _19147_/CLK _17821_/D vssd1 vssd1 vccd1 vccd1 _17821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ _10156_/A vssd1 vssd1 vccd1 vccd1 _18703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_248_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17752_ _19327_/CLK _17752_/D vssd1 vssd1 vccd1 vccd1 _17752_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14964_ _14964_/A _14964_/B _14964_/C _14964_/D vssd1 vssd1 vccd1 vccd1 _14965_/B
+ sky130_fd_sc_hd__or4_1
X_10087_ _10087_/A vssd1 vssd1 vccd1 vccd1 _18730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13915_ _17948_/Q _13902_/X _13914_/Y vssd1 vssd1 vccd1 vccd1 _17948_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17683_ _17703_/CLK _17683_/D vssd1 vssd1 vccd1 vccd1 _17683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ _18453_/Q _15059_/A _14894_/Y vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__a21o_1
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13846_ input73/X _13845_/B _13845_/Y _13841_/X vssd1 vssd1 vccd1 vccd1 _17926_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16565_ _16567_/A _19016_/Q _16564_/X vssd1 vssd1 vccd1 vccd1 _16565_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_188_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13777_ _13777_/A vssd1 vssd1 vccd1 vccd1 _13777_/X sky130_fd_sc_hd__clkbuf_4
X_10989_ _11004_/S vssd1 vssd1 vccd1 vccd1 _10998_/S sky130_fd_sc_hd__clkbuf_2
X_18304_ _18304_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
X_15516_ _17839_/Q _15516_/B vssd1 vssd1 vccd1 vccd1 _15517_/C sky130_fd_sc_hd__nand2_1
X_12728_ _12727_/A _12726_/A _12718_/X vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__o21ai_1
X_19284_ _19288_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ _18982_/Q _16497_/B vssd1 vssd1 vccd1 vccd1 _16498_/B sky130_fd_sc_hd__nor2_1
XFILLER_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18235_ _18235_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
X_12659_ _12387_/X _12658_/A _17606_/Q vssd1 vssd1 vccd1 vccd1 _12660_/C sky130_fd_sc_hd__a21o_1
XFILLER_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15447_ _15447_/A vssd1 vssd1 vccd1 vccd1 _15447_/X sky130_fd_sc_hd__buf_1
XFILLER_175_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18166_ _18166_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_1
X_15795__116 _15796__117/A vssd1 vssd1 vccd1 vccd1 _18788_/CLK sky130_fd_sc_hd__inv_2
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ _19074_/Q _19066_/Q _19058_/Q _19012_/Q _15208_/A _09605_/A vssd1 vssd1 vccd1
+ vccd1 _15379_/A sky130_fd_sc_hd__mux4_1
XFILLER_184_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17117_ _17117_/A _17117_/B _17117_/C vssd1 vssd1 vccd1 vccd1 _17118_/C sky130_fd_sc_hd__nand3_1
XFILLER_117_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18097_ _18097_/CLK _18097_/D vssd1 vssd1 vccd1 vccd1 _18097_/Q sky130_fd_sc_hd__dfxtp_1
X_14432__600 _14434__602/A vssd1 vssd1 vccd1 vccd1 _18235_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _15808_/B vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15727__1017 _15727__1017/A vssd1 vssd1 vccd1 vccd1 _18734_/CLK sky130_fd_sc_hd__inv_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14389__565 _14391__567/A vssd1 vssd1 vccd1 vccd1 _18200_/CLK sky130_fd_sc_hd__inv_2
XFILLER_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18999_ _18999_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_18 _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_29 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ hold14/X vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17032__25 _17033__26/A vssd1 vssd1 vccd1 vccd1 _19174_/CLK sky130_fd_sc_hd__inv_2
XFILLER_179_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _08910_/X _19107_/Q _09312_/S vssd1 vssd1 vccd1 vccd1 _09305_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13118__421 _13120__423/A vssd1 vssd1 vccd1 vccd1 _17717_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ _09235_/A _18562_/Q vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__and2_1
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ _19172_/Q _09116_/X _09166_/S vssd1 vssd1 vccd1 vccd1 _09167_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09097_ _19193_/Q _09096_/X _09105_/S vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10010_ _18759_/Q _09967_/X _10010_/S vssd1 vssd1 vccd1 vccd1 _10011_/A sky130_fd_sc_hd__mux2_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _18765_/D sky130_fd_sc_hd__clkbuf_1
X_15396__898 _15397__899/A vssd1 vssd1 vccd1 vccd1 _18585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11961_ _12007_/S vssd1 vssd1 vccd1 vccd1 _11961_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13880_/A sky130_fd_sc_hd__clkbuf_2
X_10912_ _10912_/A vssd1 vssd1 vccd1 vccd1 _18315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _18589_/Q _18303_/Q _17569_/Q _18840_/Q _14615_/X _14641_/X vssd1 vssd1 vccd1
+ vccd1 _14680_/X sky130_fd_sc_hd__mux4_1
X_11892_ _17216_/B _19247_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ _17855_/Q _13635_/B vssd1 vssd1 vccd1 vccd1 _13631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10843_ _18350_/Q _10803_/X _10843_/S vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ _17832_/Q _13568_/B vssd1 vssd1 vccd1 vccd1 _13562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10774_ _10774_/A vssd1 vssd1 vccd1 vccd1 _18378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12513_ _12717_/A _17624_/Q _17625_/Q _17626_/Q _12555_/A _12441_/S vssd1 vssd1 vccd1
+ vccd1 _12513_/X sky130_fd_sc_hd__mux4_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15301_ _15301_/A vssd1 vssd1 vccd1 vccd1 _15301_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16281_ _18452_/Q _19090_/Q _19127_/Q _18436_/Q _16106_/X _16108_/X vssd1 vssd1 vccd1
+ vccd1 _16281_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _13493_/A vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__buf_4
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18020_ _18021_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12444_ _18011_/Q vssd1 vssd1 vccd1 vccd1 _12464_/S sky130_fd_sc_hd__clkbuf_2
X_15232_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _15232_/X sky130_fd_sc_hd__buf_2
X_12340__400 _12344__404/A vssd1 vssd1 vccd1 vccd1 _17581_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12375_ _17610_/Q _17611_/Q _12443_/A vssd1 vssd1 vccd1 vccd1 _12375_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14114_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__clkbuf_2
X_11326_ _11326_/A vssd1 vssd1 vccd1 vccd1 _11326_/X sky130_fd_sc_hd__clkbuf_2
X_15094_ _15100_/A vssd1 vssd1 vccd1 vccd1 _15094_/X sky130_fd_sc_hd__buf_1
XFILLER_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16705__328 _16706__329/A vssd1 vssd1 vccd1 vccd1 _19103_/CLK sky130_fd_sc_hd__inv_2
X_14045_ _17996_/Q _14032_/X _14044_/Y vssd1 vssd1 vccd1 vccd1 _17996_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18922_ _18922_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11257_ _11165_/X _18171_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11258_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10208_ _10208_/A vssd1 vssd1 vccd1 vccd1 _18684_/D sky130_fd_sc_hd__clkbuf_1
X_18853_ _18853_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_1
X_11188_ _18202_/Q _11042_/X _11196_/S vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17804_ _19135_/CLK _17804_/D vssd1 vssd1 vccd1 vccd1 _17804_/Q sky130_fd_sc_hd__dfxtp_1
X_10139_ _10528_/B _10620_/B vssd1 vssd1 vccd1 vccd1 _10155_/S sky130_fd_sc_hd__nor2_2
XFILLER_212_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18784_ _18784_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15996_ _16002_/B _16002_/C _15963_/X vssd1 vssd1 vccd1 vccd1 _15996_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _19147_/CLK _17735_/D vssd1 vssd1 vccd1 vccd1 _17735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14947_ _14940_/A _17858_/Q _17857_/Q vssd1 vssd1 vccd1 vccd1 _14948_/B sky130_fd_sc_hd__o21ai_1
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17666_ _19027_/CLK _17666_/D vssd1 vssd1 vccd1 vccd1 _17666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_100 _11755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_111 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_122 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_133 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16617_ _19037_/Q _16614_/B _16616_/Y vssd1 vssd1 vccd1 vccd1 _19037_/D sky130_fd_sc_hd__o21a_1
XFILLER_90_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_144 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ _13829_/A vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__clkbuf_2
X_17597_ _17602_/CLK _17597_/D vssd1 vssd1 vccd1 vccd1 _17597_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_155 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_166 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19336_ _19336_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_177 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_188 _09861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_199 _11846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15803__123 _15804__124/A vssd1 vssd1 vccd1 vccd1 _18795_/CLK sky130_fd_sc_hd__inv_2
X_19267_ _19267_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
X_16479_ _18978_/Q _16440_/A _16478_/Y _16427_/X vssd1 vssd1 vccd1 vccd1 _16480_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09020_ _11457_/A vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__clkbuf_4
X_18218_ _18218_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19198_ _19198_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18149_ _18149_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03807_ clkbuf_0__03807_/X vssd1 vssd1 vccd1 vccd1 _15453__943/A sky130_fd_sc_hd__clkbuf_16
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _18788_/Q _09265_/X _09926_/S vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09853_ _18807_/Q vssd1 vssd1 vccd1 vccd1 _16893_/A sky130_fd_sc_hd__clkbuf_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _18880_/Q vssd1 vssd1 vccd1 vccd1 _08804_/X sky130_fd_sc_hd__clkbuf_2
X_09784_ _09784_/A vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08735_ _13540_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__nor2_2
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172__878 _15172__878/A vssd1 vssd1 vccd1 vccd1 _18554_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16095__207 _16096__208/A vssd1 vssd1 vccd1 vccd1 _18912_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14439__606 _14440__607/A vssd1 vssd1 vccd1 vccd1 _18241_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ _09218_/A vssd1 vssd1 vccd1 vccd1 _19150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _18532_/Q _10351_/X _10490_/S vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09149_ _11565_/A vssd1 vssd1 vccd1 vccd1 _10691_/B sky130_fd_sc_hd__buf_4
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _17525_/Q _17726_/Q _12170_/S vssd1 vssd1 vccd1 vccd1 _12161_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _11111_/A vssd1 vssd1 vccd1 vccd1 _18233_/D sky130_fd_sc_hd__clkbuf_1
X_12091_ _12091_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12091_/X sky130_fd_sc_hd__or2_1
X_14782__718 _14782__718/A vssd1 vssd1 vccd1 vccd1 _18361_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _18668_/Q vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__buf_2
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _17954_/Q _17683_/Q _12993_/S vssd1 vssd1 vccd1 vccd1 _12994_/B sky130_fd_sc_hd__mux2_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _19339_/CLK _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _14732_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14732_/Y sky130_fd_sc_hd__nor2_1
X_11944_ _11944_/A vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669__970 _15671__972/A vssd1 vssd1 vccd1 vccd1 _18687_/CLK sky130_fd_sc_hd__inv_2
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17451_ _17744_/Q _19332_/Q _17451_/S vssd1 vssd1 vccd1 vccd1 _17452_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _14659_/X _14662_/X _14730_/S vssd1 vssd1 vccd1 vccd1 _14664_/B sky130_fd_sc_hd__mux2_2
X_11875_ _17421_/A vssd1 vssd1 vccd1 vccd1 _11875_/X sky130_fd_sc_hd__buf_1
XFILLER_233_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _17805_/Q _16402_/B vssd1 vssd1 vccd1 vccd1 _16403_/B sky130_fd_sc_hd__nand2_1
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13614_ _17849_/Q _13621_/B vssd1 vssd1 vccd1 vccd1 _13614_/Y sky130_fd_sc_hd__nor2_1
X_10826_ _10826_/A vssd1 vssd1 vccd1 vccd1 _18358_/D sky130_fd_sc_hd__clkbuf_1
X_17382_ _17382_/A vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__clkbuf_1
X_14594_ _14594_/A vssd1 vssd1 vccd1 vccd1 _14594_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15726__1016 _15727__1017/A vssd1 vssd1 vccd1 vccd1 _18733_/CLK sky130_fd_sc_hd__inv_2
X_19121_ _19121_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ _16333_/A vssd1 vssd1 vccd1 vccd1 _16333_/X sky130_fd_sc_hd__buf_1
X_15446__939 _15446__939/A vssd1 vssd1 vccd1 vccd1 _18626_/CLK sky130_fd_sc_hd__inv_2
X_13545_ _17827_/Q _13545_/B vssd1 vssd1 vccd1 vccd1 _13545_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10757_ _10757_/A vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19052_ _19052_/CLK _19052_/D vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16264_ _16191_/X _16257_/Y _16259_/Y _16261_/Y _16263_/Y vssd1 vssd1 vccd1 vccd1
+ _16264_/X sky130_fd_sc_hd__o32a_2
X_13476_ _16058_/A _13463_/B _13475_/Y _13472_/X vssd1 vssd1 vccd1 vccd1 _17805_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_200_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10688_ _18413_/Q _09741_/X _10688_/S vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__mux2_1
X_18003_ _18014_/CLK _18003_/D vssd1 vssd1 vccd1 vccd1 _18003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12427_ _12435_/A vssd1 vssd1 vccd1 vccd1 _12440_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15215_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15215_/X sky130_fd_sc_hd__buf_2
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16195_ _16195_/A vssd1 vssd1 vccd1 vccd1 _16195_/X sky130_fd_sc_hd__buf_2
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12358_ _18011_/Q vssd1 vssd1 vccd1 vccd1 _12359_/A sky130_fd_sc_hd__buf_2
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04572_ clkbuf_0__04572_/X vssd1 vssd1 vccd1 vccd1 _16649__287/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _11150_/X _18152_/Q _11313_/S vssd1 vssd1 vccd1 vccd1 _11310_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15077_ _15079_/B vssd1 vssd1 vccd1 vccd1 _15077_/Y sky130_fd_sc_hd__inv_2
X_12289_ _12289_/A vssd1 vssd1 vccd1 vccd1 _17561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ _17990_/Q _14012_/X _14027_/Y vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__o21a_1
X_18905_ _18905_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18836_ _18836_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18767_ _18767_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
X_15979_ _15985_/B _15985_/C _15963_/X vssd1 vssd1 vccd1 vccd1 _15979_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_247_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17718_ _17718_/CLK _17718_/D vssd1 vssd1 vccd1 vccd1 _17718_/Q sky130_fd_sc_hd__dfxtp_1
X_18698_ _18698_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04006_ clkbuf_0__04006_/X vssd1 vssd1 vccd1 vccd1 _15833__136/A sky130_fd_sc_hd__clkbuf_16
X_17649_ _18012_/CLK _17649_/D vssd1 vssd1 vccd1 vccd1 _17649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12347__406 _12348__407/A vssd1 vssd1 vccd1 vccd1 _17587_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17389__84 _17389__84/A vssd1 vssd1 vccd1 vccd1 _19297_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19319_ _19319_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09003_ hold22/A hold26/A _18802_/Q vssd1 vssd1 vccd1 vccd1 _09011_/A sky130_fd_sc_hd__and3_1
XFILLER_247_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04839_ clkbuf_0__04839_/X vssd1 vssd1 vccd1 vccd1 _17018__14/A sky130_fd_sc_hd__clkbuf_16
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11885__366 _11886__367/A vssd1 vssd1 vccd1 vccd1 _17513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_191_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__07558_ clkbuf_0__07558_/X vssd1 vssd1 vccd1 vccd1 _12338__399/A sky130_fd_sc_hd__clkbuf_16
XFILLER_144_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09905_ _18795_/Q _09729_/X _09907_/S vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _09688_/X _18815_/Q _09836_/S vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17077__61 _17078__62/A vssd1 vssd1 vccd1 vccd1 _19210_/CLK sky130_fd_sc_hd__inv_2
XFILLER_246_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09767_ _18880_/Q vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__buf_2
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09697_/X _18898_/Q _09698_/S vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04592_ clkbuf_0__04592_/X vssd1 vssd1 vccd1 vccd1 _16999__349/A sky130_fd_sc_hd__clkbuf_16
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11660_ _11660_/A vssd1 vssd1 vccd1 vccd1 _17513_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10611_ _10611_/A vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11591_ _17577_/Q _10701_/A _11593_/S vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13330_ _13330_/A vssd1 vssd1 vccd1 vccd1 _13330_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10542_ _18509_/Q _10348_/X _10544_/S vssd1 vssd1 vccd1 vccd1 _10543_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _13184_/X _13259_/X _13260_/X vssd1 vssd1 vccd1 vccd1 _13261_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10473_ _10473_/A vssd1 vssd1 vccd1 vccd1 _18540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12212_ _12212_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__clkbuf_2
X_15000_ _18459_/Q _14991_/X _14999_/Y _14993_/X vssd1 vssd1 vccd1 vccd1 _15001_/B
+ sky130_fd_sc_hd__a22o_1
X_12224__370 _12226__372/A vssd1 vssd1 vccd1 vccd1 _17534_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13192_ _14079_/A vssd1 vssd1 vccd1 vccd1 _13192_/X sky130_fd_sc_hd__buf_6
XFILLER_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12143_ _17520_/Q _17731_/Q _12153_/S vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16628__270 _16631__273/A vssd1 vssd1 vccd1 vccd1 _19044_/CLK sky130_fd_sc_hd__inv_2
XFILLER_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12074_ _11977_/X _11953_/X _12091_/A vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__mux2_1
X_16951_ _16836_/X _16944_/Y _16946_/Y _16948_/Y _16950_/Y vssd1 vssd1 vccd1 vccd1
+ _16951_/X sky130_fd_sc_hd__o32a_1
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14270__470 _14271__471/A vssd1 vssd1 vccd1 vccd1 _18105_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11025_ _11040_/S vssd1 vssd1 vccd1 vccd1 _11034_/S sky130_fd_sc_hd__clkbuf_2
X_15902_ _18872_/Q _15902_/B vssd1 vssd1 vccd1 vccd1 _15945_/A sky130_fd_sc_hd__xnor2_1
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16882_ _16882_/A vssd1 vssd1 vccd1 vccd1 _16882_/X sky130_fd_sc_hd__buf_2
XFILLER_38_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18621_ _18621_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03170_ clkbuf_0__03170_/X vssd1 vssd1 vccd1 vccd1 _14412_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18552_ _18552_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _17959_/Q _17678_/Q _12976_/S vssd1 vssd1 vccd1 vccd1 _12977_/B sky130_fd_sc_hd__mux2_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14734_/A _14715_/B vssd1 vssd1 vccd1 vccd1 _14715_/Y sky130_fd_sc_hd__nor2_1
X_11927_ _11923_/X _11926_/X _12076_/S vssd1 vssd1 vccd1 vccd1 _11927_/X sky130_fd_sc_hd__mux2_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _19108_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _17749_/Q _19327_/Q _17497_/B vssd1 vssd1 vccd1 vccd1 _17435_/B sky130_fd_sc_hd__mux2_1
XFILLER_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14646_ _09433_/X _14631_/X _14645_/Y vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__a21o_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11858_ _17919_/Q _11802_/A _11812_/A _17900_/Q vssd1 vssd1 vccd1 vccd1 _11859_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17365_ _19280_/Q _17478_/B vssd1 vssd1 vccd1 vccd1 _17365_/X sky130_fd_sc_hd__or2_1
X_10809_ _18988_/Q vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_158_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11789_ _11837_/A _13278_/B vssd1 vssd1 vccd1 vccd1 _11821_/B sky130_fd_sc_hd__or2_1
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14577_ _14736_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14577_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19104_ _19104_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13528_ _16530_/A _13522_/X _13526_/X _17820_/Q _15083_/B vssd1 vssd1 vccd1 vccd1
+ _17820_/D sky130_fd_sc_hd__a221o_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19035_ _19037_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _18716_/Q _18724_/Q _18732_/Q _18497_/Q _16205_/X _16206_/X vssd1 vssd1 vccd1
+ vccd1 _16247_/X sky130_fd_sc_hd__mux4_2
XFILLER_51_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ _14072_/A vssd1 vssd1 vccd1 vccd1 _16061_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput104 _19388_/X vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_2
XFILLER_161_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput115 _11741_/X vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_2
X_16178_ _18745_/Q _18753_/Q _18761_/Q _18769_/Q _16127_/X _16128_/X vssd1 vssd1 vccd1
+ vccd1 _16178_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput126 _19391_/X vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_2
XFILLER_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput137 _19398_/X vssd1 vssd1 vccd1 vccd1 jtag_tck sky130_fd_sc_hd__buf_2
Xoutput148 _11852_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_141_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput159 _11823_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15123__839 _15123__839/A vssd1 vssd1 vccd1 vccd1 _18515_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04586_ _16701_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04586_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15650__955 _15651__956/A vssd1 vssd1 vccd1 vccd1 _18672_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09621_ _16294_/B vssd1 vssd1 vccd1 vccd1 _09649_/C sky130_fd_sc_hd__clkbuf_2
X_18819_ _18819_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09552_ _08925_/X _18955_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03399_ _14759_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03399_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09483_ _09505_/S vssd1 vssd1 vccd1 vccd1 _09496_/S sky130_fd_sc_hd__buf_2
XFILLER_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03190_ clkbuf_0__03190_/X vssd1 vssd1 vccd1 vccd1 _14492__649/A sky130_fd_sc_hd__clkbuf_16
XFILLER_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15710__1004 _15710__1004/A vssd1 vssd1 vccd1 vccd1 _18721_/CLK sky130_fd_sc_hd__inv_2
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19136_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15725__1015 _15727__1017/A vssd1 vssd1 vccd1 vccd1 _18732_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09819_ _09819_/A vssd1 vssd1 vccd1 vccd1 _18823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12830_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12812_/A vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04575_ clkbuf_0__04575_/X vssd1 vssd1 vccd1 vccd1 _16666__301/A sky130_fd_sc_hd__clkbuf_16
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11712_ _17908_/Q _18088_/Q _17843_/Q vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__mux2_8
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _17615_/Q _12687_/X _12663_/X vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__o21ai_1
X_15480_ _17828_/Q _15529_/B vssd1 vssd1 vccd1 vccd1 _15482_/B sky130_fd_sc_hd__xnor2_1
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11643_ _08789_/X _17537_/Q _11647_/S vssd1 vssd1 vccd1 vccd1 _11644_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14431_ _14443_/A vssd1 vssd1 vccd1 vccd1 _14431_/X sky130_fd_sc_hd__buf_1
XFILLER_230_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17150_ _17239_/A vssd1 vssd1 vccd1 vccd1 _17189_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11574_ _11574_/A vssd1 vssd1 vccd1 vccd1 _17585_/D sky130_fd_sc_hd__clkbuf_1
X_14362_ _14380_/A vssd1 vssd1 vccd1 vccd1 _14362_/X sky130_fd_sc_hd__buf_1
Xinput17 io_in[27] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_6
XFILLER_168_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput28 vga_hsync vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_12
X_16101_ _16276_/A vssd1 vssd1 vccd1 vccd1 _16280_/A sky130_fd_sc_hd__clkbuf_2
X_13313_ _17763_/Q _13303_/X _13312_/Y vssd1 vssd1 vccd1 vccd1 _17763_/D sky130_fd_sc_hd__o21a_1
Xinput39 wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17383__79 _17383__79/A vssd1 vssd1 vccd1 vccd1 _19292_/CLK sky130_fd_sc_hd__inv_2
X_10525_ _10525_/A vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__clkbuf_1
X_14376__556 _14379__559/A vssd1 vssd1 vccd1 vccd1 _18191_/CLK sky130_fd_sc_hd__inv_2
X_17081_ _17081_/A vssd1 vssd1 vccd1 vccd1 _17081_/X sky130_fd_sc_hd__buf_1
X_14293_ _14293_/A vssd1 vssd1 vccd1 vccd1 _14293_/X sky130_fd_sc_hd__buf_1
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ _13732_/A vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__buf_4
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16032_ _15986_/A _16035_/C _16031_/Y _16035_/B _15949_/Y vssd1 vssd1 vccd1 vccd1
+ _16033_/B sky130_fd_sc_hd__o32a_1
XFILLER_115_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10456_ _10456_/A _10492_/B vssd1 vssd1 vccd1 vccd1 _10472_/S sky130_fd_sc_hd__nor2_2
XFILLER_124_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13175_ _17729_/Q _13180_/B vssd1 vssd1 vccd1 vccd1 _13175_/Y sky130_fd_sc_hd__nor2_1
X_10387_ _10387_/A vssd1 vssd1 vccd1 vccd1 _18578_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__04009_ clkbuf_0__04009_/X vssd1 vssd1 vccd1 vccd1 _15854__154/A sky130_fd_sc_hd__clkbuf_16
XFILLER_237_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12126_ _17515_/Q _17736_/Q _12136_/S vssd1 vssd1 vccd1 vccd1 _12127_/B sky130_fd_sc_hd__mux2_1
X_17983_ _18001_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04371_ _16327_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04371_/X sky130_fd_sc_hd__clkbuf_16
X_12057_ _12006_/X _12052_/X _12115_/S vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__mux2_1
X_16934_ _16892_/X _16923_/X _16933_/Y vssd1 vssd1 vccd1 vccd1 _16934_/X sky130_fd_sc_hd__a21o_1
X_11008_ _08991_/X _18274_/Q _11016_/S vssd1 vssd1 vccd1 vccd1 _11009_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16865_ _18149_/Q _18141_/Q _18133_/Q _18277_/Q _16803_/X _16804_/X vssd1 vssd1 vccd1
+ vccd1 _16865_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ _18604_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_1
X_15816_ _18573_/Q _18574_/Q _18575_/Q _18576_/Q _18877_/Q _18878_/Q vssd1 vssd1 vccd1
+ vccd1 _15816_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1__f__03153_ clkbuf_0__03153_/X vssd1 vssd1 vccd1 vccd1 _14305__499/A sky130_fd_sc_hd__clkbuf_16
X_16796_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16797_/A sky130_fd_sc_hd__buf_2
XFILLER_225_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03184_ _14456_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03184_/X sky130_fd_sc_hd__clkbuf_16
X_18535_ _18535_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ _12957_/X _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__and2b_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18466_ _18482_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14320__511 _14320__511/A vssd1 vssd1 vccd1 vccd1 _18146_/CLK sky130_fd_sc_hd__inv_2
X_14629_ _18365_/Q _18317_/Q _18373_/Q _17706_/Q _14599_/X _14600_/X vssd1 vssd1 vccd1
+ vccd1 _14629_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18397_ _18397_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17348_ _17340_/X _17348_/B vssd1 vssd1 vccd1 vccd1 _17349_/A sky130_fd_sc_hd__and2b_1
XFILLER_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03986_ clkbuf_0__03986_/X vssd1 vssd1 vccd1 vccd1 _15778__1059/A sky130_fd_sc_hd__clkbuf_16
XFILLER_147_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17279_ _17279_/A vssd1 vssd1 vccd1 vccd1 _17288_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13112__416 _13115__419/A vssd1 vssd1 vccd1 vccd1 _17712_/CLK sky130_fd_sc_hd__inv_2
XFILLER_162_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14277__476 _14277__476/A vssd1 vssd1 vccd1 vccd1 _18111_/CLK sky130_fd_sc_hd__inv_2
X_19018_ _19027_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_216_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _08983_/A vssd1 vssd1 vccd1 vccd1 _19215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04569_ _16633_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04569_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_229_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _09605_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09535_ _09535_/A vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09466_ _10770_/A _10770_/B _10770_/C vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__nand3b_4
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _09412_/S vssd1 vssd1 vccd1 vccd1 _09406_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03173_ clkbuf_0__03173_/X vssd1 vssd1 vccd1 vccd1 _14403__577/A sky130_fd_sc_hd__clkbuf_16
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15403__904 _15403__904/A vssd1 vssd1 vccd1 vccd1 _18591_/CLK sky130_fd_sc_hd__inv_2
X_10310_ _10310_/A _10372_/A vssd1 vssd1 vccd1 vccd1 _10326_/S sky130_fd_sc_hd__or2_2
XFILLER_192_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ _11290_/A vssd1 vssd1 vccd1 vccd1 _18161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10241_ _10241_/A vssd1 vssd1 vccd1 vccd1 _18640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10172_ _10172_/A vssd1 vssd1 vccd1 vccd1 _18696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14980_ _18455_/Q _14979_/C _18456_/Q vssd1 vssd1 vccd1 vccd1 _14981_/B sky130_fd_sc_hd__a21oi_1
XFILLER_248_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _13943_/B vssd1 vssd1 vccd1 vccd1 _13941_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13862_ _17931_/Q _13850_/X _13861_/X _13857_/X vssd1 vssd1 vccd1 vccd1 _17931_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15601_ _15611_/A _15601_/B _15604_/B vssd1 vssd1 vccd1 vccd1 _15601_/X sky130_fd_sc_hd__or3_1
X_12813_ _17646_/Q _17989_/Q _12822_/S vssd1 vssd1 vccd1 vccd1 _12814_/B sky130_fd_sc_hd__mux2_1
XFILLER_216_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16581_ _19021_/Q _16578_/B _16580_/Y vssd1 vssd1 vccd1 vccd1 _19021_/D sky130_fd_sc_hd__o21a_1
X_13793_ _13792_/X _13778_/A _13789_/X vssd1 vssd1 vccd1 vccd1 _13793_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_203_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18320_ _18320_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15532_ _15535_/C vssd1 vssd1 vccd1 vccd1 _15642_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12746_/B _12742_/A _12734_/X vssd1 vssd1 vccd1 vccd1 _12745_/B sky130_fd_sc_hd__o21ai_1
XFILLER_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18251_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12673_/X _12709_/B _12675_/C vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__and3b_1
XFILLER_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17202_ _17202_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _19242_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ _11626_/A vssd1 vssd1 vccd1 vccd1 _17545_/D sky130_fd_sc_hd__clkbuf_1
X_18182_ _18182_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _19225_/Q _19224_/Q _19223_/Q _17133_/D vssd1 vssd1 vccd1 vccd1 _17149_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11557_ _17707_/Q _10901_/X _11557_/S vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10508_ _10135_/X _18524_/Q _10508_/S vssd1 vssd1 vccd1 vccd1 _10509_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11488_ _11488_/A vssd1 vssd1 vccd1 vccd1 _18050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _16018_/B _16020_/B vssd1 vssd1 vccd1 vccd1 _16015_/Y sky130_fd_sc_hd__nand2_1
X_13227_ input60/X _13650_/A vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__nand2_1
X_10439_ _10454_/S vssd1 vssd1 vccd1 vccd1 _10448_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12109_ _12024_/X _12026_/X _12109_/S vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__mux2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ _17690_/Q _12932_/X _12850_/X _17687_/Q vssd1 vssd1 vccd1 vccd1 _13097_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_17966_ _19039_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16917_ _18119_/Q _18111_/Q _18103_/Q _18095_/Q _16893_/X _16894_/X vssd1 vssd1 vccd1
+ vccd1 _16917_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17897_ _19109_/CLK _17897_/D vssd1 vssd1 vccd1 vccd1 _17897_/Q sky130_fd_sc_hd__dfxtp_1
X_14803__735 _14806__738/A vssd1 vssd1 vccd1 vccd1 _18378_/CLK sky130_fd_sc_hd__inv_2
XFILLER_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16848_ _16844_/X _16847_/X _16875_/S vssd1 vssd1 vccd1 vccd1 _16848_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16779_ _16765_/X _16776_/Y _16778_/Y _14079_/A _16762_/X vssd1 vssd1 vccd1 vccd1
+ _16780_/B sky130_fd_sc_hd__o32a_1
XFILLER_209_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09320_ _09745_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _09336_/S sky130_fd_sc_hd__nor2_2
XFILLER_206_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18518_ _18518_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03167_ _14374_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03167_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _13488_/A _18079_/Q _13540_/A _18078_/Q vssd1 vssd1 vccd1 vccd1 _09252_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_55_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03098_ _14178_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03098_/X sky130_fd_sc_hd__clkbuf_16
X_18449_ _18449_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15465__953 _15648__954/A vssd1 vssd1 vccd1 vccd1 _18640_/CLK sky130_fd_sc_hd__inv_2
X_09182_ _19165_/Q _09112_/X _09184_/S vssd1 vssd1 vccd1 vccd1 _09183_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16314__214 _16314__214/A vssd1 vssd1 vccd1 vccd1 _18930_/CLK sky130_fd_sc_hd__inv_2
XFILLER_239_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03969_ clkbuf_0__03969_/X vssd1 vssd1 vccd1 vccd1 _15691__989/A sky130_fd_sc_hd__clkbuf_16
XFILLER_162_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15852__152 _15854__154/A vssd1 vssd1 vccd1 vccd1 _18827_/CLK sky130_fd_sc_hd__inv_2
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ _08966_/A vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08897_ _19305_/Q _08789_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136__849 _15136__849/A vssd1 vssd1 vccd1 vccd1 _18525_/CLK sky130_fd_sc_hd__inv_2
XFILLER_216_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09518_ _19000_/Q _09495_/X _09518_/S vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__mux2_1
X_10790_ _11565_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _10813_/S sky130_fd_sc_hd__nor2_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09449_/X sky130_fd_sc_hd__or2_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15663__965 _15664__966/A vssd1 vssd1 vccd1 vccd1 _18682_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ _12474_/A vssd1 vssd1 vccd1 vccd1 _12768_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ _11411_/A vssd1 vssd1 vccd1 vccd1 _18111_/D sky130_fd_sc_hd__clkbuf_1
X_12391_ _12386_/X _12390_/X _12448_/A vssd1 vssd1 vccd1 vccd1 _12392_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _13755_/A _14120_/X _14123_/X vssd1 vssd1 vccd1 vccd1 _14130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11342_ _11341_/X _18140_/Q _11345_/S vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19329_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03156_ clkbuf_0__03156_/X vssd1 vssd1 vccd1 vccd1 _14320__511/A sky130_fd_sc_hd__clkbuf_16
XFILLER_180_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ _13783_/X _14055_/X _14060_/X vssd1 vssd1 vccd1 vccd1 _14061_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_181_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11273_ _18664_/Q vssd1 vssd1 vccd1 vccd1 _11273_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_180_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13012_ _17683_/Q _13090_/B vssd1 vssd1 vccd1 vccd1 _13020_/A sky130_fd_sc_hd__xnor2_1
XFILLER_152_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10224_ _18677_/Q _09749_/X _10230_/S vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17820_ _19146_/CLK _17820_/D vssd1 vssd1 vccd1 vccd1 _17820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10155_ _18703_/Q _10072_/X _10155_/S vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__mux2_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ _19327_/CLK _17751_/D vssd1 vssd1 vccd1 vccd1 _17751_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14963_ _14963_/A _14963_/B _14963_/C _14963_/D vssd1 vssd1 vccd1 vccd1 _14964_/D
+ sky130_fd_sc_hd__or4_1
X_10086_ _18730_/Q _10063_/X _10086_/S vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13914_ _13411_/X _13908_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13914_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_0__f__03989_ clkbuf_0__03989_/X vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__clkbuf_16
X_17682_ _17959_/CLK _17682_/D vssd1 vssd1 vccd1 vccd1 _17682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14894_ _15059_/A _16097_/B vssd1 vssd1 vccd1 vccd1 _14894_/Y sky130_fd_sc_hd__nor2_2
XFILLER_235_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16633_/X sky130_fd_sc_hd__buf_1
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _13845_/A _13845_/B vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16564_ _16570_/A vssd1 vssd1 vccd1 vccd1 _16564_/X sky130_fd_sc_hd__clkbuf_2
X_13776_ _17902_/Q _13770_/X _13775_/Y vssd1 vssd1 vccd1 vccd1 _17902_/D sky130_fd_sc_hd__o21a_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10988_ _11204_/B _11347_/B vssd1 vssd1 vccd1 vccd1 _11004_/S sky130_fd_sc_hd__nor2_2
XFILLER_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18303_ _18303_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
X_15515_ _15543_/C _17842_/Q _15515_/S vssd1 vssd1 vccd1 vccd1 _15524_/C sky130_fd_sc_hd__mux2_1
XFILLER_245_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ _12727_/A _12727_/B _12727_/C _12727_/D vssd1 vssd1 vccd1 vccd1 _12737_/D
+ sky130_fd_sc_hd__and4_1
X_19283_ _19288_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
X_16495_ _16493_/X _16494_/Y _16469_/X vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18234_ _18234_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12658_ _12658_/A _12666_/D vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__and2_1
XFILLER_176_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11609_ _17569_/Q _10701_/A _11611_/S vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__mux2_1
X_18165_ _18165_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 _18165_/Q sky130_fd_sc_hd__dfxtp_1
X_15377_ _19219_/Q _19107_/Q _18290_/Q _19099_/Q _15308_/X _09613_/A vssd1 vssd1 vccd1
+ vccd1 _15377_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12589_ _18007_/Q _14067_/B _14065_/B _12840_/A _12775_/B vssd1 vssd1 vccd1 vccd1
+ _12589_/X sky130_fd_sc_hd__a41o_1
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _17117_/A _17117_/C _17117_/B vssd1 vssd1 vccd1 vccd1 _17118_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18096_ _18096_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08820_ _19320_/Q _08792_/X _08822_/S vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _18998_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_19 _11773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ _08807_/A vssd1 vssd1 vccd1 vccd1 _16294_/B sky130_fd_sc_hd__clkbuf_4
X_17949_ _17951_/CLK _17949_/D vssd1 vssd1 vccd1 vccd1 _17949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09303_ _09318_/S vssd1 vssd1 vccd1 vccd1 _09312_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09234_ _09235_/A _18562_/Q _09238_/A vssd1 vssd1 vccd1 vccd1 _09244_/A sky130_fd_sc_hd__o21ai_1
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _09165_/A vssd1 vssd1 vccd1 vccd1 _19173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09096_ _10698_/A vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__buf_2
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14333__521 _14334__522/A vssd1 vssd1 vccd1 vccd1 _18156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ _18765_/Q _09943_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _09679_/A vssd1 vssd1 vccd1 vccd1 _08949_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_218_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _19252_/Q vssd1 vssd1 vccd1 vccd1 _17237_/B sky130_fd_sc_hd__clkbuf_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _18315_/Q _10910_/X _10911_/S vssd1 vssd1 vccd1 vccd1 _10912_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11891_ _11975_/S vssd1 vssd1 vccd1 vccd1 _11936_/S sky130_fd_sc_hd__buf_2
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13630_ _13630_/A vssd1 vssd1 vccd1 vccd1 _17854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10842_ _10842_/A vssd1 vssd1 vccd1 vccd1 _18351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13561_ _13561_/A vssd1 vssd1 vccd1 vccd1 _17831_/D sky130_fd_sc_hd__clkbuf_1
X_10773_ _18378_/Q _10690_/X _10781_/S vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15300_ _18831_/Q _18823_/Q _18815_/Q _18682_/Q _15299_/X _15225_/X vssd1 vssd1 vccd1
+ vccd1 _15300_/X sky130_fd_sc_hd__mux4_2
X_12512_ _12496_/X _12494_/X _12493_/X _12485_/X _12538_/A _12567_/S vssd1 vssd1 vccd1
+ vccd1 _12512_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16280_ _16280_/A _16280_/B vssd1 vssd1 vccd1 vccd1 _16280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13492_ _17809_/Q _13490_/Y _13491_/Y vssd1 vssd1 vccd1 vccd1 _17809_/D sky130_fd_sc_hd__o21a_1
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14494__650 _14496__652/A vssd1 vssd1 vccd1 vccd1 _18285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15231_ _19212_/Q _19100_/Q _18283_/Q _19092_/Q _15230_/X _09631_/X vssd1 vssd1 vccd1
+ vccd1 _15231_/X sky130_fd_sc_hd__mux4_2
X_12443_ _12443_/A vssd1 vssd1 vccd1 vccd1 _12443_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15859__158 _15859__158/A vssd1 vssd1 vccd1 vccd1 _18833_/CLK sky130_fd_sc_hd__inv_2
XFILLER_201_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15162_ _15168_/A vssd1 vssd1 vccd1 vccd1 _15162_/X sky130_fd_sc_hd__buf_1
X_12374_ _17608_/Q _17609_/Q _12435_/A vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14113_ _14113_/A _14113_/B _16052_/C vssd1 vssd1 vccd1 vccd1 _14120_/A sky130_fd_sc_hd__and3_1
XFILLER_154_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11325_ _11325_/A vssd1 vssd1 vccd1 vccd1 _18146_/D sky130_fd_sc_hd__clkbuf_1
X_15093_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__buf_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14044_ _13750_/A _14039_/X _14034_/X vssd1 vssd1 vccd1 vccd1 _14044_/Y sky130_fd_sc_hd__a21oi_1
X_18921_ _18921_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11256_ _11256_/A vssd1 vssd1 vccd1 vccd1 _18172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10207_ _18684_/Q _09752_/X _10211_/S vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11187_ _11202_/S vssd1 vssd1 vccd1 vccd1 _11196_/S sky130_fd_sc_hd__clkbuf_2
X_18852_ _18922_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10138_ _10049_/A _10424_/A _10138_/C vssd1 vssd1 vccd1 vccd1 _10620_/B sky130_fd_sc_hd__nand3b_4
X_17803_ _19133_/CLK _17803_/D vssd1 vssd1 vccd1 vccd1 _17803_/Q sky130_fd_sc_hd__dfxtp_1
X_18783_ _18783_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _18868_/Q vssd1 vssd1 vccd1 vccd1 _16002_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17734_ _19147_/CLK _17734_/D vssd1 vssd1 vccd1 vccd1 _17734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _14940_/A _14944_/X _14945_/X vssd1 vssd1 vccd1 vccd1 _14950_/C sky130_fd_sc_hd__a21bo_1
X_10069_ _10132_/A vssd1 vssd1 vccd1 vccd1 _10069_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17665_ _19016_/CLK _17665_/D vssd1 vssd1 vccd1 vccd1 _17665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14877_ _15086_/A vssd1 vssd1 vccd1 vccd1 _14877_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_101 _11751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_112 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16616_ _19037_/Q _16614_/B _14184_/A vssd1 vssd1 vccd1 vccd1 _16616_/Y sky130_fd_sc_hd__a21oi_1
XINSDIODE2_123 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ _13830_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13829_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17596_ _17602_/CLK _17596_/D vssd1 vssd1 vccd1 vccd1 _17596_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_134 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_145 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_156 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_167 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19335_ _19339_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13759_ _13759_/A _13759_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13855_/B sky130_fd_sc_hd__and3_1
XINSDIODE2_178 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_189 _09879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19266_ _19266_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16478_ _18978_/Q _16482_/C vssd1 vssd1 vccd1 vccd1 _16478_/Y sky130_fd_sc_hd__xnor2_1
X_18217_ _18217_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15429_ _15429_/A vssd1 vssd1 vccd1 vccd1 _15429_/X sky130_fd_sc_hd__buf_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19197_ _19197_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
X_14395__570 _14396__571/A vssd1 vssd1 vccd1 vccd1 _18205_/CLK sky130_fd_sc_hd__inv_2
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18148_ _18148_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03806_ clkbuf_0__03806_/X vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18079_ _18869_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09921_ _09921_/A vssd1 vssd1 vccd1 vccd1 _18789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09852_/A vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_217_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03599_ clkbuf_0__03599_/X vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_219_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _08803_/A vssd1 vssd1 vccd1 vccd1 _19342_/D sky130_fd_sc_hd__clkbuf_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _08880_/X _18838_/Q _09787_/S vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _13520_/B vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__inv_2
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14816__745 _14818__747/A vssd1 vssd1 vccd1 vccd1 _18388_/CLK sky130_fd_sc_hd__inv_2
XFILLER_167_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ _19150_/Q _09108_/X _09221_/S vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09148_ _09476_/A _09148_/B _09148_/C vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__or3_4
XFILLER_135_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ _18994_/Q vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11110_ _18233_/Q _11047_/X _11116_/S vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12090_ _11957_/X _11962_/X _11966_/X _12085_/X _11907_/S _12075_/A vssd1 vssd1 vccd1
+ vccd1 _12090_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ _11041_/A vssd1 vssd1 vccd1 vccd1 _18259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _13066_/A vssd1 vssd1 vccd1 vccd1 _12992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _19155_/Q _18420_/Q _18314_/Q _18298_/Q _14563_/X _14564_/X vssd1 vssd1 vccd1
+ vccd1 _14732_/B sky130_fd_sc_hd__mux4_1
X_11943_ _17777_/Q vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__inv_2
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17450_ _17450_/A vssd1 vssd1 vccd1 vccd1 _19331_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865__162 _15867__164/A vssd1 vssd1 vccd1 vccd1 _18837_/CLK sky130_fd_sc_hd__inv_2
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14660_/X _14661_/X _14662_/S vssd1 vssd1 vccd1 vccd1 _14662_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11874_ _17390_/A vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__buf_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _18973_/Q _16401_/B vssd1 vssd1 vccd1 vccd1 _16417_/A sky130_fd_sc_hd__xnor2_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _13613_/A vssd1 vssd1 vccd1 vccd1 _17848_/D sky130_fd_sc_hd__clkbuf_1
X_17381_ _11888_/X _17381_/B _17381_/C vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__and3b_1
X_10825_ _18358_/Q _10803_/X _10825_/S vssd1 vssd1 vccd1 vccd1 _10826_/A sky130_fd_sc_hd__mux2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14593_ _19173_/Q _19165_/Q _19197_/Q _18332_/Q _14591_/X _14592_/X vssd1 vssd1 vccd1
+ vccd1 _14593_/X sky130_fd_sc_hd__mux4_2
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19120_ _19120_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13544_ _14078_/A _13544_/B vssd1 vssd1 vccd1 vccd1 _17826_/D sky130_fd_sc_hd__nor2_1
XFILLER_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10756_ _18385_/Q _10695_/X _10762_/S vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _19051_/CLK _19051_/D vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16263_ _16171_/A _16262_/X _16162_/S vssd1 vssd1 vccd1 vccd1 _16263_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ _17805_/Q _13477_/B vssd1 vssd1 vccd1 vccd1 _13475_/Y sky130_fd_sc_hd__nor2_1
XFILLER_201_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ _10687_/A vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__clkbuf_1
X_18002_ _18013_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
X_15214_ _15301_/A vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__clkbuf_4
X_12426_ _12672_/B _17610_/Q _12426_/S vssd1 vssd1 vccd1 vccd1 _12426_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17503__1 _17506__4/A vssd1 vssd1 vccd1 vccd1 _19345_/CLK sky130_fd_sc_hd__inv_2
XFILLER_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16194_ _16194_/A vssd1 vssd1 vccd1 vccd1 _16278_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ _12707_/A _17619_/Q _12426_/S vssd1 vssd1 vccd1 vccd1 _12357_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__04571_ clkbuf_0__04571_/X vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11308_ _11308_/A vssd1 vssd1 vccd1 vccd1 _18153_/D sky130_fd_sc_hd__clkbuf_1
X_15076_ _15076_/A _15076_/B vssd1 vssd1 vccd1 vccd1 _15079_/B sky130_fd_sc_hd__and2_1
X_12288_ _12280_/X _12288_/B vssd1 vssd1 vccd1 vccd1 _12289_/A sky130_fd_sc_hd__and2b_1
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14027_ _13733_/A _14017_/X _14020_/X vssd1 vssd1 vccd1 vccd1 _14027_/Y sky130_fd_sc_hd__a21oi_1
X_18904_ _18904_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_1
X_11239_ _11165_/X _18179_/Q _11239_/S vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18835_ _18835_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18766_ _18766_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
X_15978_ _18865_/Q vssd1 vssd1 vccd1 vccd1 _15985_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14929_ _17855_/Q _14942_/B _17854_/Q vssd1 vssd1 vccd1 vccd1 _14930_/B sky130_fd_sc_hd__o21ai_1
X_17717_ _17717_/CLK _17717_/D vssd1 vssd1 vccd1 vccd1 _17717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18697_ _18697_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04005_ clkbuf_0__04005_/X vssd1 vssd1 vccd1 vccd1 _15855_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_223_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17648_ _18012_/CLK _17648_/D vssd1 vssd1 vccd1 vccd1 _17648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17579_ _17579_/CLK _17579_/D vssd1 vssd1 vccd1 vccd1 _17579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19318_ _19318_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19249_ _19251_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09002_ hold25/X vssd1 vssd1 vccd1 vccd1 _11068_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04838_ clkbuf_0__04838_/X vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_247_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__07557_ clkbuf_0__07557_/X vssd1 vssd1 vccd1 vccd1 _12332__394/A sky130_fd_sc_hd__clkbuf_16
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09904_ _09904_/A vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09835_ _09835_/A vssd1 vssd1 vccd1 vccd1 _18816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ _09766_/A vssd1 vssd1 vccd1 vccd1 _18845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14445__611 _14447__613/A vssd1 vssd1 vccd1 vccd1 _18246_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09697_ _09697_/A vssd1 vssd1 vccd1 vccd1 _09697_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04591_ clkbuf_0__04591_/X vssd1 vssd1 vccd1 vccd1 _16728__342/A sky130_fd_sc_hd__clkbuf_16
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10123_/X _18449_/Q _10612_/S vssd1 vssd1 vccd1 vccd1 _10611_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ _11590_/A vssd1 vssd1 vccd1 vccd1 _17578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17395__88 _17395__88/A vssd1 vssd1 vccd1 vccd1 _19301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ _10541_/A vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13260_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13260_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10472_ _18540_/Q _10351_/X _10472_/S vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12211_ _17521_/Q _12202_/X _12204_/X _17522_/Q _12210_/X vssd1 vssd1 vccd1 vccd1
+ _12217_/B sky130_fd_sc_hd__o221ai_1
XFILLER_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13191_ _13368_/A vssd1 vssd1 vccd1 vccd1 _14079_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _12142_/A vssd1 vssd1 vccd1 vccd1 _17519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12073_ _11974_/X _12091_/B _11982_/X _12072_/X _12018_/X _12045_/S vssd1 vssd1 vccd1
+ vccd1 _12073_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16950_ _09859_/A _16949_/X _16886_/X vssd1 vssd1 vccd1 vccd1 _16950_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ _11024_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11040_/S sky130_fd_sc_hd__nor2_2
X_15901_ _17814_/Q _15943_/B vssd1 vssd1 vccd1 vccd1 _15902_/B sky130_fd_sc_hd__xor2_1
X_16881_ _16881_/A vssd1 vssd1 vccd1 vccd1 _16881_/X sky130_fd_sc_hd__buf_2
XFILLER_238_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18620_ _18620_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18551_ _18551_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_1
X_12975_ _13066_/A vssd1 vssd1 vccd1 vccd1 _12975_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03809_ clkbuf_0__03809_/X vssd1 vssd1 vccd1 vccd1 _15648__954/A sky130_fd_sc_hd__clkbuf_16
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _19081_/Q _18345_/Q _17579_/Q _18797_/Q _14568_/X _14569_/X vssd1 vssd1 vccd1
+ vccd1 _14715_/B sky130_fd_sc_hd__mux4_2
X_11926_ _11924_/X _11925_/X _12067_/S vssd1 vssd1 vccd1 vccd1 _11926_/X sky130_fd_sc_hd__mux2_1
X_18482_ _18482_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17433_/A vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14645_ _14664_/A _14644_/X _14619_/X vssd1 vssd1 vccd1 vccd1 _14645_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _13420_/B vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__buf_2
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17364_ _19280_/Q _17478_/B vssd1 vssd1 vccd1 vccd1 _17364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10808_ _10808_/A vssd1 vssd1 vccd1 vccd1 _18365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14576_ _17581_/Q _18379_/Q _18387_/Q _18421_/Q _14574_/X _14575_/X vssd1 vssd1 vccd1
+ vccd1 _14577_/B sky130_fd_sc_hd__mux4_1
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11788_ _18066_/Q _13216_/C vssd1 vssd1 vccd1 vccd1 _13278_/B sky130_fd_sc_hd__or2b_4
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19103_ _19103_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16315_ _16315_/A vssd1 vssd1 vccd1 vccd1 _16315_/X sky130_fd_sc_hd__buf_1
X_13527_ _13951_/A vssd1 vssd1 vccd1 vccd1 _15083_/B sky130_fd_sc_hd__buf_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10739_ _10739_/A vssd1 vssd1 vccd1 vccd1 _18393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19034_ _19037_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16246_ _18748_/Q _18756_/Q _18764_/Q _18772_/Q _16149_/X _16150_/X vssd1 vssd1 vccd1
+ vccd1 _16246_/X sky130_fd_sc_hd__mux4_1
X_13458_ _13165_/X _13444_/B _13457_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _17801_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _18008_/Q vssd1 vssd1 vccd1 vccd1 _12515_/A sky130_fd_sc_hd__inv_2
XFILLER_12_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16177_ _10406_/A _16169_/Y _16171_/Y _16174_/Y _16176_/Y vssd1 vssd1 vccd1 vccd1
+ _16177_/X sky130_fd_sc_hd__o32a_2
Xoutput105 _19389_/X vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_2
X_13389_ _13247_/X _13388_/Y _13337_/X vssd1 vssd1 vccd1 vccd1 _13389_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 _11736_/X vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_2
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput127 _19392_/X vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput138 _19399_/X vssd1 vssd1 vccd1 vccd1 jtag_tdi sky130_fd_sc_hd__buf_2
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput149 _11855_/X vssd1 vssd1 vccd1 vccd1 wb_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15059_ _15059_/A _15060_/B _15059_/C vssd1 vssd1 vccd1 vccd1 _18470_/D sky130_fd_sc_hd__nor3_1
Xclkbuf_0__04585_ _16695_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04585_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _09620_/A _09628_/A vssd1 vssd1 vccd1 vccd1 _09622_/B sky130_fd_sc_hd__or2_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18818_ _18818_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509__663 _14509__663/A vssd1 vssd1 vccd1 vccd1 _18298_/CLK sky130_fd_sc_hd__inv_2
XFILLER_243_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09551_ _09551_/A vssd1 vssd1 vccd1 vccd1 _18956_/D sky130_fd_sc_hd__clkbuf_1
X_18749_ _18749_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03398_ _14753_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03398_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09482_ _09745_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09505_/S sky130_fd_sc_hd__nor2_2
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04019_ _15890_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04019_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17301__77 _17302__78/A vssd1 vssd1 vccd1 vccd1 _19273_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09818_ _09688_/X _18823_/Q _09818_/S vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_55_wb_clk_i clkbuf_leaf_55_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17621_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _18886_/Q vssd1 vssd1 vccd1 vccd1 _09749_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ _12760_/A vssd1 vssd1 vccd1 vccd1 _17635_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04574_ clkbuf_0__04574_/X vssd1 vssd1 vccd1 vccd1 _16663__299/A sky130_fd_sc_hd__clkbuf_16
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/A vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_opt_8_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _17615_/Q _12694_/C _12694_/D vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__and3_1
XFILLER_215_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A vssd1 vssd1 vccd1 vccd1 _17538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _17585_/Q _10898_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput18 io_in[28] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_6
XFILLER_156_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16100_ _16152_/A vssd1 vssd1 vccd1 vccd1 _16276_/A sky130_fd_sc_hd__buf_2
X_13312_ _13184_/X _13311_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _13312_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 vga_r[0] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_8
X_10524_ _18517_/Q _10348_/X _10526_/S vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16031_ _18875_/Q _16031_/B vssd1 vssd1 vccd1 vccd1 _16031_/Y sky130_fd_sc_hd__nor2_1
X_13243_ _17742_/Q _13219_/X _13242_/Y vssd1 vssd1 vccd1 vccd1 _17742_/D sky130_fd_sc_hd__o21a_1
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10455_ _10455_/A vssd1 vssd1 vccd1 vccd1 _18548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13174_ _13212_/B vssd1 vssd1 vccd1 vccd1 _13180_/B sky130_fd_sc_hd__clkbuf_2
X_10386_ _08801_/X _18578_/Q _10388_/S vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__04008_ clkbuf_0__04008_/X vssd1 vssd1 vccd1 vccd1 _15846__147/A sky130_fd_sc_hd__clkbuf_16
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12125_ _12176_/S vssd1 vssd1 vccd1 vccd1 _12136_/S sky130_fd_sc_hd__buf_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17982_ _18001_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04370_ _16321_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04370_/X sky130_fd_sc_hd__clkbuf_16
X_12056_ _11994_/X _12004_/X _12005_/X _12008_/X _12116_/A _12018_/X vssd1 vssd1 vccd1
+ vccd1 _12056_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16933_ _16818_/X _16932_/X _16860_/X vssd1 vssd1 vccd1 vccd1 _16933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11007_ _11022_/S vssd1 vssd1 vccd1 vccd1 _11016_/S sky130_fd_sc_hd__buf_2
XFILLER_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16864_ _18117_/Q _18109_/Q _18101_/Q _18093_/Q _16799_/X _16801_/X vssd1 vssd1 vccd1
+ vccd1 _16864_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18603_ _18603_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03152_ clkbuf_0__03152_/X vssd1 vssd1 vccd1 vccd1 _14297__492/A sky130_fd_sc_hd__clkbuf_16
X_15815_ _18569_/Q _18570_/Q _18571_/Q _18572_/Q _18877_/Q _16044_/A vssd1 vssd1 vccd1
+ vccd1 _15815_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16795_ _16795_/A _16795_/B vssd1 vssd1 vccd1 vccd1 _19136_/D sky130_fd_sc_hd__nor2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14795__729 _14795__729/A vssd1 vssd1 vccd1 vccd1 _18372_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18534_ _18534_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03183_ _14450_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03183_/X sky130_fd_sc_hd__clkbuf_16
X_12958_ _17964_/Q _17673_/Q _13022_/B vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__mux2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17071__57 _17071__57/A vssd1 vssd1 vccd1 vccd1 _19206_/CLK sky130_fd_sc_hd__inv_2
X_11909_ _19240_/Q vssd1 vssd1 vccd1 vccd1 _17194_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18465_ _18465_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12889_ _12877_/X _12889_/B vssd1 vssd1 vccd1 vccd1 _12890_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ _18855_/Q _18349_/Q _19190_/Q _18357_/Q _14637_/A _14627_/X vssd1 vssd1 vccd1
+ vccd1 _14628_/X sky130_fd_sc_hd__mux4_1
X_18396_ _18396_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17347_ _17756_/Q _19287_/Q _17350_/S vssd1 vssd1 vccd1 vccd1 _17348_/B sky130_fd_sc_hd__mux2_1
XFILLER_202_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14559_ _19049_/Q vssd1 vssd1 vccd1 vccd1 _14730_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__03985_ clkbuf_0__03985_/X vssd1 vssd1 vccd1 vccd1 _15771__1053/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _17278_/A vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__clkbuf_1
X_19017_ _19027_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
X_16229_ _16227_/X _16228_/X _16248_/S vssd1 vssd1 vccd1 vccd1 _16229_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08982_ _19215_/Q _08958_/X _08982_/S vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04568_ _16627_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04568_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03419_ clkbuf_0__03419_/X vssd1 vssd1 vccd1 vccd1 _14866__786/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ _15303_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__buf_2
XFILLER_84_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _18963_/Q _09492_/X _09536_/S vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09465_ _10770_/B _09449_/A _09464_/Y vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__o21bai_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09396_ _10967_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09412_/S sky130_fd_sc_hd__or2_2
XFILLER_212_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_102_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18886_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03172_ clkbuf_0__03172_/X vssd1 vssd1 vccd1 vccd1 _14399__574/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _18640_/Q _10175_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10171_ _18696_/Q _10069_/X _10173_/S vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _13441_/X _13925_/X _13929_/Y _13636_/X vssd1 vssd1 vccd1 vccd1 _17953_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ input68/X _13867_/B vssd1 vssd1 vccd1 vccd1 _13861_/X sky130_fd_sc_hd__and2_1
X_15600_ _18654_/Q _15605_/C vssd1 vssd1 vccd1 vccd1 _15604_/B sky130_fd_sc_hd__and2_1
XFILLER_234_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12812_/A vssd1 vssd1 vccd1 vccd1 _12812_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16580_ _16602_/A _16585_/C vssd1 vssd1 vccd1 vccd1 _16580_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13792_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13792_/X sky130_fd_sc_hd__clkbuf_4
X_14382__561 _14382__561/A vssd1 vssd1 vccd1 vccd1 _18196_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15531_ _15481_/Y _15482_/X _15485_/X _15528_/X _15530_/Y vssd1 vssd1 vccd1 vccd1
+ _15535_/C sky130_fd_sc_hd__a2111oi_4
X_12743_ _12746_/B _12746_/C _12746_/D vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__and3_1
XFILLER_231_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18250_ _18250_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12674_ _12672_/B _12673_/A _17610_/Q vssd1 vssd1 vccd1 vccd1 _12675_/C sky130_fd_sc_hd__a21o_1
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _19242_/Q _17195_/X _17164_/X vssd1 vssd1 vccd1 vccd1 _17202_/B sky130_fd_sc_hd__o21ai_1
XFILLER_163_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14458__621 _14461__624/A vssd1 vssd1 vccd1 vccd1 _18256_/CLK sky130_fd_sc_hd__inv_2
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _17545_/Q _09682_/A _11629_/S vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__mux2_1
X_18181_ _18181_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17132_ _17132_/A vssd1 vssd1 vccd1 vccd1 _19224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _11556_/A vssd1 vssd1 vccd1 vccd1 _17708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _10507_/A vssd1 vssd1 vccd1 vccd1 _18525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _14287_/A vssd1 vssd1 vccd1 vccd1 _14275_/X sky130_fd_sc_hd__buf_1
XFILLER_13_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _09139_/X _18050_/Q _11491_/S vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16014_ _16018_/B _16018_/C _16013_/Y vssd1 vssd1 vccd1 vccd1 _16014_/Y sky130_fd_sc_hd__o21ai_1
X_13226_ _17737_/Q _13218_/X _13225_/Y vssd1 vssd1 vccd1 vccd1 _17737_/D sky130_fd_sc_hd__o21a_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10438_ _10638_/B _10492_/B vssd1 vssd1 vccd1 vccd1 _10454_/S sky130_fd_sc_hd__or2_2
XFILLER_124_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13157_ _13428_/A vssd1 vssd1 vccd1 vccd1 _13472_/A sky130_fd_sc_hd__buf_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10369_/A vssd1 vssd1 vccd1 vccd1 _18586_/D sky130_fd_sc_hd__clkbuf_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12108_ _12108_/A vssd1 vssd1 vccd1 vccd1 _12108_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _17687_/Q _12850_/X _12932_/X _17690_/Q vssd1 vssd1 vccd1 vccd1 _13088_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_17965_ _19039_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12039_ _12099_/S _12030_/X _12034_/Y _12038_/Y vssd1 vssd1 vccd1 vccd1 _12207_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_16916_ _19140_/Q _16797_/X _16914_/X _16915_/X vssd1 vssd1 vccd1 vccd1 _19140_/D
+ sky130_fd_sc_hd__o211a_1
X_17896_ _19109_/CLK _17896_/D vssd1 vssd1 vccd1 vccd1 _17896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12237__381 _12239__383/A vssd1 vssd1 vccd1 vccd1 _17545_/CLK sky130_fd_sc_hd__inv_2
XFILLER_226_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16847_ _16845_/X _16846_/X _16984_/A vssd1 vssd1 vccd1 vccd1 _16847_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16778_ _16783_/A _16778_/B vssd1 vssd1 vccd1 vccd1 _16778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _18517_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03166_ _14368_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03166_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_234_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14283__481 _14284__482/A vssd1 vssd1 vccd1 vccd1 _18116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18072_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_233_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09250_ _09250_/A _13520_/B vssd1 vssd1 vccd1 vccd1 _09252_/A sky130_fd_sc_hd__or2_1
XFILLER_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03097_ _14172_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03097_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18448_ _18448_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09181_/A vssd1 vssd1 vccd1 vccd1 _19166_/D sky130_fd_sc_hd__clkbuf_1
X_18379_ _18379_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03968_ clkbuf_0__03968_/X vssd1 vssd1 vccd1 vccd1 _15685__984/A sky130_fd_sc_hd__clkbuf_16
XFILLER_174_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891__180 _15893__182/A vssd1 vssd1 vccd1 vccd1 _18856_/CLK sky130_fd_sc_hd__inv_2
XFILLER_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ _19268_/Q _08964_/X _08968_/S vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08896_ _08896_/A vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09517_ _09517_/A vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _09433_/X _09449_/B _09447_/Y vssd1 vssd1 vccd1 vccd1 _19050_/D sky130_fd_sc_hd__o21a_1
XFILLER_227_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09394_/S vssd1 vssd1 vccd1 vccd1 _09388_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_149_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11410_ _11332_/X _18111_/Q _11412_/S vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12390_ _12388_/X _12389_/X _12390_/S vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ _11341_/A vssd1 vssd1 vccd1 vccd1 _11341_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03155_ clkbuf_0__03155_/X vssd1 vssd1 vccd1 vccd1 _14317__509/A sky130_fd_sc_hd__clkbuf_16
XFILLER_181_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14060_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14060_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11272_ _11272_/A vssd1 vssd1 vccd1 vccd1 _18167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13011_ _17670_/Q _12850_/X _12932_/X _17673_/Q vssd1 vssd1 vccd1 vccd1 _13011_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_238_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10223_ _10223_/A vssd1 vssd1 vccd1 vccd1 _18678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_wb_clk_i _18455_/CLK vssd1 vssd1 vccd1 vccd1 _18462_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14865__785 _14866__786/A vssd1 vssd1 vccd1 vccd1 _18430_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _10154_/A vssd1 vssd1 vccd1 vccd1 _18704_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ _19327_/CLK _17750_/D vssd1 vssd1 vccd1 vccd1 _17750_/Q sky130_fd_sc_hd__dfxtp_1
X_14962_ _14962_/A _14962_/B _14962_/C _14962_/D vssd1 vssd1 vccd1 vccd1 _14963_/D
+ sky130_fd_sc_hd__or4_1
X_10085_ _10085_/A vssd1 vssd1 vccd1 vccd1 _18731_/D sky130_fd_sc_hd__clkbuf_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _16707_/A vssd1 vssd1 vccd1 vccd1 _16701_/X sky130_fd_sc_hd__buf_1
XFILLER_48_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03988_ clkbuf_0__03988_/X vssd1 vssd1 vccd1 vccd1 _16308_/A sky130_fd_sc_hd__clkbuf_16
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13913_ _17947_/Q _13902_/X _13912_/Y vssd1 vssd1 vccd1 vccd1 _17947_/D sky130_fd_sc_hd__o21a_1
X_17681_ _17959_/CLK _17681_/D vssd1 vssd1 vccd1 vccd1 _17681_/Q sky130_fd_sc_hd__dfxtp_1
X_14893_ _09253_/A _15064_/A _14244_/X _13428_/A vssd1 vssd1 vccd1 vccd1 _15059_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ _17925_/Q _13829_/A _13843_/X _13841_/X vssd1 vssd1 vccd1 vccd1 _17925_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16563_ _16567_/A _16715_/B vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__nor2_1
X_13775_ _13285_/X _13771_/X _13774_/X vssd1 vssd1 vccd1 vccd1 _13775_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_245_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ _11383_/A _10987_/B _09025_/A vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__or3b_4
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18302_ _18302_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
X_12726_ _12726_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _17625_/D sky130_fd_sc_hd__nor2_1
XFILLER_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15514_ _18643_/Q _17841_/Q vssd1 vssd1 vccd1 vccd1 _15515_/S sky130_fd_sc_hd__xnor2_1
XFILLER_203_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19282_ _19288_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16494_ _18981_/Q _16499_/B vssd1 vssd1 vccd1 vccd1 _16494_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18233_ _18233_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
X_12657_ _17606_/Q _17605_/Q vssd1 vssd1 vccd1 vccd1 _12666_/D sky130_fd_sc_hd__and2_1
XFILLER_203_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079__194 _16079__194/A vssd1 vssd1 vccd1 vccd1 _18899_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11608_ _11608_/A vssd1 vssd1 vccd1 vccd1 _17570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18164_ _18164_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
X_15376_ _15298_/X _15373_/X _15375_/X _15305_/X vssd1 vssd1 vccd1 vccd1 _15376_/X
+ sky130_fd_sc_hd__o211a_1
X_12588_ _12588_/A _13090_/B vssd1 vssd1 vccd1 vccd1 _12775_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17115_ _17191_/A vssd1 vssd1 vccd1 vccd1 _17289_/A sky130_fd_sc_hd__buf_2
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18095_ _18095_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _08877_/X _17715_/Q _11539_/S vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13209_ _13180_/B _16055_/A _13208_/Y _13187_/X vssd1 vssd1 vccd1 vccd1 _17735_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14189_/A vssd1 vssd1 vccd1 vccd1 _18066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18997_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08728_/X _08749_/X input74/X vssd1 vssd1 vccd1 vccd1 _08807_/A sky130_fd_sc_hd__a21oi_1
X_17948_ _19109_/CLK _17948_/D vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17879_ _18029_/CLK _17879_/D vssd1 vssd1 vccd1 vccd1 _17879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17017__13 _17018__14/A vssd1 vssd1 vccd1 vccd1 _19162_/CLK sky130_fd_sc_hd__inv_2
XFILLER_242_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04167_ clkbuf_0__04167_/X vssd1 vssd1 vccd1 vccd1 _16096__208/A sky130_fd_sc_hd__clkbuf_16
XFILLER_81_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09302_ _09826_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _09318_/S sky130_fd_sc_hd__or2_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03149_ _14281_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03149_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09233_ _18568_/Q _18563_/Q vssd1 vssd1 vccd1 vccd1 _09238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_194_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09164_ _19173_/Q _09112_/X _09166_/S vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _10698_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142__854 _15142__854/A vssd1 vssd1 vccd1 vccd1 _18530_/CLK sky130_fd_sc_hd__inv_2
XFILLER_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ _09997_/A vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _08948_/A vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _08879_/A vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _18987_/Q vssd1 vssd1 vccd1 vccd1 _10910_/X sky130_fd_sc_hd__buf_2
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11890_ _17781_/Q vssd1 vssd1 vccd1 vccd1 _11975_/S sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ _18351_/Q _10800_/X _10843_/S vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__mux2_1
X_13560_ _13560_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__or2_1
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10772_ _10787_/S vssd1 vssd1 vccd1 vccd1 _10781_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _18005_/Q vssd1 vssd1 vccd1 vccd1 _12511_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13491_ _13709_/A _13490_/Y _13408_/X vssd1 vssd1 vccd1 vccd1 _13491_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_240_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15230_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15230_/X sky130_fd_sc_hd__buf_4
X_12442_ _12438_/X _12441_/X _12536_/A vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14112_ _18021_/Q _14092_/X _14111_/Y vssd1 vssd1 vccd1 vccd1 _18021_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11324_ _11321_/X _18146_/Q _11336_/S vssd1 vssd1 vccd1 vccd1 _11325_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _15447_/A vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__buf_1
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14043_ _17995_/Q _14032_/X _14042_/Y vssd1 vssd1 vccd1 vccd1 _17995_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18920_ _18921_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_1
X_11255_ _11162_/X _18172_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11256_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10206_ _10206_/A vssd1 vssd1 vccd1 vccd1 _18685_/D sky130_fd_sc_hd__clkbuf_1
X_18851_ _18851_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11260_/A hold18/X vssd1 vssd1 vccd1 vccd1 _11202_/S sky130_fd_sc_hd__nor2_2
XFILLER_192_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17802_ _19135_/CLK _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10137_ _10137_/A vssd1 vssd1 vccd1 vccd1 _18711_/D sky130_fd_sc_hd__clkbuf_1
X_18782_ _18782_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _15992_/X _15993_/Y _15982_/X vssd1 vssd1 vccd1 vccd1 _18867_/D sky130_fd_sc_hd__a21oi_1
XFILLER_95_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _19147_/CLK _17733_/D vssd1 vssd1 vccd1 vccd1 _17733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14945_ _14940_/A _14944_/X _18454_/Q vssd1 vssd1 vccd1 vccd1 _14945_/X sky130_fd_sc_hd__mux2_1
X_10068_ _10068_/A vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17664_ _18010_/CLK _17664_/D vssd1 vssd1 vccd1 vccd1 _17664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_102 _19385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16615_ _19036_/Q _16613_/B _16614_/Y vssd1 vssd1 vccd1 vccd1 _19036_/D sky130_fd_sc_hd__o21a_1
XINSDIODE2_113 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13827_ _17919_/Q _13820_/Y _13825_/X _13826_/X vssd1 vssd1 vccd1 vccd1 _17919_/D
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_124 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17595_ _17602_/CLK _17595_/D vssd1 vssd1 vccd1 vccd1 _17595_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_135 _17720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_146 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19334_ _19336_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_157 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14503__658 _14503__658/A vssd1 vssd1 vccd1 vccd1 _18293_/CLK sky130_fd_sc_hd__inv_2
X_13758_ _17897_/Q _13743_/B _13757_/Y _13753_/X vssd1 vssd1 vccd1 vccd1 _17897_/D
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_168 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_179 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ _12717_/D _12709_/B _12709_/C vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__and3b_1
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19265_ _19266_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13689_ _13689_/A vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16477_ _16474_/X _16476_/Y _16469_/X vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__a21oi_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18216_ _18216_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
X_19196_ _19196_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18147_ _18147_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
X_15359_ _15298_/X _15356_/X _15358_/X _15305_/X vssd1 vssd1 vccd1 vccd1 _15359_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__03805_ clkbuf_0__03805_/X vssd1 vssd1 vccd1 vccd1 _15754_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18078_ _18869_/CLK _18078_/D vssd1 vssd1 vccd1 vccd1 _18078_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _18789_/Q _09262_/X _09926_/S vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _16871_/A vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03598_ clkbuf_0__03598_/X vssd1 vssd1 vccd1 vccd1 _15153__863/A sky130_fd_sc_hd__clkbuf_16
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _19342_/Q _08801_/X _08805_/S vssd1 vssd1 vccd1 vccd1 _08803_/A sky130_fd_sc_hd__mux2_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A vssd1 vssd1 vccd1 vccd1 _18839_/D sky130_fd_sc_hd__clkbuf_1
X_16541__253 _16541__253/A vssd1 vssd1 vccd1 vccd1 _18999_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08733_ _18080_/Q _18081_/Q _13386_/B _13386_/C vssd1 vssd1 vccd1 vccd1 _13520_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404__578 _14405__579/A vssd1 vssd1 vccd1 vccd1 _18213_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ _09216_/A vssd1 vssd1 vccd1 vccd1 _19151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ _09147_/A vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14296__491 _14297__492/A vssd1 vssd1 vccd1 vccd1 _18126_/CLK sky130_fd_sc_hd__inv_2
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _09078_/A vssd1 vssd1 vccd1 vccd1 _19196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11040_ _18259_/Q _09145_/X _11040_/S vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A vssd1 vssd1 vccd1 vccd1 _17682_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ _12116_/A vssd1 vssd1 vccd1 vccd1 _12016_/S sky130_fd_sc_hd__buf_2
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14730_ _14726_/X _14729_/X _14730_/S vssd1 vssd1 vccd1 vccd1 _14730_/X sky130_fd_sc_hd__mux2_2
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _18856_/Q _18350_/Q _19191_/Q _18358_/Q _14575_/A _09443_/A vssd1 vssd1 vccd1
+ vccd1 _14661_/X sky130_fd_sc_hd__mux4_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _11873_/A vssd1 vssd1 vccd1 vccd1 _11873_/X sky130_fd_sc_hd__buf_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13629_/A _13612_/B vssd1 vssd1 vccd1 vccd1 _13613_/A sky130_fd_sc_hd__or2_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _17803_/Q _16413_/A vssd1 vssd1 vccd1 vccd1 _16401_/B sky130_fd_sc_hd__xnor2_1
X_10824_ _10824_/A vssd1 vssd1 vccd1 vccd1 _18359_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17380_ _17363_/X _17369_/Y _17379_/X _19291_/Q vssd1 vssd1 vccd1 vccd1 _17381_/C
+ sky130_fd_sc_hd__a31o_1
X_14592_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__buf_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13543_ _11742_/B _13425_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13544_/B sky130_fd_sc_hd__mux2_1
X_10755_ _10755_/A vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _18451_/Q _19089_/Q _19126_/Q _18435_/Q _16106_/X _16108_/X vssd1 vssd1 vccd1
+ vccd1 _16262_/X sky130_fd_sc_hd__mux4_2
X_19050_ _19050_/CLK _19050_/D vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfxtp_1
X_13474_ _14079_/A vssd1 vssd1 vccd1 vccd1 _16058_/A sky130_fd_sc_hd__buf_8
XFILLER_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ _18414_/Q _09738_/X _10688_/S vssd1 vssd1 vccd1 vccd1 _10687_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18001_ _18001_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15213_ _19112_/Q _18943_/Q _18601_/Q _19341_/Q _15209_/X _15212_/X vssd1 vssd1 vccd1
+ vccd1 _15213_/X sky130_fd_sc_hd__mux4_1
X_12425_ _17609_/Q vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16193_ _16257_/A _16193_/B vssd1 vssd1 vccd1 vccd1 _16193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12356_ _12435_/A vssd1 vssd1 vccd1 vccd1 _12426_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__04570_ clkbuf_0__04570_/X vssd1 vssd1 vccd1 vccd1 _16644__284/A sky130_fd_sc_hd__clkbuf_16
XFILLER_154_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11147_/X _18153_/Q _11313_/S vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15075_ _14965_/A _16097_/A _15074_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _15075_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12287_ _17561_/Q _18016_/Q _12287_/S vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__mux2_1
XFILLER_84_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15676__976 _15677__977/A vssd1 vssd1 vccd1 vccd1 _18693_/CLK sky130_fd_sc_hd__inv_2
X_14026_ _17989_/Q _14012_/X _14025_/Y vssd1 vssd1 vccd1 vccd1 _17989_/D sky130_fd_sc_hd__o21a_1
X_18903_ _18903_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_1
X_11238_ _11238_/A vssd1 vssd1 vccd1 vccd1 _18180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18834_ _18834_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ _11184_/S vssd1 vssd1 vccd1 vccd1 _11178_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18765_ _18765_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _15974_/X _15976_/Y _16033_/A vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__a21oi_1
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17716_ _17716_/CLK _17716_/D vssd1 vssd1 vccd1 vccd1 _17716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14928_ _18458_/Q _14928_/B vssd1 vssd1 vccd1 vccd1 _14961_/B sky130_fd_sc_hd__xnor2_1
XFILLER_224_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18696_ _18696_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04004_ clkbuf_0__04004_/X vssd1 vssd1 vccd1 vccd1 _15829__134/A sky130_fd_sc_hd__clkbuf_16
X_17647_ _18012_/CLK _17647_/D vssd1 vssd1 vccd1 vccd1 _17647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14878__795 _14882__799/A vssd1 vssd1 vccd1 vccd1 _18440_/CLK sky130_fd_sc_hd__inv_2
XFILLER_247_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _17578_/CLK _17578_/D vssd1 vssd1 vccd1 vccd1 _17578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19317_ _19317_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
X_16529_ _16529_/A vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19248_ _19248_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09001_ _18810_/Q vssd1 vssd1 vccd1 vccd1 _09001_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19179_ _19179_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__04837_ clkbuf_0__04837_/X vssd1 vssd1 vccd1 vccd1 _17011__359/A sky130_fd_sc_hd__clkbuf_16
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__07556_ clkbuf_0__07556_/X vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__clkbuf_16
X_16727__341 _16730__344/A vssd1 vssd1 vccd1 vccd1 _19120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09903_ _18796_/Q _09726_/X _09907_/S vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09834_ _09685_/X _18816_/Q _09836_/S vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09765_ _18845_/Q _09764_/X _09768_/S vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14822__750 _14824__752/A vssd1 vssd1 vccd1 vccd1 _18393_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _09696_/A vssd1 vssd1 vccd1 vccd1 _18899_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04590_ clkbuf_0__04590_/X vssd1 vssd1 vccd1 vccd1 _16724__339/A sky130_fd_sc_hd__clkbuf_16
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _18510_/Q _10345_/X _10544_/S vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ _10471_/A vssd1 vssd1 vccd1 vccd1 _18541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12210_ _17519_/Q _12206_/X _12199_/A _17526_/Q _12209_/Y vssd1 vssd1 vccd1 vccd1
+ _12210_/X sky130_fd_sc_hd__o221a_1
X_14452__616 _14455__619/A vssd1 vssd1 vccd1 vccd1 _18251_/CLK sky130_fd_sc_hd__inv_2
X_13190_ input68/X _13483_/B vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12141_ _12132_/X _12141_/B vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__and2b_1
X_16548__259 _16548__259/A vssd1 vssd1 vccd1 vccd1 _19005_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _19223_/Q _17129_/A _19225_/Q _17142_/B _11980_/X _11981_/X vssd1 vssd1 vccd1
+ vccd1 _12072_/X sky130_fd_sc_hd__mux4_2
XFILLER_173_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15900_ _17817_/Q _17816_/Q _17815_/Q _15937_/B vssd1 vssd1 vccd1 vccd1 _15943_/B
+ sky130_fd_sc_hd__or4_2
X_11023_ _11023_/A vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16880_ _16927_/A _16880_/B vssd1 vssd1 vccd1 vccd1 _16880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _15855_/A vssd1 vssd1 vccd1 vccd1 _15831_/X sky130_fd_sc_hd__buf_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _18550_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
X_12974_ _17303_/A vssd1 vssd1 vccd1 vccd1 _13066_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346__532 _14347__533/A vssd1 vssd1 vccd1 vccd1 _18167_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03808_ clkbuf_0__03808_/X vssd1 vssd1 vccd1 vccd1 _15457__946/A sky130_fd_sc_hd__clkbuf_16
X_15194__880 _15195__881/A vssd1 vssd1 vccd1 vccd1 _18559_/CLK sky130_fd_sc_hd__inv_2
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17083__66 _17083__66/A vssd1 vssd1 vccd1 vccd1 _19215_/CLK sky130_fd_sc_hd__inv_2
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713_ _14732_/A _14713_/B vssd1 vssd1 vccd1 vccd1 _14713_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ _19236_/Q _19237_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__mux2_1
X_18481_ _18482_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15693_/X sky130_fd_sc_hd__buf_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231__376 _12234__379/A vssd1 vssd1 vccd1 vccd1 _17540_/CLK sky130_fd_sc_hd__inv_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17356_/X _17432_/B vssd1 vssd1 vccd1 vccd1 _17433_/A sky130_fd_sc_hd__and2b_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _19147_/Q vssd1 vssd1 vccd1 vccd1 _13820_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14644_ _14607_/X _14634_/Y _14636_/Y _14639_/Y _14643_/Y vssd1 vssd1 vccd1 vccd1
+ _14644_/X sky130_fd_sc_hd__o32a_1
XFILLER_221_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16635__276 _16635__276/A vssd1 vssd1 vccd1 vccd1 _19050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_246_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10807_ _18365_/Q _10806_/X _10813_/S vssd1 vssd1 vccd1 vccd1 _10808_/A sky130_fd_sc_hd__mux2_1
X_17363_ _19281_/Q _12202_/X _12204_/X _19282_/Q _17362_/X vssd1 vssd1 vccd1 vccd1
+ _17363_/X sky130_fd_sc_hd__o221a_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14575_ _14575_/A vssd1 vssd1 vccd1 vccd1 _14575_/X sky130_fd_sc_hd__buf_4
X_11787_ _13873_/A _11787_/B _11826_/A vssd1 vssd1 vccd1 vccd1 _13216_/C sky130_fd_sc_hd__and3_1
XFILLER_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19102_ _19102_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13526_ _13681_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13526_/X sky130_fd_sc_hd__or2_1
X_10738_ _18393_/Q _10695_/X _10744_/S vssd1 vssd1 vccd1 vccd1 _10739_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033_ _19037_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16245_ _16191_/X _16238_/Y _16240_/Y _16242_/Y _16244_/Y vssd1 vssd1 vccd1 vccd1
+ _16245_/X sky130_fd_sc_hd__o32a_2
X_13457_ _17801_/Q _13457_/B vssd1 vssd1 vccd1 vccd1 _13457_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10669_ _10669_/A vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__clkbuf_1
X_12408_ _12408_/A vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ _13769_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13388_/Y sky130_fd_sc_hd__nor2_1
X_16176_ _16143_/X _16175_/X _16119_/X vssd1 vssd1 vccd1 vccd1 _16176_/Y sky130_fd_sc_hd__o21ai_1
Xoutput106 _11771_/X vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_2
XFILLER_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput117 _11732_/X vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_2
XFILLER_142_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput128 _19393_/X vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_2
X_12339_ _13103_/A vssd1 vssd1 vccd1 vccd1 _12339_/X sky130_fd_sc_hd__buf_1
XFILLER_115_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput139 _19400_/X vssd1 vssd1 vccd1 vccd1 jtag_tms sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15058_ _14965_/A _15076_/A _14965_/B _15055_/Y vssd1 vssd1 vccd1 vccd1 _15059_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_141_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _17983_/Q _13989_/X _14008_/Y vssd1 vssd1 vccd1 vccd1 _17983_/D sky130_fd_sc_hd__o21a_1
XFILLER_141_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18817_ _18817_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09550_ _08921_/X _18956_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09551_/A sky130_fd_sc_hd__mux2_1
X_18748_ _18748_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03397_ _14747_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03397_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_110_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09481_ _18887_/Q vssd1 vssd1 vccd1 vccd1 _09481_/X sky130_fd_sc_hd__buf_4
X_18679_ _18679_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14516__668 _14517__669/A vssd1 vssd1 vccd1 vccd1 _18303_/CLK sky130_fd_sc_hd__inv_2
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15098__818 _15099__819/A vssd1 vssd1 vccd1 vccd1 _18494_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ _09817_/A vssd1 vssd1 vccd1 vccd1 _18824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09748_ _09748_/A vssd1 vssd1 vccd1 vccd1 _18851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A vssd1 vssd1 vccd1 vccd1 _09679_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04573_ clkbuf_0__04573_/X vssd1 vssd1 vccd1 vccd1 _16655__292/A sky130_fd_sc_hd__clkbuf_16
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _17927_/Q _11714_/B vssd1 vssd1 vccd1 vccd1 _11711_/A sky130_fd_sc_hd__and2_4
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12690_ _12690_/A vssd1 vssd1 vccd1 vccd1 _17614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _17923_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16554__263 _16555__264/A vssd1 vssd1 vccd1 vccd1 _19009_/CLK sky130_fd_sc_hd__inv_2
X_11641_ _08786_/X _17538_/Q _11647_/S vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__mux2_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _11572_/A vssd1 vssd1 vccd1 vccd1 _17586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13311_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 io_in[29] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_6
XFILLER_183_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10523_ _10523_/A vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13242_ _13240_/X _13232_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _13242_/Y sky130_fd_sc_hd__a21oi_1
X_16030_ _18875_/Q _16031_/B vssd1 vssd1 vccd1 vccd1 _16035_/C sky130_fd_sc_hd__and2_1
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10454_ _10135_/X _18548_/Q _10454_/S vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16073__189 _16073__189/A vssd1 vssd1 vccd1 vccd1 _18894_/CLK sky130_fd_sc_hd__inv_2
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13173_ _14072_/A vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__buf_6
X_10385_ _10385_/A vssd1 vssd1 vccd1 vccd1 _18579_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__04007_ clkbuf_0__04007_/X vssd1 vssd1 vccd1 vccd1 _15842__144/A sky130_fd_sc_hd__clkbuf_16
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12124_ _17770_/Q _17423_/B vssd1 vssd1 vccd1 vccd1 _12176_/S sky130_fd_sc_hd__nand2_2
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14829__756 _14829__756/A vssd1 vssd1 vccd1 vccd1 _18399_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17981_ _18001_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12055_ _12053_/X _12054_/X _12069_/A vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__mux2_2
X_16932_ _16819_/X _16925_/Y _16927_/Y _16929_/Y _16931_/Y vssd1 vssd1 vccd1 vccd1
+ _16932_/X sky130_fd_sc_hd__o32a_1
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _11024_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11022_/S sky130_fd_sc_hd__or2_2
X_16863_ _19138_/Q _16797_/X _16862_/X _15628_/X vssd1 vssd1 vccd1 vccd1 _19138_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_238_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18602_ _18602_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03151_ clkbuf_0__03151_/X vssd1 vssd1 vccd1 vccd1 _14318_/A sky130_fd_sc_hd__clkbuf_16
X_15814_ _18878_/Q vssd1 vssd1 vccd1 vccd1 _16044_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_237_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794_ _13853_/A _16762_/A _16793_/Y _16687_/B vssd1 vssd1 vccd1 vccd1 _16795_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03182_ _14449_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03182_/X sky130_fd_sc_hd__clkbuf_16
X_18533_ _18533_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12957_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07559_ clkbuf_0__07559_/X vssd1 vssd1 vccd1 vccd1 _12342__402/A sky130_fd_sc_hd__clkbuf_16
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11908_ _19238_/Q _19239_/Q _11924_/S vssd1 vssd1 vccd1 vccd1 _11908_/X sky130_fd_sc_hd__mux2_1
X_18464_ _18465_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _17976_/Q _17660_/Q _12891_/S vssd1 vssd1 vccd1 vccd1 _12889_/B sky130_fd_sc_hd__mux2_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17415_ _17415_/A vssd1 vssd1 vccd1 vccd1 _17415_/X sky130_fd_sc_hd__buf_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14627_ _14627_/A vssd1 vssd1 vccd1 vccd1 _14627_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ _11839_/A vssd1 vssd1 vccd1 vccd1 _11839_/X sky130_fd_sc_hd__clkbuf_2
X_18395_ _18395_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17346_ _17346_/A vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14558_ _14555_/X _14557_/X _14729_/S vssd1 vssd1 vccd1 vccd1 _14558_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03984_ clkbuf_0__03984_/X vssd1 vssd1 vccd1 vccd1 _15763__1046/A sky130_fd_sc_hd__clkbuf_16
XFILLER_202_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13509_ _13509_/A vssd1 vssd1 vccd1 vccd1 _17814_/D sky130_fd_sc_hd__clkbuf_1
X_17277_ _17284_/C _17277_/B _17277_/C vssd1 vssd1 vccd1 vccd1 _17278_/A sky130_fd_sc_hd__and3b_1
XFILLER_158_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15878__173 _15878__173/A vssd1 vssd1 vccd1 vccd1 _18848_/CLK sky130_fd_sc_hd__inv_2
XFILLER_220_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19016_ _19016_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
X_16228_ _18715_/Q _18723_/Q _18731_/Q _18496_/Q _16205_/X _16206_/X vssd1 vssd1 vccd1
+ vccd1 _16228_/X sky130_fd_sc_hd__mux4_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _18776_/Q _18634_/Q _18784_/Q _18618_/Q _16158_/X _16138_/A vssd1 vssd1 vccd1
+ vccd1 _16159_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08981_ _08981_/A vssd1 vssd1 vccd1 vccd1 _19216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03418_ clkbuf_0__03418_/X vssd1 vssd1 vccd1 vccd1 _14863__784/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _18932_/Q vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_244_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09533_ _09533_/A vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09464_ _10770_/C _09467_/B _09449_/A vssd1 vssd1 vccd1 vccd1 _09464_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09395_ _09395_/A vssd1 vssd1 vccd1 vccd1 _19067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03171_ clkbuf_0__03171_/X vssd1 vssd1 vccd1 vccd1 _14393__569/A sky130_fd_sc_hd__clkbuf_16
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10170_ _10170_/A vssd1 vssd1 vccd1 vccd1 _18697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _17930_/Q _13850_/X _13859_/X _13857_/X vssd1 vssd1 vccd1 vccd1 _17930_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ _12811_/A vssd1 vssd1 vccd1 vccd1 _17645_/D sky130_fd_sc_hd__clkbuf_1
X_13791_ _17907_/Q _13771_/X _13790_/Y vssd1 vssd1 vccd1 vccd1 _17907_/D sky130_fd_sc_hd__o21a_1
XFILLER_43_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15530_ _18657_/Q _15530_/B vssd1 vssd1 vccd1 vccd1 _15530_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12742_ _12742_/A _12742_/B vssd1 vssd1 vccd1 vccd1 _17630_/D sky130_fd_sc_hd__nor2_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ _12673_/A _12680_/D vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__and2_1
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _15655_/A vssd1 vssd1 vccd1 vccd1 _15461_/X sky130_fd_sc_hd__buf_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _19242_/Q _17203_/C _17203_/D vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__and3_1
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11624_/A vssd1 vssd1 vccd1 vccd1 _17546_/D sky130_fd_sc_hd__clkbuf_1
X_14412_ _14412_/A vssd1 vssd1 vccd1 vccd1 _14412_/X sky130_fd_sc_hd__buf_1
X_18180_ _18180_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
X_15392_ _15410_/A vssd1 vssd1 vccd1 vccd1 _15392_/X sky130_fd_sc_hd__buf_1
XFILLER_168_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17131_ _17135_/B _17131_/B _17277_/B vssd1 vssd1 vccd1 vccd1 _17132_/A sky130_fd_sc_hd__and3b_1
XFILLER_211_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11555_ _17708_/Q _10898_/X _11557_/S vssd1 vssd1 vccd1 vccd1 _11556_/A sky130_fd_sc_hd__mux2_1
X_14343_ _14349_/A vssd1 vssd1 vccd1 vccd1 _14343_/X sky130_fd_sc_hd__buf_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _10132_/X _18525_/Q _10508_/S vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__mux2_1
X_17062_ _17062_/A vssd1 vssd1 vccd1 vccd1 _17062_/X sky130_fd_sc_hd__buf_1
X_11486_ _11486_/A vssd1 vssd1 vccd1 vccd1 _18051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13225_ _13219_/X _13717_/A _13224_/X vssd1 vssd1 vccd1 vccd1 _13225_/Y sky130_fd_sc_hd__a21oi_1
X_16013_ _16018_/B _16018_/C _15963_/X vssd1 vssd1 vccd1 vccd1 _16013_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_195_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10437_ _18563_/Q _10437_/B _10075_/B vssd1 vssd1 vccd1 vccd1 _10492_/B sky130_fd_sc_hd__or3b_4
XFILLER_48_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13156_ _17726_/Q _14134_/B vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _18586_/Q _09738_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12102_/Y _12103_/Y _12104_/Y _12106_/Y _12016_/S _12099_/S vssd1 vssd1 vccd1
+ vccd1 _12189_/A sky130_fd_sc_hd__mux4_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13087_ _13087_/A _13087_/B _13087_/C _13087_/D vssd1 vssd1 vccd1 vccd1 _13087_/X
+ sky130_fd_sc_hd__and4_1
X_17964_ _19037_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10299_ _10299_/A vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12038_ _12016_/S _12037_/X _12020_/A vssd1 vssd1 vccd1 vccd1 _12038_/Y sky130_fd_sc_hd__a21oi_1
X_16915_ _16915_/A vssd1 vssd1 vccd1 vccd1 _16915_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17895_ _19109_/CLK _17895_/D vssd1 vssd1 vccd1 vccd1 _17895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16846_ _19205_/Q _19157_/Q _18268_/Q _18260_/Q _16828_/A _16813_/X vssd1 vssd1 vccd1
+ vccd1 _16846_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ _19134_/Q _19132_/Q _16787_/S vssd1 vssd1 vccd1 vccd1 _16778_/B sky130_fd_sc_hd__mux2_1
XFILLER_241_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13989_ _13995_/A vssd1 vssd1 vccd1 vccd1 _13989_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03165_ _14362_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03165_/X sky130_fd_sc_hd__clkbuf_16
X_18516_ _18516_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03096_ _14166_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03096_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18447_ _18447_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ _19166_/Q _09108_/X _09184_/S vssd1 vssd1 vccd1 vccd1 _09181_/A sky130_fd_sc_hd__mux2_1
X_18378_ _18378_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ _17329_/A vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__clkbuf_1
X_14359__542 _14361__544/A vssd1 vssd1 vccd1 vccd1 _18177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03967_ clkbuf_0__03967_/X vssd1 vssd1 vccd1 vccd1 _15677__977/A sky130_fd_sc_hd__clkbuf_16
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16648__286 _16649__287/A vssd1 vssd1 vccd1 vccd1 _19060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739__1027 _15741__1029/A vssd1 vssd1 vccd1 vccd1 _18744_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17412__102 _17412__102/A vssd1 vssd1 vccd1 vccd1 _19315_/CLK sky130_fd_sc_hd__inv_2
X_08964_ _09694_/A vssd1 vssd1 vccd1 vccd1 _08964_/X sky130_fd_sc_hd__buf_2
XFILLER_248_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08895_ _19306_/Q _08786_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _08896_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__07169_ clkbuf_0__07169_/X vssd1 vssd1 vccd1 vccd1 _17506__4/A sky130_fd_sc_hd__clkbuf_16
XFILLER_204_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ _19001_/Q _09492_/X _09518_/S vssd1 vssd1 vccd1 vccd1 _09517_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09433_/X _09449_/B _09449_/A vssd1 vssd1 vccd1 vccd1 _09447_/Y sky130_fd_sc_hd__a21oi_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09378_ _09508_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09394_/S sky130_fd_sc_hd__nor2_2
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11340_ _11340_/A vssd1 vssd1 vccd1 vccd1 _18141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03154_ clkbuf_0__03154_/X vssd1 vssd1 vccd1 vccd1 _14310__503/A sky130_fd_sc_hd__clkbuf_16
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _18167_/Q _11270_/X _11274_/S vssd1 vssd1 vccd1 vccd1 _11272_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13010_ _13010_/A _13010_/B _13010_/C _13010_/D vssd1 vssd1 vccd1 vccd1 _13010_/X
+ sky130_fd_sc_hd__and4_1
X_10222_ _18678_/Q _09744_/X _10230_/S vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10153_ _18704_/Q _10069_/X _10155_/S vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__mux2_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14961_ _14961_/A _14961_/B _14961_/C _14961_/D vssd1 vssd1 vccd1 vccd1 _14962_/D
+ sky130_fd_sc_hd__or4_1
X_10084_ _18731_/Q _10060_/X _10086_/S vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03987_ clkbuf_0__03987_/X vssd1 vssd1 vccd1 vccd1 _15784__1064/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13912_ _13407_/X _13908_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13912_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ _17963_/CLK _17680_/D vssd1 vssd1 vccd1 vccd1 _17680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ input56/X _13847_/B vssd1 vssd1 vccd1 vccd1 _13843_/X sky130_fd_sc_hd__and2_1
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15829__134 _15829__134/A vssd1 vssd1 vccd1 vccd1 _18809_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16562_ _19015_/Q vssd1 vssd1 vccd1 vccd1 _16567_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13774_ _13880_/A vssd1 vssd1 vccd1 vccd1 _13774_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10986_ _11511_/A vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_216_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18301_ _18301_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15513_ _18642_/Q vssd1 vssd1 vccd1 vccd1 _15543_/C sky130_fd_sc_hd__clkbuf_2
X_12725_ _12727_/B _12723_/A _12718_/X vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__o21ai_1
X_19281_ _19281_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
X_14163__442 _14165__444/A vssd1 vssd1 vccd1 vccd1 _18050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_188_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _16498_/A _16493_/B _16497_/B vssd1 vssd1 vccd1 vccd1 _16493_/X sky130_fd_sc_hd__or3_1
XFILLER_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18232_ _18232_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12656_ _12387_/X _12658_/A _12655_/Y vssd1 vssd1 vccd1 vccd1 _17605_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _17570_/Q _10698_/A _11611_/S vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__mux2_1
X_18163_ _18163_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 _18163_/Q sky130_fd_sc_hd__dfxtp_1
X_12587_ _12587_/A vssd1 vssd1 vccd1 vccd1 _13090_/B sky130_fd_sc_hd__buf_4
X_15375_ _15375_/A _15303_/X vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__or2b_1
XFILLER_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17114_ _17114_/A vssd1 vssd1 vccd1 vccd1 _17191_/A sky130_fd_sc_hd__clkbuf_2
X_18094_ _18094_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
X_11538_ _11538_/A vssd1 vssd1 vccd1 vccd1 _17716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11469_ _11338_/X _18058_/Q _11473_/S vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13208_ _17735_/Q _13208_/B vssd1 vssd1 vccd1 vccd1 _13208_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14188_ _18066_/Q input46/X _14196_/S vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__mux2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13139_ input59/X _13210_/B vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__nand2_4
XFILLER_48_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16721__336 _16724__339/A vssd1 vssd1 vccd1 vccd1 _19115_/CLK sky130_fd_sc_hd__inv_2
X_18996_ _18996_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17947_ _19109_/CLK _17947_/D vssd1 vssd1 vccd1 vccd1 _17947_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17878_ _17878_/CLK _17878_/D vssd1 vssd1 vccd1 vccd1 _17878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16829_ _18203_/Q _18123_/Q _19180_/Q _18251_/Q _16827_/X _16828_/X vssd1 vssd1 vccd1
+ vccd1 _16830_/B sky130_fd_sc_hd__mux4_1
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04166_ clkbuf_0__04166_/X vssd1 vssd1 vccd1 vccd1 _16090__203/A sky130_fd_sc_hd__clkbuf_16
XFILLER_242_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09301_ _10372_/A vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__03148_ _14275_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03148_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _18567_/Q vssd1 vssd1 vccd1 vccd1 _09235_/A sky130_fd_sc_hd__inv_2
XFILLER_210_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09163_ _09163_/A vssd1 vssd1 vccd1 vccd1 _19174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09094_ _09094_/A vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09996_ _18766_/Q _09935_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__mux2_1
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _19274_/Q _08944_/X _08959_/S vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ _19311_/Q _08877_/X _08878_/S vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__mux2_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10840_ _10840_/A vssd1 vssd1 vccd1 vccd1 _18352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10771_ _11601_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _10787_/S sky130_fd_sc_hd__nor2_2
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340__527 _14342__529/A vssd1 vssd1 vccd1 vccd1 _18162_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12510_ _13093_/B _12510_/B _12510_/C _12920_/A vssd1 vssd1 vccd1 vccd1 _12510_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_197_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13490_ _13761_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13490_/Y sky130_fd_sc_hd__nor2_2
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12441_ _12439_/X _12440_/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12372_ _12360_/X _12369_/X _12448_/A vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17419__108 _17419__108/A vssd1 vssd1 vccd1 vccd1 _19321_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14111_ _13792_/X _14099_/A _14108_/X vssd1 vssd1 vccd1 vccd1 _14111_/Y sky130_fd_sc_hd__a21oi_1
X_11323_ _11345_/S vssd1 vssd1 vccd1 vccd1 _11336_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_165_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14042_ _13748_/A _14039_/X _14034_/X vssd1 vssd1 vccd1 vccd1 _14042_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11254_ _11254_/A vssd1 vssd1 vccd1 vccd1 _18173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10205_ _18685_/Q _09749_/X _10211_/S vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18850_ _18850_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11185_ _11185_/A vssd1 vssd1 vccd1 vccd1 _18203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17801_ _19135_/CLK _17801_/D vssd1 vssd1 vccd1 vccd1 _17801_/Q sky130_fd_sc_hd__dfxtp_1
X_10136_ _10135_/X _18711_/Q _10136_/S vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18781_ _18781_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _18867_/Q _15993_/B vssd1 vssd1 vccd1 vccd1 _15993_/Y sky130_fd_sc_hd__nand2_1
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _19147_/CLK _17732_/D vssd1 vssd1 vccd1 vccd1 _17732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14944_ _18455_/Q _17858_/Q vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__xor2_1
X_10067_ _18737_/Q _10066_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__mux2_1
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17663_ _18010_/CLK _17663_/D vssd1 vssd1 vccd1 vccd1 _17663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15119__835 _15122__838/A vssd1 vssd1 vccd1 vccd1 _18511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_103 _19394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16614_ _16620_/A _16614_/B vssd1 vssd1 vccd1 vccd1 _16614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13826_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_114 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17594_ _19016_/CLK _17594_/D vssd1 vssd1 vccd1 vccd1 _17594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_125 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_136 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_147 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19333_ _19337_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
X_15738__1026 _15741__1029/A vssd1 vssd1 vccd1 vccd1 _18743_/CLK sky130_fd_sc_hd__inv_2
XFILLER_232_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13757_ _13815_/A _13757_/B vssd1 vssd1 vccd1 vccd1 _13757_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_158 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10969_ _18290_/Q _09744_/X _10977_/S vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_169 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12708_ _12706_/B _12703_/A _12706_/A vssd1 vssd1 vccd1 vccd1 _12709_/C sky130_fd_sc_hd__a21o_1
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19264_ _19266_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
X_16476_ _18977_/Q _16499_/B vssd1 vssd1 vccd1 vccd1 _16476_/Y sky130_fd_sc_hd__nand2_1
X_13688_ _13688_/A vssd1 vssd1 vccd1 vccd1 _13688_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18215_ _18215_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12639_ _12638_/A _12634_/X _12617_/X vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__o21ai_1
XFILLER_176_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19195_ _19195_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__04853_ clkbuf_0__04853_/X vssd1 vssd1 vccd1 vccd1 _17296__73/A sky130_fd_sc_hd__clkbuf_16
X_15085__809 _15085__809/A vssd1 vssd1 vccd1 vccd1 _18485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18146_ _18146_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03804_ clkbuf_0__03804_/X vssd1 vssd1 vccd1 vccd1 _15446__939/A sky130_fd_sc_hd__clkbuf_16
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _15358_/A _15303_/X vssd1 vssd1 vccd1 vccd1 _15358_/X sky130_fd_sc_hd__or2b_1
XFILLER_184_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18077_ _19146_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15289_ _15244_/X _15276_/X _15288_/X _15267_/X vssd1 vssd1 vccd1 vccd1 _15289_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_160_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _18808_/Q vssd1 vssd1 vccd1 vccd1 _16871_/A sky130_fd_sc_hd__buf_2
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03597_ clkbuf_0__03597_/X vssd1 vssd1 vccd1 vccd1 _15148__859/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _18881_/Q vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__clkbuf_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _08877_/X _18839_/Q _09781_/S vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__mux2_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18979_ _18987_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08732_ _18082_/Q _18083_/Q vssd1 vssd1 vccd1 vccd1 _13386_/C sky130_fd_sc_hd__or2_2
XFILLER_22_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09215_ _19151_/Q _09104_/X _09215_/S vssd1 vssd1 vccd1 vccd1 _09216_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09146_ _19180_/Q _09145_/X _09146_/S vssd1 vssd1 vccd1 vccd1 _09147_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _19196_/Q _08886_/X _09077_/S vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ _09979_/A vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12990_ _12975_/X _12990_/B vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__and2b_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11941_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _18366_/Q _18318_/Q _18374_/Q _17707_/Q _14575_/A _09443_/A vssd1 vssd1 vccd1
+ vccd1 _14660_/X sky130_fd_sc_hd__mux4_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _14922_/B _13446_/X _13611_/S vssd1 vssd1 vccd1 vccd1 _13612_/B sky130_fd_sc_hd__mux2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10823_ _18359_/Q _10800_/X _10825_/S vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14591_ _14594_/A vssd1 vssd1 vccd1 vccd1 _14591_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13542_ _13705_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__nor2_1
XFILLER_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _18386_/Q _10690_/X _10762_/S vssd1 vssd1 vccd1 vccd1 _10755_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14305__499 _14305__499/A vssd1 vssd1 vccd1 vccd1 _18134_/CLK sky130_fd_sc_hd__inv_2
X_16261_ _16280_/A _16261_/B vssd1 vssd1 vccd1 vccd1 _16261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10685_ _10685_/A vssd1 vssd1 vccd1 vccd1 _18415_/D sky130_fd_sc_hd__clkbuf_1
X_13473_ _16059_/A _13463_/B _13471_/Y _13472_/X vssd1 vssd1 vccd1 vccd1 _17804_/D
+ sky130_fd_sc_hd__a211oi_1
X_18000_ _18013_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15212_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15212_/X sky130_fd_sc_hd__clkbuf_4
X_12424_ _12418_/X _12421_/X _12765_/S vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16192_ _18527_/Q _18535_/Q _18543_/Q _18551_/Q _10404_/A _16102_/X vssd1 vssd1 vccd1
+ vccd1 _16193_/B sky130_fd_sc_hd__mux4_1
XFILLER_51_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _15149_/A vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__buf_1
X_12355_ _18012_/Q vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__03620_ _15199_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03620_/X sky130_fd_sc_hd__clkbuf_16
X_11306_ _11306_/A vssd1 vssd1 vccd1 vccd1 _18154_/D sky130_fd_sc_hd__clkbuf_1
X_12286_ _12286_/A vssd1 vssd1 vccd1 vccd1 _17560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15074_ _18472_/Q _18470_/Q _15074_/C vssd1 vssd1 vccd1 vccd1 _15074_/X sky130_fd_sc_hd__and3_1
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15872__168 _15872__168/A vssd1 vssd1 vccd1 vccd1 _18843_/CLK sky130_fd_sc_hd__inv_2
X_14025_ _13786_/X _14017_/X _14020_/X vssd1 vssd1 vccd1 vccd1 _14025_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11237_ _11162_/X _18180_/Q _11239_/S vssd1 vssd1 vccd1 vccd1 _11238_/A sky130_fd_sc_hd__mux2_1
X_18902_ _18902_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11168_ _11223_/A _11365_/A vssd1 vssd1 vccd1 vccd1 _11184_/S sky130_fd_sc_hd__or2_2
X_18833_ _18833_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10119_ _10119_/A vssd1 vssd1 vccd1 vccd1 _18717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18764_ _18764_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ _11099_/A vssd1 vssd1 vccd1 vccd1 _18238_/D sky130_fd_sc_hd__clkbuf_1
X_15976_ _18864_/Q _15993_/B vssd1 vssd1 vccd1 vccd1 _15976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _17715_/CLK _17715_/D vssd1 vssd1 vccd1 vccd1 _17715_/Q sky130_fd_sc_hd__dfxtp_1
X_14927_ _17855_/Q _14942_/B vssd1 vssd1 vccd1 vccd1 _14928_/B sky130_fd_sc_hd__xor2_1
XFILLER_212_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18695_ _18695_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _18012_/CLK _17646_/D vssd1 vssd1 vccd1 vccd1 _17646_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__05083_ _17421_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05083_/X sky130_fd_sc_hd__clkbuf_16
X_14858_ _14864_/A vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__buf_1
XFILLER_91_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ _17913_/Q _13796_/X _13808_/Y vssd1 vssd1 vccd1 vccd1 _17913_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17577_ _17577_/CLK _17577_/D vssd1 vssd1 vccd1 vccd1 _17577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19316_ _19316_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16528_ input69/X _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16529_/A sky130_fd_sc_hd__and3_1
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19247_ _19247_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16459_ _16467_/A _16459_/B _16466_/C vssd1 vssd1 vccd1 vccd1 _16459_/X sky130_fd_sc_hd__or3_1
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ _18808_/Q hold26/A vssd1 vssd1 vccd1 vccd1 _09856_/B sky130_fd_sc_hd__xnor2_1
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19178_ _19178_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__04836_ clkbuf_0__04836_/X vssd1 vssd1 vccd1 vccd1 _17002__351/A sky130_fd_sc_hd__clkbuf_16
XFILLER_192_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18129_ _18129_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__07555_ clkbuf_0__07555_/X vssd1 vssd1 vccd1 vccd1 _12322__386/A sky130_fd_sc_hd__clkbuf_16
XFILLER_247_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09902_ _09902_/A vssd1 vssd1 vccd1 vccd1 _18797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09833_ _09833_/A vssd1 vssd1 vccd1 vccd1 _18817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ _18881_/Q vssd1 vssd1 vccd1 vccd1 _09764_/X sky130_fd_sc_hd__buf_2
XFILLER_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14410__583 _14410__583/A vssd1 vssd1 vccd1 vccd1 _18218_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09695_ _09694_/X _18899_/Q _09698_/S vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144__429 _14144__429/A vssd1 vssd1 vccd1 vccd1 _18037_/CLK sky130_fd_sc_hd__inv_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15722__1014 _15722__1014/A vssd1 vssd1 vccd1 vccd1 _18731_/CLK sky130_fd_sc_hd__inv_2
X_10470_ _18541_/Q _10348_/X _10472_/S vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ _09129_/A vssd1 vssd1 vccd1 vccd1 _19186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _17519_/Q _17732_/Q _12153_/S vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__mux2_1
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _19226_/Q vssd1 vssd1 vccd1 vccd1 _17142_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15737__1025 _15737__1025/A vssd1 vssd1 vccd1 vccd1 _18742_/CLK sky130_fd_sc_hd__inv_2
XFILLER_173_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _09055_/X _18267_/Q _11022_/S vssd1 vssd1 vccd1 vccd1 _11023_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _16308_/A vssd1 vssd1 vccd1 vccd1 _15830_/X sky130_fd_sc_hd__buf_1
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _15767_/A vssd1 vssd1 vccd1 vccd1 _15761_/X sky130_fd_sc_hd__buf_1
X_12973_ _12973_/A vssd1 vssd1 vccd1 vccd1 _17677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03807_ clkbuf_0__03807_/X vssd1 vssd1 vccd1 vccd1 _15454__944/A sky130_fd_sc_hd__clkbuf_16
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _19154_/Q _18419_/Q _18313_/Q _18297_/Q _14563_/X _14564_/X vssd1 vssd1 vccd1
+ vccd1 _14713_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11924_ _19234_/Q _19235_/Q _11924_/S vssd1 vssd1 vccd1 vccd1 _11924_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _15785_/A _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15754_/A vssd1 vssd1 vccd1 vccd1 _15692_/X sky130_fd_sc_hd__buf_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17431_ _17750_/Q _19326_/Q _17497_/B vssd1 vssd1 vccd1 vccd1 _17432_/B sky130_fd_sc_hd__mux2_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14643_ _14640_/X _14642_/X _14561_/X vssd1 vssd1 vccd1 vccd1 _14643_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11855_/A vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17362_ _19279_/Q _12206_/X _12199_/X _19286_/Q _17361_/Y vssd1 vssd1 vccd1 vccd1
+ _17362_/X sky130_fd_sc_hd__o221a_1
X_10806_ _18989_/Q vssd1 vssd1 vccd1 vccd1 _10806_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14574_ _14627_/A vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11786_ _11786_/A vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_201_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19101_ _19101_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15682__981 _15682__981/A vssd1 vssd1 vccd1 vccd1 _18698_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _17819_/Q _13522_/X _13524_/Y vssd1 vssd1 vccd1 vccd1 _17819_/D sky130_fd_sc_hd__o21a_1
X_17293_ _17291_/Y _17289_/C _17292_/X _17109_/A _17109_/B vssd1 vssd1 vccd1 vccd1
+ _19266_/D sky130_fd_sc_hd__o2111a_1
X_10737_ _10737_/A vssd1 vssd1 vccd1 vccd1 _18394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19032_ _19040_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16244_ _16143_/X _16243_/X _16162_/S vssd1 vssd1 vccd1 vccd1 _16244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13456_ _13161_/X _13444_/B _13455_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _17800_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10668_ _18422_/Q _09738_/X _10670_/S vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _12407_/A vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__clkbuf_2
X_16175_ _18447_/Q _19085_/Q _19122_/Q _18431_/Q _16144_/X _10420_/X vssd1 vssd1 vccd1
+ vccd1 _16175_/X sky130_fd_sc_hd__mux4_2
XFILLER_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13387_ _14069_/B _13387_/B vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__or2_1
X_10599_ _10599_/A vssd1 vssd1 vccd1 vccd1 _18485_/D sky130_fd_sc_hd__clkbuf_1
Xoutput107 _11767_/X vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_2
XFILLER_217_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput118 _11728_/X vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_2
XFILLER_154_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput129 _19394_/X vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__buf_2
XFILLER_182_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15057_ _15057_/A _15057_/B vssd1 vssd1 vccd1 vccd1 _15060_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12269_ _12269_/A vssd1 vssd1 vccd1 vccd1 _17555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14008_ _13815_/X _13995_/A _14005_/X vssd1 vssd1 vccd1 vccd1 _14008_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15203__888 _15203__888/A vssd1 vssd1 vccd1 vccd1 _18567_/CLK sky130_fd_sc_hd__inv_2
XFILLER_229_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18816_ _18816_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18747_ _18747_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03396_ _14746_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03396_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15959_ _15962_/A vssd1 vssd1 vccd1 vccd1 _16035_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18678_ _18678_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_1
X_09480_ _09480_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _19041_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17629_ _17629_/CLK _17629_/D vssd1 vssd1 vccd1 vccd1 _17629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09816_ _09685_/X _18824_/Q _09818_/S vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09747_ _18851_/Q _09744_/X _09759_/S vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09678_/A vssd1 vssd1 vccd1 vccd1 _18905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__04572_ clkbuf_0__04572_/X vssd1 vssd1 vccd1 vccd1 _16651__289/A sky130_fd_sc_hd__clkbuf_16
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A vssd1 vssd1 vccd1 vccd1 _17539_/D sky130_fd_sc_hd__clkbuf_1
X_15823__129 _15823__129/A vssd1 vssd1 vccd1 vccd1 _18804_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11571_ _17586_/Q _10895_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13310_ _17762_/Q _13303_/X _13309_/Y vssd1 vssd1 vccd1 vccd1 _17762_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_64_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _17703_/CLK sky130_fd_sc_hd__clkbuf_16
X_10522_ _18518_/Q _10345_/X _10526_/S vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13241_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__clkbuf_2
X_10453_ _10453_/A vssd1 vssd1 vccd1 vccd1 _18549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13172_ input71/X _13650_/A vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__nand2_4
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10384_ _08798_/X _18579_/Q _10388_/S vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__04006_ clkbuf_0__04006_/X vssd1 vssd1 vccd1 vccd1 _15836__139/A sky130_fd_sc_hd__clkbuf_16
XFILLER_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14417__589 _14417__589/A vssd1 vssd1 vccd1 vccd1 _18224_/CLK sky130_fd_sc_hd__inv_2
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12123_ _17490_/B _12123_/B _12123_/C _12122_/X vssd1 vssd1 vccd1 vccd1 _17423_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_237_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17980_ _18001_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12054_ _11994_/X _11996_/X _12004_/X _12005_/X _12076_/S _12045_/S vssd1 vssd1 vccd1
+ vccd1 _12054_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16931_ _09859_/A _16930_/X _16886_/X vssd1 vssd1 vccd1 vccd1 _16931_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11005_ _11005_/A vssd1 vssd1 vccd1 vccd1 _18275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16862_ _09845_/X _16848_/X _16861_/Y vssd1 vssd1 vccd1 vccd1 _16862_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16641__281 _16644__284/A vssd1 vssd1 vccd1 vccd1 _19055_/CLK sky130_fd_sc_hd__inv_2
XFILLER_238_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18601_ _18601_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15813_ _18879_/Q vssd1 vssd1 vccd1 vccd1 _15813_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03150_ clkbuf_0__03150_/X vssd1 vssd1 vccd1 vccd1 _14292__489/A sky130_fd_sc_hd__clkbuf_16
X_16793_ _19136_/Q _16771_/B _16792_/X vssd1 vssd1 vccd1 vccd1 _16793_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04839_ clkbuf_0__04839_/X vssd1 vssd1 vccd1 vccd1 _17016__12/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18532_ _18532_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03181_ _14443_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03181_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_206_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12956_ _12956_/A vssd1 vssd1 vccd1 vccd1 _17672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__07558_ clkbuf_0__07558_/X vssd1 vssd1 vccd1 vccd1 _12335__396/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _11898_/X _11903_/X _11907_/S vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18463_ _19039_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12887_/A vssd1 vssd1 vccd1 vccd1 _17659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14624_/X _14625_/X _14688_/S vssd1 vssd1 vccd1 vccd1 _14626_/X sky130_fd_sc_hd__mux2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _17925_/Q _13326_/B _11836_/Y _13830_/A _11837_/Y vssd1 vssd1 vccd1 vccd1
+ _11838_/X sky130_fd_sc_hd__o2111a_2
X_18394_ _18394_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17345_ _17340_/X _17345_/B vssd1 vssd1 vccd1 vccd1 _17346_/A sky130_fd_sc_hd__and2b_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14557_ _18853_/Q _18347_/Q _19188_/Q _18355_/Q _14575_/A _14554_/X vssd1 vssd1 vccd1
+ vccd1 _14557_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11769_ _11769_/A vssd1 vssd1 vccd1 vccd1 _11769_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03983_ clkbuf_0__03983_/X vssd1 vssd1 vccd1 vccd1 _15760__1044/A sky130_fd_sc_hd__clkbuf_16
XFILLER_159_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _13560_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__or2_1
X_17276_ _17276_/A _17276_/B vssd1 vssd1 vccd1 vccd1 _17277_/C sky130_fd_sc_hd__or2_1
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19015_ _19016_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16227_ _18747_/Q _18755_/Q _18763_/Q _18771_/Q _16127_/X _16128_/X vssd1 vssd1 vccd1
+ vccd1 _16227_/X sky130_fd_sc_hd__mux4_1
X_13439_ _17794_/Q _13444_/B vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16158_ _18565_/Q vssd1 vssd1 vccd1 vccd1 _16158_/X sky130_fd_sc_hd__buf_2
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _19216_/Q _08955_/X _08982_/S vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03417_ clkbuf_0__03417_/X vssd1 vssd1 vccd1 vccd1 _14853__775/A sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09601_ _18933_/Q vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15721__1013 _15722__1014/A vssd1 vssd1 vccd1 vccd1 _18730_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09532_ _18964_/Q _09489_/X _09536_/S vssd1 vssd1 vccd1 vccd1 _09533_/A sky130_fd_sc_hd__mux2_1
X_15689__987 _15689__987/A vssd1 vssd1 vccd1 vccd1 _18704_/CLK sky130_fd_sc_hd__inv_2
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ _09476_/A _09480_/A vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__and2_2
XFILLER_58_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14522__673 _14523__674/A vssd1 vssd1 vccd1 vccd1 _18308_/CLK sky130_fd_sc_hd__inv_2
X_09394_ _19067_/Q _08967_/X _09394_/S vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03170_ clkbuf_0__03170_/X vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325__389 _12325__389/A vssd1 vssd1 vccd1 vccd1 _17570_/CLK sky130_fd_sc_hd__inv_2
XFILLER_153_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12810_ _12795_/X _12810_/B vssd1 vssd1 vccd1 vccd1 _12811_/A sky130_fd_sc_hd__and2b_1
X_13790_ _13244_/X _13778_/X _13789_/X vssd1 vssd1 vccd1 vccd1 _13790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12741_ _12746_/C _12746_/D _12734_/X vssd1 vssd1 vccd1 vccd1 _12742_/B sky130_fd_sc_hd__o21ai_1
XFILLER_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _17610_/Q _12672_/B vssd1 vssd1 vccd1 vccd1 _12680_/D sky130_fd_sc_hd__and2_1
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423__593 _14423__593/A vssd1 vssd1 vccd1 vccd1 _18228_/CLK sky130_fd_sc_hd__inv_2
XFILLER_231_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _17546_/Q _09679_/A _11629_/S vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14835__761 _14835__761/A vssd1 vssd1 vccd1 vccd1 _18404_/CLK sky130_fd_sc_hd__inv_2
X_17130_ _17129_/B _17129_/C _17129_/A vssd1 vssd1 vccd1 vccd1 _17131_/B sky130_fd_sc_hd__a21o_1
XFILLER_168_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11554_ _11554_/A vssd1 vssd1 vccd1 vccd1 _17709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10505_ _10505_/A vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__clkbuf_1
X_11485_ _09136_/X _18051_/Q _11485_/S vssd1 vssd1 vccd1 vccd1 _11486_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16012_ _18871_/Q vssd1 vssd1 vccd1 vccd1 _16018_/B sky130_fd_sc_hd__clkbuf_1
X_13224_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10436_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13155_ _13786_/A vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__buf_6
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10367_ _10367_/A vssd1 vssd1 vccd1 vccd1 _18587_/D sky130_fd_sc_hd__clkbuf_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12106_ _12106_/A vssd1 vssd1 vccd1 vccd1 _12106_/Y sky130_fd_sc_hd__clkinv_2
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13086_ _17694_/Q _12921_/X _12838_/X _17702_/Q _13085_/X vssd1 vssd1 vccd1 vccd1
+ _13087_/D sky130_fd_sc_hd__a221oi_1
X_17963_ _17963_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _18614_/Q _10183_/X _10302_/S vssd1 vssd1 vccd1 vccd1 _10299_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12037_ _12035_/X _12036_/X _12037_/S vssd1 vssd1 vccd1 vccd1 _12037_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16914_ _16892_/X _16903_/X _16913_/Y vssd1 vssd1 vccd1 vccd1 _16914_/X sky130_fd_sc_hd__a21o_1
XFILLER_238_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17894_ _19109_/CLK _17894_/D vssd1 vssd1 vccd1 vccd1 _17894_/Q sky130_fd_sc_hd__dfxtp_1
X_14465__627 _14467__629/A vssd1 vssd1 vccd1 vccd1 _18262_/CLK sky130_fd_sc_hd__inv_2
XFILLER_239_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17029__23 _17030__24/A vssd1 vssd1 vccd1 vccd1 _19172_/CLK sky130_fd_sc_hd__inv_2
XFILLER_226_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16845_ _18057_/Q _18049_/Q _18041_/Q _18033_/Q _16809_/X _16810_/X vssd1 vssd1 vccd1
+ vccd1 _16845_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16776_ _19133_/Q _16786_/B vssd1 vssd1 vccd1 vccd1 _16776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_230_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13988_ _13995_/A vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18515_ _18515_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03164_ _14356_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03164_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_248_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12939_ _17658_/Q _13095_/B vssd1 vssd1 vccd1 vccd1 _12941_/C sky130_fd_sc_hd__xnor2_1
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03095_ _14160_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03095_/X sky130_fd_sc_hd__clkbuf_16
X_18446_ _18446_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ _14736_/A _14609_/B vssd1 vssd1 vccd1 vccd1 _14609_/Y sky130_fd_sc_hd__nor2_1
X_18377_ _18377_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
X_15589_ _18652_/Q vssd1 vssd1 vccd1 vccd1 _15595_/B sky130_fd_sc_hd__clkbuf_1
X_17328_ _17323_/X _17328_/B vssd1 vssd1 vccd1 vccd1 _17329_/A sky130_fd_sc_hd__and2b_1
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03966_ clkbuf_0__03966_/X vssd1 vssd1 vccd1 vccd1 _15673__974/A sky130_fd_sc_hd__clkbuf_16
XFILLER_239_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17259_ _17262_/C _17258_/C _17262_/B vssd1 vssd1 vccd1 vccd1 _17260_/C sky130_fd_sc_hd__a21o_1
XFILLER_175_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15695__991 _15696__992/A vssd1 vssd1 vccd1 vccd1 _18708_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14290__487 _14290__487/A vssd1 vssd1 vccd1 vccd1 _18122_/CLK sky130_fd_sc_hd__inv_2
X_08963_ _08963_/A vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08894_ _08894_/A vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__07168_ clkbuf_0__07168_/X vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09515_ _09515_/A vssd1 vssd1 vccd1 vccd1 _19002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12331__393 _12332__394/A vssd1 vssd1 vccd1 vccd1 _17574_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09446_/A _09453_/B vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__nor2_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ _09377_/A _09639_/A _09789_/A vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__or3b_4
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_4_1_wb_clk_i clkbuf_opt_4_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _11873_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03153_ clkbuf_0__03153_/X vssd1 vssd1 vccd1 vccd1 _14302__496/A sky130_fd_sc_hd__clkbuf_16
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11270_ _18665_/Q vssd1 vssd1 vccd1 vccd1 _11270_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10221_ hold3/A vssd1 vssd1 vccd1 vccd1 _10230_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_234_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10152_ _10152_/A vssd1 vssd1 vccd1 vccd1 _18705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ _14960_/A _14960_/B _14960_/C vssd1 vssd1 vccd1 vccd1 _14964_/C sky130_fd_sc_hd__or3_1
X_10083_ _10083_/A vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _17946_/Q _13902_/X _13910_/Y vssd1 vssd1 vccd1 vccd1 _17946_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f__03986_ clkbuf_0__03986_/X vssd1 vssd1 vccd1 vccd1 _15776__1057/A sky130_fd_sc_hd__clkbuf_16
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529__679 _14529__679/A vssd1 vssd1 vccd1 vccd1 _18314_/CLK sky130_fd_sc_hd__inv_2
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13842_ _17924_/Q _13829_/X _13840_/X _13841_/X vssd1 vssd1 vccd1 vccd1 _17924_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16561_ _13430_/Y _09084_/C _11816_/X _16530_/B vssd1 vssd1 vccd1 vccd1 _19014_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_244_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13773_ _17901_/Q _13770_/X _13772_/Y vssd1 vssd1 vccd1 vccd1 _17901_/D sky130_fd_sc_hd__o21a_1
XFILLER_245_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10985_ _15808_/B _10985_/B vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__nand2_8
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15512_ _18646_/Q _15512_/B vssd1 vssd1 vccd1 vccd1 _15524_/B sky130_fd_sc_hd__xnor2_1
X_18300_ _18300_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _12727_/B _12727_/C _12727_/D vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__and3_1
X_19280_ _19281_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16492_ _18981_/Q _18980_/Q _16492_/C vssd1 vssd1 vccd1 vccd1 _16497_/B sky130_fd_sc_hd__and3_1
XFILLER_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18231_ _18231_/CLK _18231_/D vssd1 vssd1 vccd1 vccd1 _18231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ _12387_/X _12658_/A _12755_/A vssd1 vssd1 vccd1 vccd1 _12655_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_231_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11606_ _11606_/A vssd1 vssd1 vccd1 vccd1 _17571_/D sky130_fd_sc_hd__clkbuf_1
X_18162_ _18162_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15374_ _18678_/Q _18584_/Q _17539_/Q _17514_/Q _15308_/A _15301_/X vssd1 vssd1 vccd1
+ vccd1 _15375_/A sky130_fd_sc_hd__mux4_1
X_12586_ _12584_/X _12585_/X _12586_/S vssd1 vssd1 vccd1 vccd1 _12587_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17113_ _17113_/A vssd1 vssd1 vccd1 vccd1 _19220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14325_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14325_/X sky130_fd_sc_hd__buf_1
XFILLER_102_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11537_ _08874_/X _17716_/Q _11539_/S vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__mux2_1
X_18093_ _18093_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15720__1012 _15720__1012/A vssd1 vssd1 vccd1 vccd1 _18729_/CLK sky130_fd_sc_hd__inv_2
X_17044_ _17068_/A vssd1 vssd1 vccd1 vccd1 _17044_/X sky130_fd_sc_hd__buf_1
XFILLER_116_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14256_ _14256_/A vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__buf_1
X_11468_ _11468_/A vssd1 vssd1 vccd1 vccd1 _18059_/D sky130_fd_sc_hd__clkbuf_1
X_15836__139 _15836__139/A vssd1 vssd1 vccd1 vccd1 _18814_/CLK sky130_fd_sc_hd__inv_2
X_13207_ _13755_/A vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__buf_12
XFILLER_125_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10419_ _16182_/A vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14187_ _14231_/A vssd1 vssd1 vccd1 vccd1 _14196_/S sky130_fd_sc_hd__clkbuf_2
X_11399_ _11399_/A vssd1 vssd1 vccd1 vccd1 _18116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13138_ _13446_/B vssd1 vssd1 vccd1 vccd1 _13210_/B sky130_fd_sc_hd__clkbuf_4
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _18996_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13069_ _13069_/A vssd1 vssd1 vccd1 vccd1 _17699_/D sky130_fd_sc_hd__clkbuf_1
X_17946_ _19109_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17877_ _17878_/CLK _17877_/D vssd1 vssd1 vccd1 vccd1 _17877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16828_ _16828_/A vssd1 vssd1 vccd1 vccd1 _16828_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__04165_ clkbuf_0__04165_/X vssd1 vssd1 vccd1 vccd1 _16081__195/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16759_ _16788_/A vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ _09300_/A vssd1 vssd1 vccd1 vccd1 _19112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03147_ _14269_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03147_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16654__291 _16655__292/A vssd1 vssd1 vccd1 vccd1 _19065_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09231_ _18561_/Q _18560_/Q _18559_/Q vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__and3_1
XFILLER_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18429_ _18429_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09162_ _19174_/Q _09108_/X _09166_/S vssd1 vssd1 vccd1 vccd1 _09163_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09093_ _19194_/Q _09092_/X _09105_/S vssd1 vssd1 vccd1 vccd1 _09094_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09995_ _10010_/S vssd1 vssd1 vccd1 vccd1 _10004_/S sky130_fd_sc_hd__buf_2
XFILLER_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _08968_/S vssd1 vssd1 vccd1 vccd1 _08959_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _18990_/Q vssd1 vssd1 vccd1 vccd1 _08877_/X sky130_fd_sc_hd__buf_6
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023__18 _17024__19/A vssd1 vssd1 vccd1 vccd1 _19167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_241_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _10770_/A _10770_/B _10770_/C vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__nand3_4
XFILLER_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09429_ _09429_/A vssd1 vssd1 vccd1 vccd1 _19052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ _17607_/Q _17608_/Q _12440_/S vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12371_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12448_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ _18020_/Q _14092_/X _14109_/Y vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__o21a_1
XFILLER_176_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _11475_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11345_/S sky130_fd_sc_hd__or2_2
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _17994_/Q _14032_/X _14040_/Y vssd1 vssd1 vccd1 vccd1 _17994_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11253_ _11159_/X _18173_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11254_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _10204_/A vssd1 vssd1 vccd1 vccd1 _18686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _11165_/X _18203_/Q _11184_/S vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17800_ _19135_/CLK _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Q sky130_fd_sc_hd__dfxtp_1
X_10135_ _10135_/A vssd1 vssd1 vccd1 vccd1 _10135_/X sky130_fd_sc_hd__clkbuf_4
X_18780_ _18780_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_1
X_15992_ _16024_/A _15992_/B _16002_/C vssd1 vssd1 vccd1 vccd1 _15992_/X sky130_fd_sc_hd__or3_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338__399 _12338__399/A vssd1 vssd1 vccd1 vccd1 _17580_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14943_ _14942_/B _14942_/C _18457_/Q vssd1 vssd1 vccd1 vccd1 _14950_/B sky130_fd_sc_hd__a21oi_1
X_17731_ _19147_/CLK _17731_/D vssd1 vssd1 vccd1 vccd1 _17731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10066_ _10129_/A vssd1 vssd1 vccd1 vccd1 _10066_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03969_ clkbuf_0__03969_/X vssd1 vssd1 vccd1 vccd1 _15689__987/A sky130_fd_sc_hd__clkbuf_16
XFILLER_208_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17662_ _17969_/CLK _17662_/D vssd1 vssd1 vccd1 vccd1 _17662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16613_ _16613_/A _16613_/B _16613_/C vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__nor3_1
X_13825_ _19147_/Q input62/X _13828_/B vssd1 vssd1 vccd1 vccd1 _13825_/X sky130_fd_sc_hd__and3_1
X_17593_ _19016_/CLK _17593_/D vssd1 vssd1 vccd1 vccd1 _17593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_104 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_115 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_126 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19332_ _19336_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_137 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_148 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13756_ _17896_/Q _13743_/B _13755_/Y _13753_/X vssd1 vssd1 vccd1 vccd1 _17896_/D
+ sky130_fd_sc_hd__a211o_1
X_10968_ hold11/A vssd1 vssd1 vccd1 vccd1 _10977_/S sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_159 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12707_ _12707_/A _12707_/B _12707_/C _12707_/D vssd1 vssd1 vccd1 vccd1 _12717_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_189_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19263_ _19266_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16475_ _16475_/A vssd1 vssd1 vccd1 vccd1 _16499_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13687_ _17872_/Q _13682_/X _13686_/Y vssd1 vssd1 vccd1 vccd1 _17872_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10899_ _18319_/Q _10898_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18214_ _18214_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
X_12638_ _12638_/A _12638_/B _12641_/D vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__and3_1
X_19194_ _19194_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__04852_ clkbuf_0__04852_/X vssd1 vssd1 vccd1 vccd1 _17083__66/A sky130_fd_sc_hd__clkbuf_16
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18145_ _18145_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
X_15357_ _18677_/Q _18583_/Q _17538_/Q _17513_/Q _15308_/A _15301_/X vssd1 vssd1 vccd1
+ vccd1 _15358_/A sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1__f__03803_ clkbuf_0__03803_/X vssd1 vssd1 vccd1 vccd1 _15439__933/A sky130_fd_sc_hd__clkbuf_16
X_12569_ _12458_/X _12459_/X _12569_/S vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18076_ _19146_/CLK _18076_/D vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15288_ _15280_/X _15287_/X _09615_/A vssd1 vssd1 vccd1 vccd1 _15288_/X sky130_fd_sc_hd__o21a_1
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14239_ _18914_/Q _18915_/Q _18916_/Q _18917_/Q _18470_/Q _15060_/A vssd1 vssd1 vccd1
+ vccd1 _14239_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14848__771 _14851__774/A vssd1 vssd1 vccd1 vccd1 _18416_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03596_ clkbuf_0__03596_/X vssd1 vssd1 vccd1 vccd1 _15138__850/A sky130_fd_sc_hd__clkbuf_16
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08800_/A vssd1 vssd1 vccd1 vccd1 _19343_/D sky130_fd_sc_hd__clkbuf_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09780_/A vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18987_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08731_ _18084_/Q _18085_/Q _18086_/Q _18087_/Q vssd1 vssd1 vccd1 vccd1 _13386_/B
+ sky130_fd_sc_hd__or4_4
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _19136_/CLK _17929_/D vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09214_ _09214_/A vssd1 vssd1 vccd1 vccd1 _19152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09145_ _18661_/Q vssd1 vssd1 vccd1 vccd1 _09145_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09076_ _09076_/A vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14749__691 _14749__691/A vssd1 vssd1 vccd1 vccd1 _18334_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _18774_/Q _09935_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__mux2_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _17922_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08929_ _09688_/A vssd1 vssd1 vccd1 vccd1 _08929_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _17778_/Q vssd1 vssd1 vccd1 vccd1 _12044_/A sky130_fd_sc_hd__inv_2
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _17935_/Q _17826_/Q vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__or2_4
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _17848_/Q vssd1 vssd1 vccd1 vccd1 _14922_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _10822_/A vssd1 vssd1 vccd1 vccd1 _18360_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _18323_/Q _14543_/X _14586_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18323_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _13541_/A _13541_/B _13541_/C _08741_/D vssd1 vssd1 vccd1 vccd1 _13571_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_213_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10753_ _10768_/S vssd1 vssd1 vccd1 vccd1 _10762_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16260_ _18443_/Q _18693_/Q _18701_/Q _18709_/Q _16198_/X _16172_/X vssd1 vssd1 vccd1
+ vccd1 _16261_/B sky130_fd_sc_hd__mux4_2
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13472_/X sky130_fd_sc_hd__buf_4
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10684_ _18415_/Q _09735_/X _10688_/S vssd1 vssd1 vccd1 vccd1 _10685_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15308_/A vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__buf_2
X_12423_ _12474_/A vssd1 vssd1 vccd1 vccd1 _12765_/S sky130_fd_sc_hd__clkbuf_2
X_16191_ _16290_/S vssd1 vssd1 vccd1 vccd1 _16191_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12354_ _17618_/Q vssd1 vssd1 vccd1 vccd1 _12707_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11305_ _11142_/X _18154_/Q _11313_/S vssd1 vssd1 vccd1 vccd1 _11306_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15073_ _16061_/A _15177_/A vssd1 vssd1 vccd1 vccd1 _18480_/D sky130_fd_sc_hd__nor2_1
X_12285_ _12280_/X _12285_/B vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _17988_/Q _14011_/X _14023_/Y vssd1 vssd1 vccd1 vccd1 _17988_/D sky130_fd_sc_hd__o21a_1
X_18901_ _18901_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11236_ _11236_/A vssd1 vssd1 vccd1 vccd1 _18181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18832_ _18832_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_1
X_11167_ _11167_/A vssd1 vssd1 vccd1 vccd1 _18211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10118_ _10117_/X _18717_/Q _10127_/S vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18763_ _18763_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ _09043_/X _18238_/Q _11098_/S vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__mux2_1
X_15975_ _16025_/B vssd1 vssd1 vccd1 vccd1 _15993_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17714_ _17714_/CLK _17714_/D vssd1 vssd1 vccd1 vccd1 _17714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14926_ _18460_/Q _14952_/B vssd1 vssd1 vccd1 vccd1 _14962_/B sky130_fd_sc_hd__and2_1
XFILLER_49_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10049_ _10049_/A _10437_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__or3_4
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18694_ _18694_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__05082_ _17415_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05082_/X sky130_fd_sc_hd__clkbuf_16
X_15091__814 _15091__814/A vssd1 vssd1 vccd1 vccd1 _18490_/CLK sky130_fd_sc_hd__inv_2
X_17645_ _17991_/CLK _17645_/D vssd1 vssd1 vccd1 vccd1 _17645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _13411_/X _13802_/X _13805_/X vssd1 vssd1 vccd1 vccd1 _13808_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17576_ _17576_/CLK _17576_/D vssd1 vssd1 vccd1 vccd1 _17576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19315_ _19315_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13739_ _13757_/B vssd1 vssd1 vccd1 vccd1 _13743_/B sky130_fd_sc_hd__clkbuf_2
X_16527_ _16527_/A vssd1 vssd1 vccd1 vccd1 _18991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19246_ _19246_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ _18974_/Q _16458_/B vssd1 vssd1 vccd1 vccd1 _16466_/C sky130_fd_sc_hd__and2_1
XFILLER_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17400__92 _17402__94/A vssd1 vssd1 vccd1 vccd1 _19305_/CLK sky130_fd_sc_hd__inv_2
X_19177_ _19177_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_1
X_16389_ _18977_/Q _16389_/B _16389_/C vssd1 vssd1 vccd1 vccd1 _16420_/B sky130_fd_sc_hd__and3_1
XFILLER_129_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18128_ _18128_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176__453 _14177__454/A vssd1 vssd1 vccd1 vccd1 _18061_/CLK sky130_fd_sc_hd__inv_2
X_18059_ _18059_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _18797_/Q _09723_/X _09907_/S vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09832_ _09682_/X _18817_/Q _09836_/S vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09763_ _09763_/A vssd1 vssd1 vccd1 vccd1 _18846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _09694_/A vssd1 vssd1 vccd1 vccd1 _09694_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_230_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16734__347 _16735__348/A vssd1 vssd1 vccd1 vccd1 _19126_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ _19186_/Q _09127_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09059_ _09770_/A vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_151_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12070_ _12099_/S _12064_/X _12069_/X vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__o21ai_4
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11021_ _11021_/A vssd1 vssd1 vccd1 vccd1 _18268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12972_ _12957_/X _12972_/B vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__and2b_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03806_ clkbuf_0__03806_/X vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11923_ _11920_/X _11921_/X _11957_/S vssd1 vssd1 vccd1 vccd1 _11923_/X sky130_fd_sc_hd__mux2_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14707_/X _14710_/X _14730_/S vssd1 vssd1 vccd1 vccd1 _14711_/X sky130_fd_sc_hd__mux2_2
XFILLER_206_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _17430_/A vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _18587_/Q _18301_/Q _17567_/Q _18838_/Q _14615_/X _14641_/X vssd1 vssd1 vccd1
+ vccd1 _14642_/X sky130_fd_sc_hd__mux4_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11854_ _13279_/A _11854_/B vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__and2_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10805_/A vssd1 vssd1 vccd1 vccd1 _18366_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17361_ _19279_/Q _12206_/X _12212_/X _19283_/Q _17360_/X vssd1 vssd1 vccd1 vccd1
+ _17361_/Y sky130_fd_sc_hd__a221oi_1
X_14573_ _14662_/S vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11785_ _11815_/A vssd1 vssd1 vccd1 vccd1 _11785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_242_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19100_ _19100_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13524_ _13394_/X _13523_/X _13513_/X vssd1 vssd1 vccd1 vccd1 _13524_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_0__f__03599_ clkbuf_0__03599_/X vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17292_ _19265_/Q _17288_/B _17288_/C _17284_/C _19266_/Q vssd1 vssd1 vccd1 vccd1
+ _17292_/X sky130_fd_sc_hd__a41o_1
XFILLER_158_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10736_ _18394_/Q _10690_/X _10744_/S vssd1 vssd1 vccd1 vccd1 _10737_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19031_ _19040_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
X_16243_ _18450_/Q _19088_/Q _19125_/Q _18434_/Q _16144_/X _16108_/X vssd1 vssd1 vccd1
+ vccd1 _16243_/X sky130_fd_sc_hd__mux4_2
X_13455_ _17800_/Q _13457_/B vssd1 vssd1 vccd1 vccd1 _13455_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _10667_/A vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12406_ _18009_/Q vssd1 vssd1 vccd1 vccd1 _12407_/A sky130_fd_sc_hd__clkinv_2
XFILLER_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16174_ _16223_/A _16174_/B vssd1 vssd1 vccd1 vccd1 _16174_/Y sky130_fd_sc_hd__nor2_1
X_13386_ _18081_/Q _13386_/B _13386_/C _13386_/D vssd1 vssd1 vccd1 vccd1 _13387_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_86_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10598_ _09051_/X _18485_/Q hold19/X vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15125_ _15131_/A vssd1 vssd1 vccd1 vccd1 _15125_/X sky130_fd_sc_hd__buf_1
XFILLER_86_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput108 _11763_/X vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_2
XFILLER_217_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput119 _11724_/X vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_2
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14353__538 _14354__539/A vssd1 vssd1 vccd1 vccd1 _18173_/CLK sky130_fd_sc_hd__inv_2
XFILLER_142_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03602_ _15168_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03602_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15056_ _18482_/Q _18472_/Q _15060_/A _15055_/Y _15076_/A vssd1 vssd1 vccd1 vccd1
+ _15057_/B sky130_fd_sc_hd__a311o_1
XFILLER_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12268_ _12263_/X _12268_/B vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__and2b_1
X_14007_ _17982_/Q _13989_/X _14006_/Y vssd1 vssd1 vccd1 vccd1 _17982_/D sky130_fd_sc_hd__o21a_1
XFILLER_218_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11219_ _11219_/A vssd1 vssd1 vccd1 vccd1 _18188_/D sky130_fd_sc_hd__clkbuf_1
X_12199_ _12199_/A vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput90 _11749_/X vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_233_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18815_ _18815_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18746_ _18746_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03395_ _14745_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03395_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15958_ _18888_/Q _15958_/B vssd1 vssd1 vccd1 vccd1 _15962_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _17847_/Q _14909_/B vssd1 vssd1 vccd1 vccd1 _14910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18677_ _18677_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17628_ _17629_/CLK _17628_/D vssd1 vssd1 vccd1 vccd1 _17628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17559_ _18027_/CLK _17559_/D vssd1 vssd1 vccd1 vccd1 _17559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19229_ _19252_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_1
X_17385__80 _17386__81/A vssd1 vssd1 vccd1 vccd1 _19293_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04849_ _17068_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04849_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14254__458 _14255__459/A vssd1 vssd1 vccd1 vccd1 _18093_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150__434 _14150__434/A vssd1 vssd1 vccd1 vccd1 _18042_/CLK sky130_fd_sc_hd__inv_2
X_09815_ _09815_/A vssd1 vssd1 vccd1 vccd1 _18825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09746_ _09768_/S vssd1 vssd1 vccd1 vccd1 _09759_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09674_/X _18905_/Q _09689_/S vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04571_ clkbuf_0__04571_/X vssd1 vssd1 vccd1 vccd1 _16658_/A sky130_fd_sc_hd__clkbuf_16
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11570_ _11570_/A vssd1 vssd1 vccd1 vccd1 _17587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ _10521_/A vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13240_ _13786_/A vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__buf_4
XFILLER_196_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10452_ _10132_/X _18549_/Q _10454_/S vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13171_ _13216_/B vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__buf_2
X_10383_ _10383_/A vssd1 vssd1 vccd1 vccd1 _18580_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__04005_ clkbuf_0__04005_/X vssd1 vssd1 vccd1 vccd1 _15843_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ _12184_/A _12199_/A _12122_/C vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_33_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _19340_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12053_ _12006_/X _12008_/X _12051_/X _12052_/X _12091_/A _12045_/S vssd1 vssd1 vccd1
+ vccd1 _12053_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16930_ _18215_/Q _18199_/Q _18488_/Q _18191_/Q _09852_/A _09858_/A vssd1 vssd1 vccd1
+ vccd1 _16930_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11004_ _18275_/Q _09145_/X _11004_/S vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__mux2_1
X_16861_ _16818_/X _16859_/X _16860_/X vssd1 vssd1 vccd1 vccd1 _16861_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18600_ _18600_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15812_ _16063_/A vssd1 vssd1 vccd1 vccd1 _15812_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16792_ _19135_/Q _16767_/S _16788_/A _16791_/X vssd1 vssd1 vccd1 vccd1 _16792_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__04838_ clkbuf_0__04838_/X vssd1 vssd1 vccd1 vccd1 _17037_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18531_ _18531_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03180_ _14437_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03180_/X sky130_fd_sc_hd__clkbuf_16
X_12955_ _12911_/X _12955_/B vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__and2b_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07557_ clkbuf_0__07557_/X vssd1 vssd1 vccd1 vccd1 _12329__391/A sky130_fd_sc_hd__clkbuf_16
XFILLER_46_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11906_ _12076_/S vssd1 vssd1 vccd1 vccd1 _11907_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _18462_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12886_ _12877_/X _12886_/B vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__and2b_1
XFILLER_179_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15686_/A vssd1 vssd1 vccd1 vccd1 _15674_/X sky130_fd_sc_hd__buf_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _11837_/A vssd1 vssd1 vccd1 vccd1 _11837_/Y sky130_fd_sc_hd__inv_2
X_14625_ _18405_/Q _18397_/Q _19310_/Q _17714_/Q _14594_/X _14595_/X vssd1 vssd1 vccd1
+ vccd1 _14625_/X sky130_fd_sc_hd__mux4_1
X_18393_ _18393_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17344_ _17757_/Q _19286_/Q _17350_/S vssd1 vssd1 vccd1 vccd1 _17345_/B sky130_fd_sc_hd__mux2_1
X_14556_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__buf_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _18003_/Q _17885_/Q vssd1 vssd1 vccd1 vccd1 _11769_/A sky130_fd_sc_hd__and2b_1
XFILLER_144_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03982_ clkbuf_0__03982_/X vssd1 vssd1 vccd1 vccd1 _15767_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13507_ _17814_/Q _13446_/X _13507_/S vssd1 vssd1 vccd1 vccd1 _13508_/B sky130_fd_sc_hd__mux2_1
X_10719_ _10719_/A vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__clkbuf_1
X_17275_ _17288_/D vssd1 vssd1 vccd1 vccd1 _17284_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14487_ _14487_/A vssd1 vssd1 vccd1 vccd1 _14487_/X sky130_fd_sc_hd__buf_1
X_11699_ _18412_/Q _11694_/C _11698_/Y vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19014_ _19014_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
X_13438_ _13447_/S vssd1 vssd1 vccd1 vccd1 _13444_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16226_ _16191_/X _16219_/Y _16221_/Y _16223_/Y _16225_/Y vssd1 vssd1 vccd1 vccd1
+ _16226_/X sky130_fd_sc_hd__o32a_2
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16157_ _18626_/Q _18501_/Q _18907_/Q _18509_/Q _16155_/X _16156_/X vssd1 vssd1 vccd1
+ vccd1 _16157_/X sky130_fd_sc_hd__mux4_1
X_13369_ _13748_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _18466_/Q _14967_/X _15038_/Y _15026_/X vssd1 vssd1 vccd1 vccd1 _15040_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03416_ clkbuf_0__03416_/X vssd1 vssd1 vccd1 vccd1 _14850__773/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09600_ _09600_/A vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _09531_/A vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18729_ _18729_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138__850 _15138__850/A vssd1 vssd1 vccd1 vccd1 _18526_/CLK sky130_fd_sc_hd__inv_2
XFILLER_243_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09462_ _09462_/A vssd1 vssd1 vccd1 vccd1 _19046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _09393_/A vssd1 vssd1 vccd1 vccd1 _19068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15442__935 _15444__937/A vssd1 vssd1 vccd1 vccd1 _18622_/CLK sky130_fd_sc_hd__inv_2
XFILLER_193_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16699__323 _16700__324/A vssd1 vssd1 vccd1 vccd1 _19098_/CLK sky130_fd_sc_hd__inv_2
XFILLER_248_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09729_ _10701_/A vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__buf_4
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _12746_/C _12746_/D vssd1 vssd1 vccd1 vccd1 _12742_/A sky130_fd_sc_hd__and2_1
XFILLER_167_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12672_/B _12673_/A _12670_/Y vssd1 vssd1 vccd1 vccd1 _17609_/D sky130_fd_sc_hd__a21oi_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11622_ _11622_/A vssd1 vssd1 vccd1 vccd1 _17547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _17709_/Q _10895_/X _11557_/S vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ _10129_/X _18526_/Q _10508_/S vssd1 vssd1 vccd1 vccd1 _10505_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ _11484_/A vssd1 vssd1 vccd1 vccd1 _18052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16011_ _16008_/X _16009_/Y _16010_/X vssd1 vssd1 vccd1 vccd1 _18870_/D sky130_fd_sc_hd__a21oi_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13223_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13293_/A sky130_fd_sc_hd__clkbuf_2
X_10435_ _09971_/A _09255_/A _10407_/X vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__o21ai_1
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13154_ input56/X _13210_/B vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__nand2_4
XFILLER_163_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _18587_/Q _09735_/X _10370_/S vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12105_ _11912_/X _11926_/X _12111_/S vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__mux2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _17697_/Q _13085_/B vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__xor2_1
X_17962_ _19037_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ _10297_/A vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12036_ _11921_/X _11924_/X _12036_/S vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__mux2_1
X_16913_ _16818_/X _16912_/X _16860_/X vssd1 vssd1 vccd1 vccd1 _16913_/Y sky130_fd_sc_hd__o21ai_1
X_17893_ _19109_/CLK _17893_/D vssd1 vssd1 vccd1 vccd1 _17893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14842__766 _14843__767/A vssd1 vssd1 vccd1 vccd1 _18409_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16842_/X _16843_/X _16982_/A vssd1 vssd1 vccd1 vccd1 _16844_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16775_ _16775_/A _16775_/B vssd1 vssd1 vccd1 vccd1 _19132_/D sky130_fd_sc_hd__nor2_1
XFILLER_93_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13987_ _14031_/A _13987_/B _14076_/C vssd1 vssd1 vccd1 vccd1 _13995_/A sky130_fd_sc_hd__and3_2
XFILLER_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18514_ _18514_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03163_ _14355_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03163_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _17662_/Q _13093_/B vssd1 vssd1 vccd1 vccd1 _12941_/B sky130_fd_sc_hd__xnor2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03094_ _14159_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03094_/X sky130_fd_sc_hd__clkbuf_16
X_18445_ _18445_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
X_15806__125 _15807__126/A vssd1 vssd1 vccd1 vccd1 _18797_/CLK sky130_fd_sc_hd__inv_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12830_/X _12869_/B vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__and2b_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14608_ _19149_/Q _18414_/Q _18308_/Q _18292_/Q _09443_/A _14575_/X vssd1 vssd1 vccd1
+ vccd1 _14609_/B sky130_fd_sc_hd__mux4_1
XFILLER_222_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18376_ _18376_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
X_15588_ _15586_/X _15587_/Y _15581_/X vssd1 vssd1 vccd1 vccd1 _18651_/D sky130_fd_sc_hd__a21oi_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ _17762_/Q _19281_/Q _17333_/S vssd1 vssd1 vccd1 vccd1 _17328_/B sky130_fd_sc_hd__mux2_1
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03965_ clkbuf_0__03965_/X vssd1 vssd1 vccd1 vccd1 _15664__966/A sky130_fd_sc_hd__clkbuf_16
XFILLER_175_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ _17262_/B _17262_/C _17258_/C vssd1 vssd1 vccd1 vccd1 _17264_/B sky130_fd_sc_hd__and3_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16209_ _18628_/Q _18503_/Q _18909_/Q _18511_/Q _16155_/X _16156_/X vssd1 vssd1 vccd1
+ vccd1 _16209_/X sky130_fd_sc_hd__mux4_1
X_17189_ _17195_/A _17189_/B _17189_/C vssd1 vssd1 vccd1 vccd1 _17190_/A sky130_fd_sc_hd__and3b_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_7_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_7_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ _19269_/Q _08961_/X _08968_/S vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08893_ _19307_/Q _08724_/X _08901_/S vssd1 vssd1 vccd1 vccd1 _08894_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__07167_ clkbuf_0__07167_/X vssd1 vssd1 vccd1 vccd1 _17043_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14366__548 _14367__549/A vssd1 vssd1 vccd1 vccd1 _18183_/CLK sky130_fd_sc_hd__inv_2
XFILLER_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09514_ _19002_/Q _09489_/X _09518_/S vssd1 vssd1 vccd1 vccd1 _09515_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _14651_/A _09456_/A vssd1 vssd1 vccd1 vccd1 _09453_/B sky130_fd_sc_hd__nand2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09376_ _09376_/A vssd1 vssd1 vccd1 vccd1 _19075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15704__999 _15704__999/A vssd1 vssd1 vccd1 vccd1 _18716_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03152_ clkbuf_0__03152_/X vssd1 vssd1 vccd1 vccd1 _14299__494/A sky130_fd_sc_hd__clkbuf_16
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10220_ _10220_/A hold2/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__nor2_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10151_ _18705_/Q _10066_/X _10155_/S vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310__503 _14310__503/A vssd1 vssd1 vccd1 vccd1 _18138_/CLK sky130_fd_sc_hd__inv_2
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10082_ _18732_/Q _10057_/X _10086_/S vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03985_ clkbuf_0__03985_/X vssd1 vssd1 vccd1 vccd1 _15772__1054/A sky130_fd_sc_hd__clkbuf_16
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13910_ _13529_/X _13908_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13910_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13841_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__buf_2
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14267__468 _14268__469/A vssd1 vssd1 vccd1 vccd1 _18103_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13772_ _13281_/X _13771_/X _13701_/X vssd1 vssd1 vccd1 vccd1 _13772_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16560_ _16560_/A vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__clkbuf_1
X_10984_ _10984_/A vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15511_ _15511_/A _15511_/B vssd1 vssd1 vccd1 vccd1 _15512_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12723_ _12723_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _17624_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16491_ _18981_/Q _16491_/B vssd1 vssd1 vccd1 vccd1 _16493_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17506__4 _17506__4/A vssd1 vssd1 vccd1 vccd1 _19348_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18230_ _18230_/CLK _18230_/D vssd1 vssd1 vccd1 vccd1 _18230_/Q sky130_fd_sc_hd__dfxtp_1
X_12654_ _12658_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _17604_/D sky130_fd_sc_hd__nor2_1
XFILLER_188_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11605_ _17571_/Q _10695_/A _11611_/S vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18161_ _18161_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
X_12585_ _12466_/X _12463_/X _12464_/X _12458_/X _12569_/S _12502_/A vssd1 vssd1 vccd1
+ vccd1 _12585_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15373_ _18835_/Q _18827_/Q _18819_/Q _18686_/Q _15299_/X _15230_/X vssd1 vssd1 vccd1
+ vccd1 _15373_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0__f__03419_ clkbuf_0__03419_/X vssd1 vssd1 vccd1 vccd1 _14869__789/A sky130_fd_sc_hd__clkbuf_16
XFILLER_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17112_ _17117_/C _17112_/B vssd1 vssd1 vccd1 vccd1 _17113_/A sky130_fd_sc_hd__and2b_1
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _11536_/A vssd1 vssd1 vccd1 vccd1 _17717_/D sky130_fd_sc_hd__clkbuf_1
X_14324_ _14355_/A vssd1 vssd1 vccd1 vccd1 _14324_/X sky130_fd_sc_hd__buf_1
X_18092_ _18092_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17043_ _17043_/A vssd1 vssd1 vccd1 vccd1 _17043_/X sky130_fd_sc_hd__buf_1
X_14471__632 _14472__633/A vssd1 vssd1 vccd1 vccd1 _18267_/CLK sky130_fd_sc_hd__inv_2
X_11467_ _11335_/X _18059_/Q _11467_/S vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _13812_/A vssd1 vssd1 vccd1 vccd1 _13755_/A sky130_fd_sc_hd__buf_4
X_10418_ _18564_/Q vssd1 vssd1 vccd1 vccd1 _16182_/A sky130_fd_sc_hd__clkbuf_4
X_14186_ _12828_/A input78/X input54/X _14186_/D vssd1 vssd1 vccd1 vccd1 _14231_/A
+ sky130_fd_sc_hd__and4b_2
X_11398_ _11341_/X _18116_/Q _11400_/S vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13137_ _13216_/B vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10349_ _18594_/Q _10348_/X _10352_/S vssd1 vssd1 vccd1 vccd1 _10350_/A sky130_fd_sc_hd__mux2_1
X_18994_ _18996_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735__1024 _15735__1024/A vssd1 vssd1 vccd1 vccd1 _18741_/CLK sky130_fd_sc_hd__inv_2
XFILLER_239_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14170__448 _14171__449/A vssd1 vssd1 vccd1 vccd1 _18056_/CLK sky130_fd_sc_hd__inv_2
X_13068_ _13066_/X _13068_/B vssd1 vssd1 vccd1 vccd1 _13069_/A sky130_fd_sc_hd__and2b_1
X_17945_ _17945_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12019_ _11912_/X _11923_/X _11926_/X _12017_/X _12116_/A _12018_/X vssd1 vssd1 vccd1
+ vccd1 _12020_/B sky130_fd_sc_hd__mux4_1
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17876_ _17878_/CLK _17876_/D vssd1 vssd1 vccd1 vccd1 _17876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16827_ _16881_/A vssd1 vssd1 vccd1 vccd1 _16827_/X sky130_fd_sc_hd__buf_2
XFILLER_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04164_ clkbuf_0__04164_/X vssd1 vssd1 vccd1 vccd1 _16079__194/A sky130_fd_sc_hd__clkbuf_16
XFILLER_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17407__98 _17408__99/A vssd1 vssd1 vccd1 vccd1 _19311_/CLK sky130_fd_sc_hd__inv_2
X_16758_ _19130_/Q _16771_/B vssd1 vssd1 vccd1 vccd1 _16758_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03146_ _14263_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03146_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_222_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16689_ _16689_/A _16689_/B _16737_/B vssd1 vssd1 vccd1 vccd1 _16689_/X sky130_fd_sc_hd__and3_1
XFILLER_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ _18559_/Q vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__inv_2
XFILLER_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18428_ _18428_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _09161_/A vssd1 vssd1 vccd1 vccd1 _19175_/D sky130_fd_sc_hd__clkbuf_1
X_18359_ _18359_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _10695_/A vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__buf_2
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03979_ _15736_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03979_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09994_ _10157_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10010_/S sky130_fd_sc_hd__nor2_2
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ _09745_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08968_/S sky130_fd_sc_hd__nor2_2
XFILLER_229_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _08876_/A vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08199_ clkbuf_0__08199_/X vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _08937_/X _19052_/Q _09430_/S vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ _10691_/B _11583_/B vssd1 vssd1 vccd1 vccd1 _09375_/S sky130_fd_sc_hd__nor2_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12370_ _18010_/Q vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ _11321_/A vssd1 vssd1 vccd1 vccd1 _11321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535__684 _14535__684/A vssd1 vssd1 vccd1 vccd1 _18319_/CLK sky130_fd_sc_hd__inv_2
X_14040_ _13746_/A _14039_/X _14034_/X vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11252_ _11252_/A vssd1 vssd1 vccd1 vccd1 _18174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10203_ _18686_/Q _09744_/X _10211_/S vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _11183_/A vssd1 vssd1 vccd1 vccd1 _18204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _10134_/A vssd1 vssd1 vccd1 vccd1 _18712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _18867_/Q _15991_/B vssd1 vssd1 vccd1 vccd1 _16002_/C sky130_fd_sc_hd__and2_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17730_ _19147_/CLK _17730_/D vssd1 vssd1 vccd1 vccd1 _17730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _18457_/Q _14942_/B _14942_/C vssd1 vssd1 vccd1 vccd1 _14950_/A sky130_fd_sc_hd__and3_1
X_10065_ _10065_/A vssd1 vssd1 vccd1 vccd1 _18738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03968_ clkbuf_0__03968_/X vssd1 vssd1 vccd1 vccd1 _15682__981/A sky130_fd_sc_hd__clkbuf_16
XFILLER_235_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _18006_/CLK _17661_/D vssd1 vssd1 vccd1 vccd1 _17661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19400_ input21/X vssd1 vssd1 vccd1 vccd1 _19400_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16612_ _19034_/Q _16608_/B _19035_/Q vssd1 vssd1 vccd1 vccd1 _16613_/C sky130_fd_sc_hd__a21oi_1
XFILLER_211_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13824_ _17918_/Q _13820_/Y _13823_/X _13753_/X vssd1 vssd1 vccd1 vccd1 _17918_/D
+ sky130_fd_sc_hd__a211o_1
X_17592_ _19016_/CLK _17592_/D vssd1 vssd1 vccd1 vccd1 _17592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_105 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_116 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19331_ _19336_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_127 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16543_ _16543_/A vssd1 vssd1 vccd1 vccd1 _16543_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_138 _11838_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13755_ _13755_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13755_/Y sky130_fd_sc_hd__nor2_1
X_10967_ _10967_/A _10967_/B vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__nor2_2
XINSDIODE2_149 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12706_/A _12706_/B vssd1 vssd1 vccd1 vccd1 _12707_/D sky130_fd_sc_hd__and2_1
X_19262_ _19266_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15842__144 _15842__144/A vssd1 vssd1 vccd1 vccd1 _18819_/CLK sky130_fd_sc_hd__inv_2
X_16474_ _16498_/A _16474_/B _16482_/C vssd1 vssd1 vccd1 vccd1 _16474_/X sky130_fd_sc_hd__or3_1
XFILLER_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13686_ _13256_/X _13683_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _13686_/Y sky130_fd_sc_hd__a21oi_1
X_10898_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _10898_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _18213_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _12637_/A vssd1 vssd1 vccd1 vccd1 _17599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__04851_ clkbuf_0__04851_/X vssd1 vssd1 vccd1 vccd1 _17078__62/A sky130_fd_sc_hd__clkbuf_16
X_19193_ _19193_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18144_ _18144_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03802_ clkbuf_0__03802_/X vssd1 vssd1 vccd1 vccd1 _15433__928/A sky130_fd_sc_hd__clkbuf_16
X_12568_ _12568_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12568_/Y sky130_fd_sc_hd__nor2_1
X_15356_ _18834_/Q _18826_/Q _18818_/Q _18685_/Q _15299_/X _15230_/X vssd1 vssd1 vccd1
+ vccd1 _15356_/X sky130_fd_sc_hd__mux4_2
XFILLER_106_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11519_ _18036_/Q _11332_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14317__509 _14317__509/A vssd1 vssd1 vccd1 vccd1 _18144_/CLK sky130_fd_sc_hd__inv_2
X_18075_ _18869_/CLK _18075_/D vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_2
X_12499_ _18006_/Q _18005_/Q _12763_/A vssd1 vssd1 vccd1 vccd1 _12510_/C sky130_fd_sc_hd__or3b_1
X_15287_ _15281_/X _15282_/X _15286_/Y vssd1 vssd1 vccd1 vccd1 _15287_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14238_ _18471_/Q vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03595_ clkbuf_0__03595_/X vssd1 vssd1 vccd1 vccd1 _15134__847/A sky130_fd_sc_hd__clkbuf_16
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18987_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08730_ _08855_/C vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17928_ _19136_/CLK _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17859_ _17953_/CLK _17859_/D vssd1 vssd1 vccd1 vccd1 _17859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478__638 _14479__639/A vssd1 vssd1 vccd1 vccd1 _18273_/CLK sky130_fd_sc_hd__inv_2
X_09213_ _19152_/Q _09100_/X _09215_/S vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09144_ _09144_/A vssd1 vssd1 vccd1 vccd1 _19181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ _19197_/Q _08883_/X _09077_/S vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09977_ _09992_/S vssd1 vssd1 vccd1 vccd1 _09986_/S sky130_fd_sc_hd__buf_2
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _18883_/Q vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_218_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16069__185 _16071__187/A vssd1 vssd1 vccd1 vccd1 _18890_/CLK sky130_fd_sc_hd__inv_2
XFILLER_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ _08728_/X _08857_/X _11675_/A vssd1 vssd1 vccd1 vccd1 _16559_/B sky130_fd_sc_hd__a21oi_4
XFILLER_242_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _11870_/A vssd1 vssd1 vccd1 vccd1 _11870_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18006_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _18360_/Q _10797_/X _10825_/S vssd1 vssd1 vccd1 vccd1 _10822_/A sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10752_ _10752_/A hold13/X vssd1 vssd1 vccd1 vccd1 _10768_/S sky130_fd_sc_hd__nor2_2
X_13540_ _13540_/A _13540_/B _13488_/A vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__or3b_1
XFILLER_197_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15734__1023 _15735__1024/A vssd1 vssd1 vccd1 vccd1 _18740_/CLK sky130_fd_sc_hd__inv_2
X_13471_ _17804_/Q _13477_/B vssd1 vssd1 vccd1 vccd1 _13471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10683_ _10683_/A vssd1 vssd1 vccd1 vccd1 _18416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12422_ _18010_/Q vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__clkbuf_2
X_15210_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _15308_/A sky130_fd_sc_hd__buf_4
X_16190_ _16291_/A vssd1 vssd1 vccd1 vccd1 _16190_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12353_ _17616_/Q _17617_/Q _12443_/A vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04167_ clkbuf_0__04167_/X vssd1 vssd1 vccd1 vccd1 _16307__209/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11304_ _11319_/S vssd1 vssd1 vccd1 vccd1 _11313_/S sky130_fd_sc_hd__clkbuf_2
X_16310__210 _16314__214/A vssd1 vssd1 vccd1 vccd1 _18926_/CLK sky130_fd_sc_hd__inv_2
XFILLER_154_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15072_ _16060_/A _15177_/A vssd1 vssd1 vccd1 vccd1 _18479_/D sky130_fd_sc_hd__nor2_1
X_12284_ _17560_/Q _18017_/Q _12287_/S vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__mux2_1
X_14023_ _13783_/X _14017_/X _14020_/X vssd1 vssd1 vccd1 vccd1 _14023_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18900_ _18900_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_1
X_11235_ _11159_/X _18181_/Q _11239_/S vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__mux2_1
X_17002__351 _17002__351/A vssd1 vssd1 vccd1 vccd1 _19150_/CLK sky130_fd_sc_hd__inv_2
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18831_ _18831_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_1
X_11166_ _11165_/X _18211_/Q _11166_/S vssd1 vssd1 vccd1 vccd1 _11167_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108__414 _13108__414/A vssd1 vssd1 vccd1 vccd1 _17710_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10117_ _10117_/A vssd1 vssd1 vccd1 vccd1 _10117_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18762_ _18762_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ _11097_/A vssd1 vssd1 vccd1 vccd1 _18239_/D sky130_fd_sc_hd__clkbuf_1
X_15974_ _15986_/A _15974_/B _15985_/C vssd1 vssd1 vccd1 vccd1 _15974_/X sky130_fd_sc_hd__or3_1
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17713_/CLK _17713_/D vssd1 vssd1 vccd1 vccd1 _17713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14925_ _17853_/Q _14930_/A vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10048_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10048_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18693_ _18693_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__05081_ _17409_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05081_/X sky130_fd_sc_hd__clkbuf_16
X_17644_ _17991_/CLK _17644_/D vssd1 vssd1 vccd1 vccd1 _17644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13807_ _17912_/Q _13796_/X _13806_/Y vssd1 vssd1 vccd1 vccd1 _17912_/D sky130_fd_sc_hd__o21a_1
X_17575_ _17575_/CLK _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ _19262_/Q vssd1 vssd1 vccd1 vccd1 _17276_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19314_ _19314_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16526_ input68/X _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16527_/A sky130_fd_sc_hd__and3_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13738_ _13757_/B vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15132__845 _15134__847/A vssd1 vssd1 vccd1 vccd1 _18521_/CLK sky130_fd_sc_hd__inv_2
XFILLER_232_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19245_ _19247_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16457_ _18974_/Q _16458_/B vssd1 vssd1 vccd1 vccd1 _16459_/B sky130_fd_sc_hd__nor2_1
X_13669_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13669_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19176_ _19176_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_1
X_16388_ _16389_/B _16389_/C _18977_/Q vssd1 vssd1 vccd1 vccd1 _16420_/A sky130_fd_sc_hd__a21oi_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18127_ _18127_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_1
X_15339_ _18833_/Q _18825_/Q _18817_/Q _18684_/Q _15299_/X _15230_/X vssd1 vssd1 vccd1
+ vccd1 _15339_/X sky130_fd_sc_hd__mux4_2
XFILLER_247_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18058_ _18058_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09900_ _09900_/A vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09831_ _09831_/A vssd1 vssd1 vccd1 vccd1 _18818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ _18846_/Q _09761_/X _09768_/S vssd1 vssd1 vccd1 vccd1 _09763_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14484__642 _14484__642/A vssd1 vssd1 vccd1 vccd1 _18277_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09693_ _09693_/A vssd1 vssd1 vccd1 vccd1 _18900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16693__318 _16694__319/A vssd1 vssd1 vccd1 vccd1 _19093_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15406__906 _15409__909/A vssd1 vssd1 vccd1 vccd1 _18593_/CLK sky130_fd_sc_hd__inv_2
XFILLER_194_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _18667_/Q vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09058_ _09770_/B vssd1 vssd1 vccd1 vccd1 _10770_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15791__113 _15792__114/A vssd1 vssd1 vccd1 vccd1 _18785_/CLK sky130_fd_sc_hd__inv_2
XFILLER_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11020_ _09051_/X _18268_/Q _11022_/S vssd1 vssd1 vccd1 vccd1 _11021_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12971_ _17960_/Q _17677_/Q _12976_/S vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__mux2_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03805_ clkbuf_0__03805_/X vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_246_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14708_/X _14709_/X _14729_/S vssd1 vssd1 vccd1 vccd1 _14710_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11922_ _12008_/S vssd1 vssd1 vccd1 vccd1 _11957_/S sky130_fd_sc_hd__buf_2
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14797__730 _14799__732/A vssd1 vssd1 vccd1 vccd1 _18373_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14641_/A vssd1 vssd1 vccd1 vccd1 _14641_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _17920_/Q _11839_/X _11840_/X _17901_/Q vssd1 vssd1 vccd1 vccd1 _11854_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17360_ _19290_/Q _12185_/A _12204_/X _19282_/Q vssd1 vssd1 vccd1 vccd1 _17360_/X
+ sky130_fd_sc_hd__a22o_1
X_10804_ _18366_/Q _10803_/X _10804_/S vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11784_ _11837_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__or2_1
X_14572_ _14572_/A vssd1 vssd1 vccd1 vccd1 _14662_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03598_ clkbuf_0__03598_/X vssd1 vssd1 vccd1 vccd1 _15154__864/A sky130_fd_sc_hd__clkbuf_16
X_13523_ _13523_/A vssd1 vssd1 vccd1 vccd1 _13523_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17291_ _19266_/Q vssd1 vssd1 vccd1 vccd1 _17291_/Y sky130_fd_sc_hd__inv_2
X_10735_ _10750_/S vssd1 vssd1 vccd1 vccd1 _10744_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19030_ _19040_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _16280_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16242_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13454_ _13155_/X _13437_/X _13453_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _17799_/D
+ sky130_fd_sc_hd__a211oi_1
X_10666_ _18423_/Q _09735_/X _10670_/S vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12405_ _12405_/A vssd1 vssd1 vccd1 vccd1 _12405_/Y sky130_fd_sc_hd__inv_2
X_13385_ _18080_/Q _13874_/B vssd1 vssd1 vccd1 vccd1 _13386_/D sky130_fd_sc_hd__nand2_1
XFILLER_16_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16173_ _18439_/Q _18689_/Q _18697_/Q _18705_/Q _16112_/X _16172_/X vssd1 vssd1 vccd1
+ vccd1 _16174_/B sky130_fd_sc_hd__mux4_1
XFILLER_126_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10597_ _10597_/A vssd1 vssd1 vccd1 vccd1 _18486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15124_/A vssd1 vssd1 vccd1 vccd1 _15124_/X sky130_fd_sc_hd__buf_1
Xoutput109 _11759_/X vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_2
XFILLER_142_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03601_ _15162_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03601_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12267_ _17555_/Q _18022_/Q _12270_/S vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__mux2_1
X_15055_ _18470_/Q vssd1 vssd1 vccd1 vccd1 _15055_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14006_ _13812_/X _13995_/X _14005_/X vssd1 vssd1 vccd1 vccd1 _14006_/Y sky130_fd_sc_hd__a21oi_1
X_11218_ _18188_/Q _11062_/X _11220_/S vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12198_ _12198_/A _12198_/B _12198_/C _12198_/D vssd1 vssd1 vccd1 vccd1 _12218_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput80 _11775_/X vssd1 vssd1 vccd1 vccd1 flash_io0_read sky130_fd_sc_hd__buf_2
Xoutput91 _11745_/X vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18814_ _18814_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_1
X_11149_ _11149_/A vssd1 vssd1 vccd1 vccd1 _18217_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18745_ _18745_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _18889_/Q _16063_/B vssd1 vssd1 vccd1 vccd1 _15958_/B sky130_fd_sc_hd__and2_1
XFILLER_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ _14922_/B _14936_/A vssd1 vssd1 vccd1 vccd1 _14909_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18676_ _18676_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17627_ _17629_/CLK _17627_/D vssd1 vssd1 vccd1 vccd1 _17627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _14870_/A vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__buf_1
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__04015_ _15880_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04015_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ _18027_/CLK _17558_/D vssd1 vssd1 vccd1 vccd1 _17558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18869_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16509_ _16511_/B _16505_/X _16508_/Y _14589_/X vssd1 vssd1 vccd1 vccd1 _18984_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16317__216 _16318__217/A vssd1 vssd1 vccd1 vccd1 _18932_/CLK sky130_fd_sc_hd__inv_2
X_17489_ _19337_/Q _17489_/B vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__xnor2_1
XFILLER_176_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19228_ _19252_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17009__357 _17011__359/A vssd1 vssd1 vccd1 vccd1 _19156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19159_ _19159_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04848_ _17062_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04848_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15659__963 _15660__964/A vssd1 vssd1 vccd1 vccd1 _18680_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _09682_/X _18825_/Q _09818_/S vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15733__1022 _15735__1024/A vssd1 vssd1 vccd1 vccd1 _18739_/CLK sky130_fd_sc_hd__inv_2
XFILLER_219_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _09745_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09768_/S sky130_fd_sc_hd__nor2_2
XFILLER_223_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09698_/S vssd1 vssd1 vccd1 vccd1 _09689_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_243_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__04570_ clkbuf_0__04570_/X vssd1 vssd1 vccd1 vccd1 _16643__283/A sky130_fd_sc_hd__clkbuf_16
XFILLER_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ _18519_/Q _10342_/X _10520_/S vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _10451_/A vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ _13212_/B vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10382_ _08795_/X _18580_/Q _10382_/S vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__04004_ clkbuf_0__04004_/X vssd1 vssd1 vccd1 vccd1 _15826__131/A sky130_fd_sc_hd__clkbuf_16
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12195_/A _12189_/A _12205_/A _12121_/D vssd1 vssd1 vccd1 vccd1 _12122_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _19229_/Q _17158_/B _17159_/A _19232_/Q _11980_/A _12005_/S vssd1 vssd1 vccd1
+ vccd1 _12052_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11003_ _11003_/A vssd1 vssd1 vccd1 vccd1 _18276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19040_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15811_ _18888_/Q vssd1 vssd1 vccd1 vccd1 _16063_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_219_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16791_ _16741_/S _17783_/Q input14/X vssd1 vssd1 vccd1 vccd1 _16791_/X sky130_fd_sc_hd__and3b_1
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04837_ clkbuf_0__04837_/X vssd1 vssd1 vccd1 vccd1 _17008__356/A sky130_fd_sc_hd__clkbuf_16
X_18530_ _18530_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15742_ _15748_/A vssd1 vssd1 vccd1 vccd1 _15742_/X sky130_fd_sc_hd__buf_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12954_ _17965_/Q _17672_/Q _13022_/B vssd1 vssd1 vccd1 vccd1 _12955_/B sky130_fd_sc_hd__mux2_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07556_ clkbuf_0__07556_/X vssd1 vssd1 vccd1 vccd1 _13103_/A sky130_fd_sc_hd__clkbuf_16
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11905_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12076_/S sky130_fd_sc_hd__clkbuf_2
X_18461_ _19039_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _17977_/Q _17659_/Q _12891_/S vssd1 vssd1 vccd1 vccd1 _12886_/B sky130_fd_sc_hd__mux2_1
XFILLER_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _19174_/Q _19166_/Q _19198_/Q _18333_/Q _14591_/X _14592_/X vssd1 vssd1 vccd1
+ vccd1 _14624_/X sky130_fd_sc_hd__mux4_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11834_/Y _13645_/B _13326_/B _11835_/X vssd1 vssd1 vccd1 vccd1 _11836_/Y
+ sky130_fd_sc_hd__o211ai_1
X_18392_ _18392_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17343_/A vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14555_ _18363_/Q _18315_/Q _18371_/Q _17704_/Q _14553_/X _14554_/X vssd1 vssd1 vccd1
+ vccd1 _14555_/X sky130_fd_sc_hd__mux4_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A vssd1 vssd1 vccd1 vccd1 _11767_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03981_ clkbuf_0__03981_/X vssd1 vssd1 vccd1 vccd1 _15750__1036/A sky130_fd_sc_hd__clkbuf_16
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15798__119 _15798__119/A vssd1 vssd1 vccd1 vccd1 _18791_/CLK sky130_fd_sc_hd__inv_2
XFILLER_186_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ _17813_/Q _13499_/X _13505_/Y vssd1 vssd1 vccd1 vccd1 _17813_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17274_ _17276_/A _17274_/B _17274_/C _17274_/D vssd1 vssd1 vccd1 vccd1 _17288_/D
+ sky130_fd_sc_hd__and4_1
X_10718_ _18402_/Q _10690_/X _10726_/S vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11698_ _18412_/Q _11694_/C _11697_/X vssd1 vssd1 vccd1 vccd1 _11698_/Y sky130_fd_sc_hd__a21oi_1
X_16091__204 _16091__204/A vssd1 vssd1 vccd1 vccd1 _18909_/CLK sky130_fd_sc_hd__inv_2
X_19013_ _19013_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
X_16225_ _16143_/X _16224_/X _16119_/X vssd1 vssd1 vccd1 vccd1 _16225_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14435__603 _14436__604/A vssd1 vssd1 vccd1 vccd1 _18238_/CLK sky130_fd_sc_hd__inv_2
X_13437_ _13457_/B vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10649_ _10649_/A vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _13368_/A vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13299_ _17759_/Q _13282_/X _13298_/Y vssd1 vssd1 vccd1 vccd1 _17759_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15038_ _15038_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03415_ clkbuf_0__03415_/X vssd1 vssd1 vccd1 vccd1 _14845__769/A sky130_fd_sc_hd__clkbuf_16
XFILLER_228_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16989_ _16836_/X _16982_/Y _16984_/Y _16986_/Y _16988_/Y vssd1 vssd1 vccd1 vccd1
+ _16989_/X sky130_fd_sc_hd__o32a_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ _18965_/Q _09486_/X _09536_/S vssd1 vssd1 vccd1 vccd1 _09531_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18728_ _18728_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09461_ _09444_/B _09461_/B _09477_/C vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__and3b_1
X_18659_ _19144_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _19068_/Q _08964_/X _09394_/S vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260__463 _14260__463/A vssd1 vssd1 vccd1 vccd1 _18098_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _09728_/A vssd1 vssd1 vccd1 vccd1 _18858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09659_ _09659_/A vssd1 vssd1 vccd1 vccd1 _18913_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12672_/B _12673_/A _12607_/X vssd1 vssd1 vccd1 vccd1 _12670_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _17547_/Q _09674_/A _11629_/S vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12343__403 _12344__404/A vssd1 vssd1 vccd1 vccd1 _17584_/CLK sky130_fd_sc_hd__inv_2
XFILLER_243_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ _11552_/A vssd1 vssd1 vccd1 vccd1 _17710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10503_ _10503_/A vssd1 vssd1 vccd1 vccd1 _18527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11483_ _09133_/X _18052_/Q _11485_/S vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16010_ _16010_/A vssd1 vssd1 vccd1 vccd1 _16010_/X sky130_fd_sc_hd__clkbuf_2
X_13222_ _13892_/A vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__buf_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10434_ _10434_/A vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13153_ _13135_/X _13150_/X _13152_/Y _16619_/A vssd1 vssd1 vccd1 vccd1 _17725_/D
+ sky130_fd_sc_hd__a211oi_1
X_10365_ _10365_/A vssd1 vssd1 vccd1 vccd1 _18588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12104_ _12104_/A vssd1 vssd1 vccd1 vccd1 _12104_/Y sky130_fd_sc_hd__clkinv_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _17693_/Q _12924_/A _12834_/X _17688_/Q _13083_/X vssd1 vssd1 vccd1 vccd1
+ _13087_/C sky130_fd_sc_hd__o221a_1
X_17961_ _19039_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _18615_/Q _10180_/X _10302_/S vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12035_ _11936_/X _11920_/X _12067_/S vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15419__916 _15419__916/A vssd1 vssd1 vccd1 vccd1 _18603_/CLK sky130_fd_sc_hd__inv_2
X_16912_ _16819_/X _16905_/Y _16907_/Y _16909_/Y _16911_/Y vssd1 vssd1 vccd1 vccd1
+ _16912_/X sky130_fd_sc_hd__o32a_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17892_ _19109_/CLK _17892_/D vssd1 vssd1 vccd1 vccd1 _17892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14430__599 _14430__599/A vssd1 vssd1 vccd1 vccd1 _18234_/CLK sky130_fd_sc_hd__inv_2
XFILLER_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16843_ _18148_/Q _18140_/Q _18132_/Q _18276_/Q _16803_/X _16804_/X vssd1 vssd1 vccd1
+ vccd1 _16843_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ _16765_/X _16771_/Y _16773_/Y _14081_/A _16762_/X vssd1 vssd1 vccd1 vccd1
+ _16775_/B sky130_fd_sc_hd__o32a_1
XFILLER_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _17975_/Q _13968_/X _13985_/Y vssd1 vssd1 vccd1 vccd1 _17975_/D sky130_fd_sc_hd__o21a_1
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18513_ _18513_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03162_ _14349_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03162_/X sky130_fd_sc_hd__clkbuf_16
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _17657_/Q _13094_/B vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__xnor2_1
XFILLER_207_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03093_ _14158_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03093_/X sky130_fd_sc_hd__clkbuf_16
X_18444_ _18444_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12868_ _17982_/Q _17654_/Q _12944_/B vssd1 vssd1 vccd1 vccd1 _12869_/B sky130_fd_sc_hd__mux2_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14607_ _19049_/Q vssd1 vssd1 vccd1 vccd1 _14607_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11819_ _17910_/Q _11812_/X _11809_/Y input15/X _11796_/X vssd1 vssd1 vccd1 vccd1
+ _11819_/X sky130_fd_sc_hd__a221o_1
X_18375_ _18375_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
X_15587_ _18651_/Q _15597_/B vssd1 vssd1 vccd1 vccd1 _15587_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _17642_/Q _17993_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12800_/B sky130_fd_sc_hd__mux2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17326_ _17326_/A vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03964_ clkbuf_0__03964_/X vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_174_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15732__1021 _15735__1024/A vssd1 vssd1 vccd1 vccd1 _18738_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _17262_/C _17258_/C _17256_/Y vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__o21a_1
XFILLER_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16208_ _16204_/X _16207_/X _16248_/S vssd1 vssd1 vccd1 vccd1 _16208_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17188_ _17186_/B _17186_/C _17186_/D _19239_/Q vssd1 vssd1 vccd1 vccd1 _17189_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _18594_/Q _18610_/Q _18736_/Q _18517_/Q _16106_/X _16138_/X vssd1 vssd1 vccd1
+ vccd1 _16140_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _09691_/A vssd1 vssd1 vccd1 vccd1 _08961_/X sky130_fd_sc_hd__buf_2
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08892_ _08907_/S vssd1 vssd1 vccd1 vccd1 _08901_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04378_ clkbuf_0__04378_/X vssd1 vssd1 vccd1 vccd1 _16541__253/A sky130_fd_sc_hd__clkbuf_16
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17035__28 _17036__29/A vssd1 vssd1 vccd1 vccd1 _19177_/CLK sky130_fd_sc_hd__inv_2
X_09513_ _09513_/A vssd1 vssd1 vccd1 vccd1 _19003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__and2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _19075_/Q _09116_/X _09375_/S vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16666__301 _16666__301/A vssd1 vssd1 vccd1 vccd1 _19075_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03151_ clkbuf_0__03151_/X vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_193_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10150_ _10150_/A vssd1 vssd1 vccd1 vccd1 _18706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ _10081_/A vssd1 vssd1 vccd1 vccd1 _18733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03984_ clkbuf_0__03984_/X vssd1 vssd1 vccd1 vccd1 _15766__1049/A sky130_fd_sc_hd__clkbuf_16
XFILLER_88_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13840_ input57/X _13847_/B vssd1 vssd1 vccd1 vccd1 _13840_/X sky130_fd_sc_hd__and2_1
XFILLER_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102__409 _13102__409/A vssd1 vssd1 vccd1 vccd1 _17705_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13771_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13771_/X sky130_fd_sc_hd__clkbuf_2
X_10983_ _18283_/Q _09767_/X hold11/X vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15510_ _17838_/Q _15517_/B vssd1 vssd1 vccd1 vccd1 _15511_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12722_ _12727_/C _12727_/D _12718_/X vssd1 vssd1 vccd1 vccd1 _12723_/B sky130_fd_sc_hd__o21ai_1
XFILLER_243_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _16488_/X _16489_/Y _16469_/X vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15441_ _15441_/A vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__buf_1
X_12653_ _17604_/Q _12647_/X _12617_/X vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11604_/A vssd1 vssd1 vccd1 vccd1 _17572_/D sky130_fd_sc_hd__clkbuf_1
X_18160_ _18160_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15372_ _15368_/X _15369_/X _15370_/X _15371_/X _15281_/X _15222_/X vssd1 vssd1 vccd1
+ vccd1 _15372_/X sky130_fd_sc_hd__mux4_1
X_12584_ _12459_/X _12453_/X _12457_/X _12583_/X _12569_/S _12502_/A vssd1 vssd1 vccd1
+ vccd1 _12584_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03418_ clkbuf_0__03418_/X vssd1 vssd1 vccd1 vccd1 _14862__783/A sky130_fd_sc_hd__clkbuf_16
XFILLER_129_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _17239_/A vssd1 vssd1 vccd1 vccd1 _17112_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11535_ _08871_/X _17717_/Q _11539_/S vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__mux2_1
X_18091_ _18091_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11466_ _11466_/A vssd1 vssd1 vccd1 vccd1 _18060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13205_ input65/X _13446_/B vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__nand2_1
X_10417_ _10417_/A _10417_/B vssd1 vssd1 vccd1 vccd1 _18565_/D sky130_fd_sc_hd__nor2_1
X_11397_ _11397_/A vssd1 vssd1 vccd1 vccd1 _18117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14185_ _18065_/Q _14186_/D _14184_/Y vssd1 vssd1 vccd1 vccd1 _18065_/D sky130_fd_sc_hd__o21a_1
XFILLER_87_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13136_ _14243_/C vssd1 vssd1 vccd1 vccd1 _13216_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _18474_/Q vssd1 vssd1 vccd1 vccd1 _10348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_225_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18993_ _18993_/CLK _18993_/D vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_140_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _17939_/Q _17699_/Q _13070_/S vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__mux2_1
X_17944_ _17945_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _10279_/A vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ _12115_/S vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17875_ _17878_/CLK _17875_/D vssd1 vssd1 vccd1 vccd1 _17875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16826_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16927_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1__f__04163_ clkbuf_0__04163_/X vssd1 vssd1 vccd1 vccd1 _16071__187/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16757_ _16775_/A _16757_/B vssd1 vssd1 vccd1 vccd1 _19129_/D sky130_fd_sc_hd__nor2_1
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13969_ _13717_/A _13968_/X _13920_/X vssd1 vssd1 vccd1 vccd1 _13969_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_62_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03145_ _14262_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03145_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16688_ _13387_/B _16688_/B vssd1 vssd1 vccd1 vccd1 _16737_/B sky130_fd_sc_hd__and2b_1
X_14890__805 _14892__807/A vssd1 vssd1 vccd1 vccd1 _18450_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18427_ _18427_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
X_15639_ _16059_/A _15641_/B vssd1 vssd1 vccd1 vccd1 _18666_/D sky130_fd_sc_hd__nor2_1
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _19175_/Q _09104_/X _09160_/S vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__mux2_1
X_18358_ _18358_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17309_ _17309_/A vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09091_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _10695_/A sky130_fd_sc_hd__buf_2
X_18289_ _18289_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03978_ _15730_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03978_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_134_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14372__553 _14373__554/A vssd1 vssd1 vccd1 vccd1 _18188_/CLK sky130_fd_sc_hd__inv_2
XFILLER_157_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09993_ _09993_/A vssd1 vssd1 vccd1 vccd1 _18767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _09674_/A vssd1 vssd1 vccd1 vccd1 _08944_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16661__297 _16663__299/A vssd1 vssd1 vccd1 vccd1 _19071_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__08198_ clkbuf_0__08198_/X vssd1 vssd1 vccd1 vccd1 _13106__412/A sky130_fd_sc_hd__clkbuf_16
X_08875_ _19312_/Q _08874_/X _08878_/S vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09427_ _09427_/A vssd1 vssd1 vccd1 vccd1 _19053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791__725 _14793__727/A vssd1 vssd1 vccd1 vccd1 _18368_/CLK sky130_fd_sc_hd__inv_2
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _09770_/A _09358_/B _09770_/B vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__or3_4
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09289_ _19117_/Q _08952_/X _09293_/S vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__mux2_1
X_12227__373 _12228__374/A vssd1 vssd1 vccd1 vccd1 _17537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11320_ _11320_/A vssd1 vssd1 vccd1 vccd1 _18147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ _11156_/X _18174_/Q _11251_/S vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ hold6/A vssd1 vssd1 vccd1 vccd1 _10211_/S sky130_fd_sc_hd__clkbuf_2
X_14273__473 _14274__474/A vssd1 vssd1 vccd1 vccd1 _18108_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ _11162_/X _18204_/Q _11184_/S vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10133_ _10132_/X _18712_/Q _10136_/S vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _18867_/Q _15991_/B vssd1 vssd1 vccd1 vccd1 _15992_/B sky130_fd_sc_hd__nor2_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ _17856_/Q _14948_/A vssd1 vssd1 vccd1 vccd1 _14942_/C sky130_fd_sc_hd__nand2_1
XFILLER_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10064_ _18738_/Q _10063_/X _10064_/S vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__mux2_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03967_ clkbuf_0__03967_/X vssd1 vssd1 vccd1 vccd1 _15679__979/A sky130_fd_sc_hd__clkbuf_16
X_15731__1020 _15731__1020/A vssd1 vssd1 vccd1 vccd1 _18737_/CLK sky130_fd_sc_hd__inv_2
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ _17969_/CLK _17660_/D vssd1 vssd1 vccd1 vccd1 _17660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16611_ _19034_/Q _16608_/B _16610_/Y vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13823_ _19147_/Q input63/X _13828_/B vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__and3_1
X_17591_ _18010_/CLK _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_106 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_117 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19330_ _19336_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_128 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ _17895_/Q _13743_/B _13752_/Y _13753_/X vssd1 vssd1 vccd1 vccd1 _17895_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_139 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ _10966_/A vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12705_ _12706_/B _12703_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _17619_/D sky130_fd_sc_hd__a21oi_1
X_19261_ _19261_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16473_ _18977_/Q _16473_/B vssd1 vssd1 vccd1 vccd1 _16482_/C sky130_fd_sc_hd__and2_1
X_13685_ _17871_/Q _13682_/X _13684_/Y vssd1 vssd1 vccd1 vccd1 _17871_/D sky130_fd_sc_hd__o21a_1
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ _10897_/A vssd1 vssd1 vccd1 vccd1 _18320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18212_ _18212_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12636_ _12634_/X _12636_/B _12695_/A vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__and3b_1
Xclkbuf_1_1__f__04850_ clkbuf_0__04850_/X vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__clkbuf_16
X_19192_ _19192_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18143_ _18143_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03801_ clkbuf_0__03801_/X vssd1 vssd1 vccd1 vccd1 _15428__924/A sky130_fd_sc_hd__clkbuf_16
XFILLER_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15355_ _15351_/X _15352_/X _15353_/X _15354_/X _15281_/X _09600_/X vssd1 vssd1 vccd1
+ vccd1 _15355_/X sky130_fd_sc_hd__mux4_1
X_12567_ _12463_/X _12464_/X _12567_/S vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__mux2_1
XFILLER_156_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__07169_ clkbuf_0__07169_/X vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_89_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _14318_/A vssd1 vssd1 vccd1 vccd1 _14306_/X sky130_fd_sc_hd__buf_1
XFILLER_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11518_ _11518_/A vssd1 vssd1 vccd1 vccd1 _18037_/D sky130_fd_sc_hd__clkbuf_1
X_18074_ _18870_/CLK _18074_/D vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
X_15286_ _09614_/A _15284_/Y _15285_/X vssd1 vssd1 vccd1 vccd1 _15286_/Y sky130_fd_sc_hd__a21oi_1
X_12498_ _12492_/X _12497_/X _12515_/A vssd1 vssd1 vccd1 vccd1 _12763_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17025_ _17037_/A vssd1 vssd1 vccd1 vccd1 _17025_/X sky130_fd_sc_hd__buf_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ _18481_/Q vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11449_ _11449_/A vssd1 vssd1 vccd1 vccd1 _18094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03594_ clkbuf_0__03594_/X vssd1 vssd1 vccd1 vccd1 _15130__844/A sky130_fd_sc_hd__clkbuf_16
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14099_ _14099_/A vssd1 vssd1 vccd1 vccd1 _14099_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _18987_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653__958 _15654__959/A vssd1 vssd1 vccd1 vccd1 _18675_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _19132_/CLK _17927_/D vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17858_ _17935_/CLK _17858_/D vssd1 vssd1 vccd1 vccd1 _17858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ _16893_/A vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__buf_2
XFILLER_187_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17789_ _19132_/CLK _17789_/D vssd1 vssd1 vccd1 vccd1 _17789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14855__777 _14857__779/A vssd1 vssd1 vccd1 vccd1 _18422_/CLK sky130_fd_sc_hd__inv_2
X_09212_ _09212_/A vssd1 vssd1 vccd1 vccd1 _19153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09143_ _19181_/Q _09142_/X _09146_/S vssd1 vssd1 vccd1 vccd1 _09144_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ _09074_/A vssd1 vssd1 vccd1 vccd1 _19198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _10528_/B _10030_/B vssd1 vssd1 vccd1 vccd1 _09992_/S sky130_fd_sc_hd__nor2_2
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08927_ _08927_/A vssd1 vssd1 vccd1 vccd1 _19296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ input74/X vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__buf_6
XFILLER_245_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08789_ _18885_/Q vssd1 vssd1 vccd1 vccd1 _08789_/X sky130_fd_sc_hd__buf_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ _10820_/A vssd1 vssd1 vccd1 vccd1 _18361_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10751_ _10751_/A vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13470_ _13529_/A vssd1 vssd1 vccd1 vccd1 _16059_/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_27_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _19339_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10682_ _18416_/Q _09732_/X _10682_/S vssd1 vssd1 vccd1 vccd1 _10683_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14379__559 _14379__559/A vssd1 vssd1 vccd1 vccd1 _18194_/CLK sky130_fd_sc_hd__inv_2
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14756__697 _14757__698/A vssd1 vssd1 vccd1 vccd1 _18340_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _17621_/Q _12717_/B _12717_/A _17624_/Q _12555_/A _12429_/S vssd1 vssd1 vccd1
+ vccd1 _12421_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12352_ _18012_/Q vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04166_ clkbuf_0__04166_/X vssd1 vssd1 vccd1 vccd1 _16091__204/A sky130_fd_sc_hd__clkbuf_16
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11303_ _11457_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11319_/S sky130_fd_sc_hd__or2_2
X_15071_ _16059_/A _15177_/A vssd1 vssd1 vccd1 vccd1 _18478_/D sky130_fd_sc_hd__nor2_1
X_12283_ _12283_/A vssd1 vssd1 vccd1 vccd1 _17559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15749__1035 _15750__1036/A vssd1 vssd1 vccd1 vccd1 _18752_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _17987_/Q _14011_/X _14021_/Y vssd1 vssd1 vccd1 vccd1 _17987_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11234_ _11234_/A vssd1 vssd1 vccd1 vccd1 _18182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18830_ _18830_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _11344_/A vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__buf_2
XFILLER_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16679__311 _16680__312/A vssd1 vssd1 vccd1 vccd1 _19085_/CLK sky130_fd_sc_hd__inv_2
XFILLER_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _10116_/A vssd1 vssd1 vccd1 vccd1 _18718_/D sky130_fd_sc_hd__clkbuf_1
X_18761_ _18761_/CLK _18761_/D vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_1
X_11096_ _09039_/X _18239_/Q _11098_/S vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__mux2_1
X_15973_ _18864_/Q _15973_/B vssd1 vssd1 vccd1 vccd1 _15985_/C sky130_fd_sc_hd__and2_1
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ _14924_/A vssd1 vssd1 vccd1 vccd1 _14964_/A sky130_fd_sc_hd__inv_2
X_10047_ _10047_/A vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__clkbuf_1
X_17712_ _17712_/CLK _17712_/D vssd1 vssd1 vccd1 vccd1 _17712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18692_ _18692_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__05080_ _17403_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__05080_/X sky130_fd_sc_hd__clkbuf_16
X_17643_ _19246_/CLK _17643_/D vssd1 vssd1 vccd1 vccd1 _17643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ _13407_/X _13802_/X _13805_/X vssd1 vssd1 vccd1 vccd1 _13806_/Y sky130_fd_sc_hd__a21oi_1
X_17574_ _17574_/CLK _17574_/D vssd1 vssd1 vccd1 vccd1 _17574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11998_ _19261_/Q vssd1 vssd1 vccd1 vccd1 _17274_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14323__514 _14323__514/A vssd1 vssd1 vccd1 vccd1 _18149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19313_ _19313_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_16525_ _16525_/A vssd1 vssd1 vccd1 vccd1 _18990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ _14069_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13757_/B sky130_fd_sc_hd__or2_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10949_ hold8/X _11529_/B vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__or2_1
XFILLER_220_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19244_ _19247_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_1
X_16456_ _16454_/X _16455_/Y _16480_/A vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__a21oi_1
XFILLER_176_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13668_ _17865_/Q _13659_/X _13667_/Y vssd1 vssd1 vccd1 vccd1 _17865_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12619_ _12622_/C _12619_/B vssd1 vssd1 vccd1 vccd1 _17594_/D sky130_fd_sc_hd__nor2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115__419 _13115__419/A vssd1 vssd1 vccd1 vccd1 _17715_/CLK sky130_fd_sc_hd__inv_2
X_19175_ _19175_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_1
X_16387_ _17800_/Q _16393_/B _17799_/Q vssd1 vssd1 vccd1 vccd1 _16389_/C sky130_fd_sc_hd__o21ai_1
X_13599_ _13599_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13611_/S sky130_fd_sc_hd__nor2_1
XFILLER_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18126_ _18126_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15338_ _15334_/X _15335_/X _15336_/X _15337_/X _09600_/A _09625_/X vssd1 vssd1 vccd1
+ vccd1 _15338_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18057_ _18057_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15269_ _18570_/Q _15207_/X _15242_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _18570_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09830_ _09679_/X _18818_/Q _09836_/S vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09761_ _18882_/Q vssd1 vssd1 vccd1 vccd1 _09761_/X sky130_fd_sc_hd__buf_2
X_18959_ _18959_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15888__178 _15889__179/A vssd1 vssd1 vccd1 vccd1 _18854_/CLK sky130_fd_sc_hd__inv_2
X_09692_ _09691_/X _18900_/Q _09698_/S vssd1 vssd1 vccd1 vccd1 _09693_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09126_ _09126_/A vssd1 vssd1 vccd1 vccd1 _19187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16075__190 _16077__192/A vssd1 vssd1 vccd1 vccd1 _18895_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _09057_/A vssd1 vssd1 vccd1 vccd1 _19204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09959_ _10129_/A vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__buf_2
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04853_ clkbuf_0__04853_/X vssd1 vssd1 vccd1 vccd1 _17297__74/A sky130_fd_sc_hd__clkbuf_16
XFILLER_44_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12970_ _12970_/A vssd1 vssd1 vccd1 vccd1 _17676_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03804_ clkbuf_0__03804_/X vssd1 vssd1 vccd1 vccd1 _15444__937/A sky130_fd_sc_hd__clkbuf_16
XFILLER_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11921_ _19232_/Q _19233_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__mux2_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14734_/A vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11852_ _11852_/A vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10803_ _18990_/Q vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14571_ _14734_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14571_/Y sky130_fd_sc_hd__nor2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _13352_/B vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__buf_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13522_ _13523_/A vssd1 vssd1 vccd1 vccd1 _13522_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__03597_ clkbuf_0__03597_/X vssd1 vssd1 vccd1 vccd1 _15147__858/A sky130_fd_sc_hd__clkbuf_16
XFILLER_242_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17290_ _17290_/A vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10734_ _10851_/A hold13/A vssd1 vssd1 vccd1 vccd1 _10750_/S sky130_fd_sc_hd__nor2_2
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16241_ _18442_/Q _18692_/Q _18700_/Q _18708_/Q _16198_/X _16172_/X vssd1 vssd1 vccd1
+ vccd1 _16242_/B sky130_fd_sc_hd__mux4_2
X_13453_ _17799_/Q _13457_/B vssd1 vssd1 vccd1 vccd1 _13453_/Y sky130_fd_sc_hd__nor2_1
X_10665_ _10665_/A vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12404_ _12398_/X _12403_/X _12448_/A vssd1 vssd1 vccd1 vccd1 _12405_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16172_ _16172_/A vssd1 vssd1 vccd1 vccd1 _16172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13384_ _13599_/A vssd1 vssd1 vccd1 vccd1 _13769_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10596_ _09047_/X _18486_/Q hold19/X vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03600_ _15156_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03600_/X sky130_fd_sc_hd__clkbuf_16
X_15054_ _14904_/A _14978_/X _15048_/Y _15053_/X _14894_/Y vssd1 vssd1 vccd1 vccd1
+ _18469_/D sky130_fd_sc_hd__o311a_1
XFILLER_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ _12266_/A vssd1 vssd1 vccd1 vccd1 _17554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14005_/X sky130_fd_sc_hd__clkbuf_2
X_11217_ _11217_/A vssd1 vssd1 vccd1 vccd1 _18189_/D sky130_fd_sc_hd__clkbuf_1
X_12197_ _17517_/Q _17490_/B vssd1 vssd1 vccd1 vccd1 _12198_/D sky130_fd_sc_hd__xor2_1
XFILLER_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput81 _11773_/X vssd1 vssd1 vccd1 vccd1 flash_io1_read sky130_fd_sc_hd__buf_2
Xoutput92 _11872_/X vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__buf_2
X_18813_ _18813_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11148_ _11147_/X _18217_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _11149_/A sky130_fd_sc_hd__mux2_1
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806__738 _14806__738/A vssd1 vssd1 vccd1 vccd1 _18381_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18744_ _18744_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _09043_/X _18246_/Q _11079_/S vssd1 vssd1 vccd1 vccd1 _11080_/A sky130_fd_sc_hd__mux2_1
X_15956_ _15989_/A vssd1 vssd1 vccd1 vccd1 _15986_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_237_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14907_ _14907_/A vssd1 vssd1 vccd1 vccd1 _14936_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18675_ _18675_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17626_ _17629_/CLK _17626_/D vssd1 vssd1 vccd1 vccd1 _17626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04014_ _15874_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04014_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17557_ _18027_/CLK _17557_/D vssd1 vssd1 vccd1 vccd1 _17557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _16514_/A _16511_/B _16507_/X vssd1 vssd1 vccd1 vccd1 _16508_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_225_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17488_ _19325_/Q _12187_/A _12185_/X _19339_/Q vssd1 vssd1 vccd1 vccd1 _17494_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_177_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19227_ _19252_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16439_ _16467_/A _16445_/B _16439_/C vssd1 vssd1 vccd1 vccd1 _16439_/X sky130_fd_sc_hd__or3_1
XFILLER_108_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19158_ _19158_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04847_ _17056_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04847_/X sky130_fd_sc_hd__clkbuf_16
X_18109_ _18109_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ _19089_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _09813_/A vssd1 vssd1 vccd1 vccd1 _18826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09744_ _18887_/Q vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_246_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09675_ _11637_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09698_/S sky130_fd_sc_hd__or2_2
XFILLER_227_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15412__911 _15413__912/A vssd1 vssd1 vccd1 vccd1 _18598_/CLK sky130_fd_sc_hd__inv_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15666__968 _15667__969/A vssd1 vssd1 vccd1 vccd1 _18685_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ _10129_/X _18550_/Q _10454_/S vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _19190_/Q _09108_/X _09117_/S vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ _10381_/A vssd1 vssd1 vccd1 vccd1 _18581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _17487_/B vssd1 vssd1 vccd1 vccd1 _12121_/D sky130_fd_sc_hd__inv_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _19225_/Q _19226_/Q _17142_/A _11978_/X _11980_/X _11981_/X vssd1 vssd1 vccd1
+ vccd1 _12051_/X sky130_fd_sc_hd__mux4_2
X_17500__7 _17501__8/A vssd1 vssd1 vccd1 vccd1 _19342_/CLK sky130_fd_sc_hd__inv_2
XFILLER_132_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11002_ _18276_/Q _09142_/X _11004_/S vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15810_ _17827_/Q _09016_/X _13681_/A _15641_/B vssd1 vssd1 vccd1 vccd1 _18800_/D
+ sky130_fd_sc_hd__a211oi_1
X_16790_ _16795_/A _16790_/B vssd1 vssd1 vccd1 vccd1 _19135_/D sky130_fd_sc_hd__nor2_1
XFILLER_219_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04836_ clkbuf_0__04836_/X vssd1 vssd1 vccd1 vccd1 _17005__354/A sky130_fd_sc_hd__clkbuf_16
X_12953_ _12953_/A vssd1 vssd1 vccd1 vccd1 _17671_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07555_ clkbuf_0__07555_/X vssd1 vssd1 vccd1 vccd1 _12325__389/A sky130_fd_sc_hd__clkbuf_16
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ _17779_/Q vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_opt_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19261_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18460_ _18462_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12884_/A vssd1 vssd1 vccd1 vccd1 _17658_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14623_ _14623_/A vssd1 vssd1 vccd1 vccd1 _14623_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _13278_/B _17722_/Q input19/X vssd1 vssd1 vccd1 vccd1 _11835_/X sky130_fd_sc_hd__or3b_4
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18391_ _18391_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17340_/X _17342_/B vssd1 vssd1 vccd1 vccd1 _17343_/A sky130_fd_sc_hd__and2b_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14554_ _14627_/A vssd1 vssd1 vccd1 vccd1 _14554_/X sky130_fd_sc_hd__buf_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _17865_/Q _17669_/Q _18002_/Q vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__mux2_2
Xclkbuf_1_1__f__03980_ clkbuf_0__03980_/X vssd1 vssd1 vccd1 vccd1 _15747__1034/A sky130_fd_sc_hd__clkbuf_16
XFILLER_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13231_/X _13500_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _13505_/Y sky130_fd_sc_hd__a21oi_1
X_17273_ _17273_/A vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10717_ _10732_/S vssd1 vssd1 vccd1 vccd1 _10726_/S sky130_fd_sc_hd__clkbuf_2
X_11697_ _13951_/A vssd1 vssd1 vccd1 vccd1 _11697_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_201_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19012_ _19012_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
X_16224_ _18449_/Q _19087_/Q _19124_/Q _18433_/Q _16144_/X _16108_/X vssd1 vssd1 vccd1
+ vccd1 _16224_/X sky130_fd_sc_hd__mux4_2
X_13436_ _13447_/S vssd1 vssd1 vccd1 vccd1 _13457_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10648_ _09271_/X _18432_/Q _10648_/S vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14812__742 _14813__743/A vssd1 vssd1 vccd1 vccd1 _18385_/CLK sky130_fd_sc_hd__inv_2
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16155_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16155_/X sky130_fd_sc_hd__buf_2
X_13367_ _16715_/B _13367_/B vssd1 vssd1 vccd1 vccd1 _17777_/D sky130_fd_sc_hd__nor2_1
XFILLER_154_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10579_ _10579_/A vssd1 vssd1 vccd1 vccd1 _18493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15106_/X sky130_fd_sc_hd__buf_1
X_12318_ _16578_/A _12318_/B _12318_/C vssd1 vssd1 vccd1 vccd1 _17564_/D sky130_fd_sc_hd__nor3_1
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16086_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16086_/X sky130_fd_sc_hd__buf_1
X_13298_ _13244_/X _13288_/X _13293_/X vssd1 vssd1 vccd1 vccd1 _13298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ _18466_/Q _15043_/C vssd1 vssd1 vccd1 vccd1 _15042_/B sky130_fd_sc_hd__and2_1
XFILLER_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12249_ _17550_/Q _18027_/Q _12318_/B vssd1 vssd1 vccd1 vccd1 _12250_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03414_ clkbuf_0__03414_/X vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16988_ _09859_/A _16987_/X _16902_/A vssd1 vssd1 vccd1 vccd1 _16988_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17047__37 _17049__39/A vssd1 vssd1 vccd1 vccd1 _19186_/CLK sky130_fd_sc_hd__inv_2
X_16323__221 _16323__221/A vssd1 vssd1 vccd1 vccd1 _18937_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18727_ _18727_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _18869_/Q _15940_/B vssd1 vssd1 vccd1 vccd1 _15939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09460_ _19013_/Q _16559_/C _09459_/X vssd1 vssd1 vccd1 vccd1 _09461_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18658_ _18670_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17609_ _17609_/CLK _17609_/D vssd1 vssd1 vccd1 vccd1 _17609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09391_ _09391_/A vssd1 vssd1 vccd1 vccd1 _19069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _18589_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14336__524 _14336__524/A vssd1 vssd1 vccd1 vccd1 _18159_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15145__856 _15148__859/A vssd1 vssd1 vccd1 vccd1 _18532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221__368 _12222__369/A vssd1 vssd1 vccd1 vccd1 _17532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_161_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16625__268 _16626__269/A vssd1 vssd1 vccd1 vccd1 _19042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ _18858_/Q _09726_/X _09733_/S vssd1 vssd1 vccd1 vccd1 _09728_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09658_ _18913_/Q _09223_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _18939_/Q _09492_/X _09591_/S vssd1 vssd1 vccd1 vccd1 _09590_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11620_ _11635_/S vssd1 vssd1 vccd1 vccd1 _11629_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14497__653 _14498__654/A vssd1 vssd1 vccd1 vccd1 _18288_/CLK sky130_fd_sc_hd__inv_2
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ _17710_/Q _10892_/X _11557_/S vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ _10126_/X _18527_/Q _10502_/S vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__mux2_1
X_11482_ _11482_/A vssd1 vssd1 vccd1 vccd1 _18053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13221_ _13434_/A vssd1 vssd1 vccd1 vccd1 _13717_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10433_ _10424_/C _10433_/B _10433_/C vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__and3b_1
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13152_ _17725_/Q _14134_/B vssd1 vssd1 vccd1 vccd1 _13152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10364_ _18588_/Q _09732_/X _10364_/S vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12103_/A vssd1 vssd1 vccd1 vccd1 _12103_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11881__364 _11881__364/A vssd1 vssd1 vccd1 vccd1 _17511_/CLK sky130_fd_sc_hd__inv_2
X_13083_ _17699_/Q _12845_/A _12838_/A _17702_/Q _13082_/Y vssd1 vssd1 vccd1 vccd1
+ _13083_/X sky130_fd_sc_hd__o221a_1
XFILLER_174_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17960_ _17963_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10295_ _10295_/A vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12034_ _12034_/A _12034_/B vssd1 vssd1 vccd1 vccd1 _12034_/Y sky130_fd_sc_hd__nand2_1
X_16911_ _09868_/X _16910_/X _16886_/X vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_238_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17891_ _19109_/CLK _17891_/D vssd1 vssd1 vccd1 vccd1 _17891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16842_ _18116_/Q _18108_/Q _18100_/Q _18092_/Q _16799_/X _16801_/X vssd1 vssd1 vccd1
+ vccd1 _16842_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13985_ _13792_/X _13973_/A _13978_/X vssd1 vssd1 vccd1 vccd1 _13985_/Y sky130_fd_sc_hd__a21oi_1
X_16773_ _16783_/A _16773_/B vssd1 vssd1 vccd1 vccd1 _16773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03161_ _14343_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03161_/X sky130_fd_sc_hd__clkbuf_16
X_18512_ _18512_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_1
X_12936_ _17656_/Q _12932_/X _12850_/A _17653_/Q vssd1 vssd1 vccd1 vccd1 _12942_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_15724_ _15730_/A vssd1 vssd1 vccd1 vccd1 _15724_/X sky130_fd_sc_hd__buf_1
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03092_ _14157_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03092_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18443_ _18443_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _12867_/A vssd1 vssd1 vccd1 vccd1 _17653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15655_ _15655_/A vssd1 vssd1 vccd1 vccd1 _15655_/X sky130_fd_sc_hd__buf_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _17930_/Q _11815_/X _11816_/X _11817_/X vssd1 vssd1 vccd1 vccd1 _11818_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14606_ _19050_/Q vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15586_ _15611_/A _15586_/B _15595_/C vssd1 vssd1 vccd1 vccd1 _15586_/X sky130_fd_sc_hd__or3_1
X_18374_ _18374_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_1
X_12798_ _12798_/A vssd1 vssd1 vccd1 vccd1 _17641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17323_/X _17325_/B vssd1 vssd1 vccd1 vccd1 _17326_/A sky130_fd_sc_hd__and2b_1
X_11749_ _11749_/A vssd1 vssd1 vccd1 vccd1 _11749_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_239_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14398__573 _14399__574/A vssd1 vssd1 vccd1 vccd1 _18208_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03963_ clkbuf_0__03963_/X vssd1 vssd1 vccd1 vccd1 _15660__964/A sky130_fd_sc_hd__clkbuf_16
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17256_ _17262_/C _17258_/C _17112_/B vssd1 vssd1 vccd1 vccd1 _17256_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468_ _14474_/A vssd1 vssd1 vccd1 vccd1 _14468_/X sky130_fd_sc_hd__buf_1
XFILLER_88_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13419_ _17791_/Q _13393_/X _13418_/Y vssd1 vssd1 vccd1 vccd1 _17791_/D sky130_fd_sc_hd__o21a_1
X_16207_ _18714_/Q _18722_/Q _18730_/Q _18495_/Q _16205_/X _16206_/X vssd1 vssd1 vccd1
+ vccd1 _16207_/X sky130_fd_sc_hd__mux4_2
X_17187_ _17203_/C vssd1 vssd1 vccd1 vccd1 _17195_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16138_ _16138_/A vssd1 vssd1 vccd1 vccd1 _16138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08960_ _08960_/A vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16544__255 _16547__258/A vssd1 vssd1 vccd1 vccd1 _19001_/CLK sky130_fd_sc_hd__inv_2
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08891_ _08945_/B _10967_/A vssd1 vssd1 vccd1 vccd1 _08907_/S sky130_fd_sc_hd__nor2_2
XFILLER_124_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04377_ clkbuf_0__04377_/X vssd1 vssd1 vccd1 vccd1 _16355__246/A sky130_fd_sc_hd__clkbuf_16
XFILLER_97_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14743__688 _14744__689/A vssd1 vssd1 vccd1 vccd1 _18331_/CLK sky130_fd_sc_hd__inv_2
XFILLER_237_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09512_ _19003_/Q _09486_/X _09518_/S vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09443_/A _19013_/Q _16559_/C vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__and3_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14819__748 _14820__749/A vssd1 vssd1 vccd1 vccd1 _18391_/CLK sky130_fd_sc_hd__inv_2
X_09374_ _09374_/A vssd1 vssd1 vccd1 vccd1 _19076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03150_ clkbuf_0__03150_/X vssd1 vssd1 vccd1 vccd1 _14290__487/A sky130_fd_sc_hd__clkbuf_16
XFILLER_123_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ _18733_/Q _10054_/X _10086_/S vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__mux2_1
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_0 _18064_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03983_ clkbuf_0__03983_/X vssd1 vssd1 vccd1 vccd1 _15758__1042/A sky130_fd_sc_hd__clkbuf_16
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10982_ _10982_/A vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12721_ _12727_/C _12727_/D vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__and2_1
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12652_ _12666_/C vssd1 vssd1 vccd1 vccd1 _12658_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_203_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11603_ _17572_/Q _10690_/A _11611_/S vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15371_ _18942_/Q _18905_/Q _18897_/Q _18851_/Q _15248_/X _15249_/X vssd1 vssd1 vccd1
+ vccd1 _15371_/X sky130_fd_sc_hd__mux4_1
X_12583_ _17630_/Q _12746_/B _12746_/A _17633_/Q _12555_/X _12556_/X vssd1 vssd1 vccd1
+ vccd1 _12583_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03417_ clkbuf_0__03417_/X vssd1 vssd1 vccd1 vccd1 _14857__779/A sky130_fd_sc_hd__clkbuf_16
XFILLER_157_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15087__810 _15089__812/A vssd1 vssd1 vccd1 vccd1 _18486_/CLK sky130_fd_sc_hd__inv_2
X_17110_ _17114_/A vssd1 vssd1 vccd1 vccd1 _17239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11534_ _11534_/A vssd1 vssd1 vccd1 vccd1 _17718_/D sky130_fd_sc_hd__clkbuf_1
X_18090_ _18922_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
X_15425__921 _15425__921/A vssd1 vssd1 vccd1 vccd1 _18608_/CLK sky130_fd_sc_hd__inv_2
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _11332_/X _18060_/Q _11467_/S vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__mux2_1
X_13204_ _13170_/X _16056_/A _13203_/Y _13187_/X vssd1 vssd1 vccd1 vccd1 _17734_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_183_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ _10405_/A _10405_/B _10407_/X vssd1 vssd1 vccd1 vccd1 _10417_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ _14184_/A _14249_/B vssd1 vssd1 vccd1 vccd1 _14184_/Y sky130_fd_sc_hd__nor2_1
X_11396_ _11338_/X _18117_/Q _11400_/S vssd1 vssd1 vccd1 vccd1 _11397_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13135_ _14136_/B vssd1 vssd1 vccd1 vccd1 _13135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10347_ _10347_/A vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18992_ _18996_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17943_ _17951_/CLK _17943_/D vssd1 vssd1 vccd1 vccd1 _17943_/Q sky130_fd_sc_hd__dfxtp_1
X_13066_ _13066_/A vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__clkbuf_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10278_ _18623_/Q _10180_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12017_ _11935_/X _11936_/X _12017_/S vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17874_ _17878_/CLK _17874_/D vssd1 vssd1 vccd1 vccd1 _17874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16825_ _16986_/A _16825_/B vssd1 vssd1 vccd1 vccd1 _16825_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__04162_ clkbuf_0__04162_/X vssd1 vssd1 vccd1 vccd1 _16092_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16756_ _13871_/A _16762_/A _16755_/Y _16687_/B vssd1 vssd1 vccd1 vccd1 _16757_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13968_ _13973_/A vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03144_ _14256_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03144_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12919_ _16690_/A vssd1 vssd1 vccd1 vccd1 _16620_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_207_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13899_ _13792_/X _13885_/A _13894_/X vssd1 vssd1 vccd1 vccd1 _13899_/Y sky130_fd_sc_hd__a21oi_1
X_16687_ _19109_/Q _16687_/B vssd1 vssd1 vccd1 vccd1 _16687_/X sky130_fd_sc_hd__and2_1
XFILLER_59_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _18426_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
X_15638_ _16058_/A _15638_/B vssd1 vssd1 vccd1 vccd1 _18665_/D sky130_fd_sc_hd__nor2_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040__32 _17042__34/A vssd1 vssd1 vccd1 vccd1 _19181_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _18357_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _15572_/B _15569_/B vssd1 vssd1 vccd1 vccd1 _15569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17308_ _17304_/X _17308_/B vssd1 vssd1 vccd1 vccd1 _17309_/A sky130_fd_sc_hd__and2b_1
X_09090_ _09090_/A vssd1 vssd1 vccd1 vccd1 _19195_/D sky130_fd_sc_hd__clkbuf_1
X_18288_ _18288_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17239_ _17239_/A vssd1 vssd1 vccd1 vccd1 _17265_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__03977_ _15724_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03977_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09992_ _18767_/Q _09967_/X _09992_/S vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08943_ _08943_/A vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__04529_ _16550_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04529_/X sky130_fd_sc_hd__clkbuf_16
X_14448__614 _14448__614/A vssd1 vssd1 vccd1 vccd1 _18249_/CLK sky130_fd_sc_hd__inv_2
XFILLER_233_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08874_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _08874_/X sky130_fd_sc_hd__buf_6
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ _08933_/X _19053_/Q _09430_/S vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09357_ _09357_/A vssd1 vssd1 vccd1 vccd1 _19083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ _09288_/A vssd1 vssd1 vccd1 vccd1 _19118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11250_/A vssd1 vssd1 vccd1 vccd1 _18175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _11655_/A hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__nor2_2
XFILLER_107_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11181_ _11181_/A vssd1 vssd1 vccd1 vccd1 _18205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10132_ _10132_/A vssd1 vssd1 vccd1 vccd1 _10132_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ _14940_/A _17858_/Q _17857_/Q vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__or3_1
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10063_ _10126_/A vssd1 vssd1 vccd1 vccd1 _10063_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03966_ clkbuf_0__03966_/X vssd1 vssd1 vccd1 vccd1 _15671__972/A sky130_fd_sc_hd__clkbuf_16
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ _14883_/A vssd1 vssd1 vccd1 vccd1 _14871_/X sky130_fd_sc_hd__buf_1
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15158__866 _15158__866/A vssd1 vssd1 vccd1 vccd1 _18542_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16610_ _19034_/Q _16608_/B _14184_/A vssd1 vssd1 vccd1 vccd1 _16610_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ _17917_/Q _13820_/Y _13821_/X _13753_/X vssd1 vssd1 vccd1 vccd1 _17917_/D
+ sky130_fd_sc_hd__a211o_1
X_17590_ _18010_/CLK _17590_/D vssd1 vssd1 vccd1 vccd1 _17590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_107 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_118 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ _13841_/A vssd1 vssd1 vccd1 vccd1 _13753_/X sky130_fd_sc_hd__buf_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_129 _19387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10965_ _08886_/X _18291_/Q hold9/X vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ _12706_/B _12703_/A _12607_/X vssd1 vssd1 vccd1 vccd1 _12704_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19260_ _19266_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13684_ _13394_/X _13683_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _13684_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16472_ _18977_/Q _16473_/B vssd1 vssd1 vccd1 vccd1 _16474_/B sky130_fd_sc_hd__nor2_1
X_10896_ _18320_/Q _10895_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10897_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18211_ _18211_/CLK _18211_/D vssd1 vssd1 vccd1 vccd1 _18211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ _12638_/B _12641_/D vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__or2_1
X_15423_ _15429_/A vssd1 vssd1 vccd1 vccd1 _15423_/X sky130_fd_sc_hd__buf_1
XFILLER_176_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19191_ _19191_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18142_ _18142_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03800_ clkbuf_0__03800_/X vssd1 vssd1 vccd1 vccd1 _15419__916/A sky130_fd_sc_hd__clkbuf_16
X_15354_ _18941_/Q _18904_/Q _18896_/Q _18850_/Q _15248_/X _15249_/X vssd1 vssd1 vccd1
+ vccd1 _15354_/X sky130_fd_sc_hd__mux4_1
X_12566_ _12465_/X _12565_/X _12466_/X _12519_/X _12407_/A _12449_/S vssd1 vssd1 vccd1
+ vccd1 _12566_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__07168_ clkbuf_0__07168_/X vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_156_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11517_ _18037_/Q _11329_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _11518_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15285_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15285_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18073_ _18870_/CLK _18073_/D vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12497_ _12493_/X _12494_/X _12495_/X _12496_/X _12768_/S _12407_/A vssd1 vssd1 vccd1
+ vccd1 _12497_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14236_ _18482_/Q _18481_/Q vssd1 vssd1 vccd1 vccd1 _16097_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11448_ _18094_/Q _11273_/X _11448_/S vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11379_ _11341_/X _18124_/Q _11381_/S vssd1 vssd1 vccd1 vccd1 _11380_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03593_ clkbuf_0__03593_/X vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_124_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _18015_/Q _14091_/X _14097_/Y vssd1 vssd1 vccd1 vccd1 _18015_/D sky130_fd_sc_hd__o21a_1
X_18975_ _18987_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15102__821 _15103__822/A vssd1 vssd1 vccd1 vccd1 _18497_/CLK sky130_fd_sc_hd__inv_2
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13066_/A vssd1 vssd1 vccd1 vccd1 _13049_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17926_ _19132_/CLK _17926_/D vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17857_ _17953_/CLK _17857_/D vssd1 vssd1 vccd1 vccd1 _17857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_3_1_wb_clk_i clkbuf_opt_3_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _16802_/X _16805_/X _16982_/A vssd1 vssd1 vccd1 vccd1 _16808_/X sky130_fd_sc_hd__mux2_1
X_17788_ _19128_/CLK _17788_/D vssd1 vssd1 vccd1 vccd1 _17788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16739_ input55/X input71/X _16787_/S vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14146__430 _14150__434/A vssd1 vssd1 vccd1 vccd1 _18038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_179_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09211_ _19153_/Q _09096_/X _09215_/S vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18409_ _18409_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ input5/X vssd1 vssd1 vccd1 vccd1 _19389_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_37_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _18662_/Q vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__buf_2
XFILLER_147_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09073_ _19198_/Q _08880_/X _09077_/S vssd1 vssd1 vccd1 vccd1 _09074_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09975_ _10437_/B _10138_/C _09975_/C vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__nand3b_4
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ _08925_/X _19296_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__mux2_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _09253_/A _08857_/B _13874_/B vssd1 vssd1 vccd1 vccd1 _08857_/X sky130_fd_sc_hd__and3_2
XFILLER_218_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _08788_/A vssd1 vssd1 vccd1 vccd1 _19347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16557__265 _16558__266/A vssd1 vssd1 vccd1 vccd1 _19011_/CLK sky130_fd_sc_hd__inv_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _18387_/Q _10713_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10751_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _09409_/A vssd1 vssd1 vccd1 vccd1 _19061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ _10681_/A vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ _18011_/Q vssd1 vssd1 vccd1 vccd1 _12429_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_200_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12351_ _18007_/Q _18006_/Q vssd1 vssd1 vccd1 vccd1 _12351_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_67_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18007_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04165_ clkbuf_0__04165_/X vssd1 vssd1 vccd1 vccd1 _16085__199/A sky130_fd_sc_hd__clkbuf_16
X_11302_ _11302_/A vssd1 vssd1 vccd1 vccd1 _18155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15070_ _16058_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _18477_/D sky130_fd_sc_hd__nor2_1
X_12282_ _12280_/X _12282_/B vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__and2b_1
XFILLER_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14021_ _13669_/X _14017_/X _14020_/X vssd1 vssd1 vccd1 vccd1 _14021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _11156_/X _18182_/Q _11233_/S vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11164_ _11164_/A vssd1 vssd1 vccd1 vccd1 _18212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10115_ _10112_/X _18718_/Q _10127_/S vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18760_ _18760_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11095_ _11095_/A vssd1 vssd1 vccd1 vccd1 _18240_/D sky130_fd_sc_hd__clkbuf_1
X_15972_ _18864_/Q _15973_/B vssd1 vssd1 vccd1 vccd1 _15974_/B sky130_fd_sc_hd__nor2_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17711_ _17711_/CLK _17711_/D vssd1 vssd1 vccd1 vccd1 _17711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ _14936_/B _14936_/C _14936_/A vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__a21o_1
X_10046_ _18743_/Q _09967_/X _10046_/S vssd1 vssd1 vccd1 vccd1 _10047_/A sky130_fd_sc_hd__mux2_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _18691_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17642_ _19246_/CLK _17642_/D vssd1 vssd1 vccd1 vccd1 _17642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13805_ _13880_/A vssd1 vssd1 vccd1 vccd1 _13805_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17573_ _17573_/CLK _17573_/D vssd1 vssd1 vccd1 vccd1 _17573_/Q sky130_fd_sc_hd__dfxtp_1
X_11997_ _19257_/Q _19258_/Q _19259_/Q _19260_/Q _11995_/X _12067_/S vssd1 vssd1 vccd1
+ vccd1 _11997_/X sky130_fd_sc_hd__mux4_2
XFILLER_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19312_ _19312_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ input67/X _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16525_/A sky130_fd_sc_hd__and3_1
XFILLER_189_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13736_ _17889_/Q _13719_/B _13735_/Y _13726_/X vssd1 vssd1 vccd1 vccd1 _17889_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10948_ _10948_/A vssd1 vssd1 vccd1 vccd1 _18299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19243_ _19247_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16455_ _18973_/Q _16468_/B vssd1 vssd1 vccd1 vccd1 _16455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ _13231_/X _13666_/X _13661_/X vssd1 vssd1 vccd1 vccd1 _13667_/Y sky130_fd_sc_hd__a21oi_1
X_10879_ _18334_/Q _10803_/X _10879_/S vssd1 vssd1 vccd1 vccd1 _10880_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ _12394_/X _12610_/X _12617_/X vssd1 vssd1 vccd1 vccd1 _12619_/B sky130_fd_sc_hd__o21ai_1
X_19174_ _19174_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _14078_/A _13598_/B vssd1 vssd1 vccd1 vccd1 _17844_/D sky130_fd_sc_hd__nor2_1
X_16386_ _18978_/Q _16386_/B vssd1 vssd1 vccd1 vccd1 _16421_/C sky130_fd_sc_hd__xnor2_1
XFILLER_191_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18125_ _18125_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_1
X_12549_ _12476_/Y _12480_/Y _12548_/Y _12478_/Y _12586_/S _12504_/A vssd1 vssd1 vccd1
+ vccd1 _12775_/D sky130_fd_sc_hd__mux4_1
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15337_ _18940_/Q _18903_/Q _18895_/Q _18849_/Q _15248_/X _15252_/X vssd1 vssd1 vccd1
+ vccd1 _15337_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18056_ _18056_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
X_15268_ _15244_/X _15254_/X _15266_/X _15267_/X vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _18080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15199_ _15199_/A vssd1 vssd1 vccd1 vccd1 _15199_/X sky130_fd_sc_hd__buf_1
XFILLER_125_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14330__519 _14330__519/A vssd1 vssd1 vccd1 vccd1 _18154_/CLK sky130_fd_sc_hd__inv_2
X_09760_ _09760_/A vssd1 vssd1 vccd1 vccd1 _18847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18958_ _18958_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17909_ _18007_/CLK _17909_/D vssd1 vssd1 vccd1 vccd1 _17909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09691_ _09691_/A vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__buf_2
XFILLER_132_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14861__782 _14862__783/A vssd1 vssd1 vccd1 vccd1 _18427_/CLK sky130_fd_sc_hd__inv_2
X_18889_ _18889_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825__130 _15826__131/A vssd1 vssd1 vccd1 vccd1 _18805_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09125_ _19187_/Q _09119_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14491__648 _14492__649/A vssd1 vssd1 vccd1 vccd1 _18283_/CLK sky130_fd_sc_hd__inv_2
XFILLER_159_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _09055_/X _19204_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__mux2_1
X_15109__827 _15109__827/A vssd1 vssd1 vccd1 vccd1 _18503_/CLK sky130_fd_sc_hd__inv_2
XFILLER_191_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09958_ _18475_/Q vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_237_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04852_ clkbuf_0__04852_/X vssd1 vssd1 vccd1 vccd1 _17086__69/A sky130_fd_sc_hd__clkbuf_16
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08909_ _18887_/Q vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03803_ clkbuf_0__03803_/X vssd1 vssd1 vccd1 vccd1 _15440__934/A sky130_fd_sc_hd__clkbuf_16
XFILLER_246_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _11383_/B _09892_/B _09888_/X _09870_/X vssd1 vssd1 vccd1 vccd1 _18804_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_218_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14385__564 _14385__564/A vssd1 vssd1 vccd1 vccd1 _18199_/CLK sky130_fd_sc_hd__inv_2
X_11920_ _19230_/Q _17159_/A _12025_/S vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__mux2_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11851_ _13279_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11852_/A sky130_fd_sc_hd__and2_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10802_/A vssd1 vssd1 vccd1 vccd1 _18367_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _19075_/Q _18339_/Q _17573_/Q _18791_/Q _14568_/X _14569_/X vssd1 vssd1 vccd1
+ vccd1 _14571_/B sky130_fd_sc_hd__mux4_2
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11782_ _18066_/Q _13873_/A _08747_/B _11786_/A vssd1 vssd1 vccd1 vccd1 _13352_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03596_ clkbuf_0__03596_/X vssd1 vssd1 vccd1 vccd1 _15142__854/A sky130_fd_sc_hd__clkbuf_16
XFILLER_213_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13521_ _16052_/A _14113_/A _14076_/B vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__and3_1
X_10733_ _10733_/A vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _13150_/X _13437_/X _13450_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _17798_/D
+ sky130_fd_sc_hd__a211oi_1
X_16240_ _16278_/A _16240_/B vssd1 vssd1 vccd1 vccd1 _16240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10664_ _18424_/Q _09732_/X _10670_/S vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12403_ _12622_/A _12626_/A _12631_/A _12638_/B _12366_/X _12368_/X vssd1 vssd1 vccd1
+ vccd1 _12403_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _19146_/Q _13420_/B vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__nand2_4
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16171_ _16171_/A _16171_/B vssd1 vssd1 vccd1 vccd1 _16171_/Y sky130_fd_sc_hd__nor2_1
X_10595_ _10595_/A vssd1 vssd1 vccd1 vccd1 _18487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14392__568 _14393__569/A vssd1 vssd1 vccd1 vccd1 _18203_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15053_ _18468_/Q _15080_/C _15049_/B _18469_/Q vssd1 vssd1 vccd1 vccd1 _15053_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12265_ _12263_/X _12265_/B vssd1 vssd1 vccd1 vccd1 _12266_/A sky130_fd_sc_hd__and2b_1
XFILLER_181_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _14095_/A vssd1 vssd1 vccd1 vccd1 _14060_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16349__241 _16349__241/A vssd1 vssd1 vccd1 vccd1 _18957_/CLK sky130_fd_sc_hd__inv_2
X_11216_ _18189_/Q _11059_/X _11220_/S vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12196_ _17525_/Q _17491_/B vssd1 vssd1 vccd1 vccd1 _12198_/C sky130_fd_sc_hd__xor2_1
Xoutput82 _18924_/Q vssd1 vssd1 vccd1 vccd1 internal_uart_tx sky130_fd_sc_hd__buf_2
X_18812_ _18812_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput93 _11739_/X vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__buf_2
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11147_ _11326_/A vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18743_ _18743_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15955_ _15955_/A _16063_/B vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__or2_1
X_11078_ _11078_/A vssd1 vssd1 vccd1 vccd1 _18247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ _18468_/Q _14906_/B vssd1 vssd1 vccd1 vccd1 _14963_/B sky130_fd_sc_hd__xnor2_1
X_10029_ _10029_/A vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__clkbuf_1
X_18674_ _18674_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15886_ _15886_/A vssd1 vssd1 vccd1 vccd1 _18852_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14286__484 _14286__484/A vssd1 vssd1 vccd1 vccd1 _18119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17625_ _17629_/CLK _17625_/D vssd1 vssd1 vccd1 vccd1 _17625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04013_ _15868_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04013_/X sky130_fd_sc_hd__clkbuf_16
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ _17776_/CLK _17556_/D vssd1 vssd1 vccd1 vccd1 _17556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16507_ _16507_/A _16505_/X vssd1 vssd1 vccd1 vccd1 _16507_/X sky130_fd_sc_hd__or2b_1
X_13719_ _13719_/A _13719_/B vssd1 vssd1 vccd1 vccd1 _13719_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17487_ _19333_/Q _17487_/B vssd1 vssd1 vccd1 vccd1 _17494_/B sky130_fd_sc_hd__xnor2_1
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14699_ _18590_/Q _18304_/Q _17570_/Q _18841_/Q _14615_/X _14641_/X vssd1 vssd1 vccd1
+ vccd1 _14699_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19226_ _19252_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16438_ _18969_/Q _16437_/C _18970_/Q vssd1 vssd1 vccd1 vccd1 _16439_/C sky130_fd_sc_hd__a21oi_1
XFILLER_165_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19157_ _19157_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_1
X_16369_ _17801_/Q _16397_/B vssd1 vssd1 vccd1 vccd1 _16393_/B sky130_fd_sc_hd__or2_1
XFILLER_145_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18108_ _18108_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04846_ _17050_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04846_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_172_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ _19088_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15894__183 _15895__184/A vssd1 vssd1 vccd1 vccd1 _18859_/CLK sky130_fd_sc_hd__inv_2
XFILLER_145_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ _18039_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09812_ _09679_/X _18826_/Q _09818_/S vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _09743_/A vssd1 vssd1 vccd1 vccd1 _18853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09674_ _09674_/A vssd1 vssd1 vccd1 vccd1 _09674_/X sky130_fd_sc_hd__buf_2
XFILLER_227_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _10707_/A vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__buf_2
XFILLER_182_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10380_ _08792_/X _18581_/Q _10382_/S vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__mux2_1
X_09039_ _11332_/A vssd1 vssd1 vccd1 vccd1 _09039_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14868__788 _14869__789/A vssd1 vssd1 vccd1 vccd1 _18433_/CLK sky130_fd_sc_hd__inv_2
X_12050_ _17098_/A vssd1 vssd1 vccd1 vccd1 _17492_/B sky130_fd_sc_hd__buf_4
XFILLER_2_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _11001_/A vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _12911_/X _12952_/B vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__and2b_1
XFILLER_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11903_ _11900_/X _11901_/X _12036_/S vssd1 vssd1 vccd1 vccd1 _11903_/X sky130_fd_sc_hd__mux2_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12877_/X _12883_/B vssd1 vssd1 vccd1 vccd1 _12884_/A sky130_fd_sc_hd__and2b_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16717__334 _16717__334/A vssd1 vssd1 vccd1 vccd1 _19113_/CLK sky130_fd_sc_hd__inv_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _18324_/Q _14543_/X _14589_/X _14621_/X vssd1 vssd1 vccd1 vccd1 _18324_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _17906_/Q vssd1 vssd1 vccd1 vccd1 _11834_/Y sky130_fd_sc_hd__inv_2
X_18390_ _18390_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17758_/Q _19285_/Q _17350_/S vssd1 vssd1 vccd1 vccd1 _17342_/B sky130_fd_sc_hd__mux2_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11765_/A vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_82_wb_clk_i clkbuf_leaf_82_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18670_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13504_ _17812_/Q _13499_/X _13503_/Y vssd1 vssd1 vccd1 vccd1 _17812_/D sky130_fd_sc_hd__o21a_1
X_10716_ _11529_/A _10752_/A vssd1 vssd1 vccd1 vccd1 _10732_/S sky130_fd_sc_hd__nor2_2
XFILLER_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17272_ _17276_/B _17277_/B _17272_/C vssd1 vssd1 vccd1 vccd1 _17273_/A sky130_fd_sc_hd__and3b_1
XFILLER_147_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11696_ _12918_/A vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18971_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19011_ _19011_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
X_16223_ _16223_/A _16223_/B vssd1 vssd1 vccd1 vccd1 _16223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_201_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13435_ _13769_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13447_/S sky130_fd_sc_hd__nor2_1
X_10647_ _10647_/A vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13366_ _11945_/X _13529_/A _13366_/S vssd1 vssd1 vccd1 vccd1 _13367_/B sky130_fd_sc_hd__mux2_1
X_16154_ _16148_/X _16151_/X _16248_/S vssd1 vssd1 vccd1 vccd1 _16154_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10578_ _10132_/X _18493_/Q _10580_/S vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12317_ _12301_/X _12316_/X _17564_/Q vssd1 vssd1 vccd1 vccd1 _12318_/C sky130_fd_sc_hd__a21oi_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13297_ _17758_/Q _13282_/X _13296_/Y vssd1 vssd1 vccd1 vccd1 _17758_/D sky130_fd_sc_hd__o21a_1
XFILLER_114_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12248_ _12248_/A vssd1 vssd1 vccd1 vccd1 _17549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _18466_/Q _15043_/C vssd1 vssd1 vccd1 vccd1 _15038_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03413_ clkbuf_0__03413_/X vssd1 vssd1 vccd1 vccd1 _14835__761/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12179_ _17531_/Q vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16987_ _18218_/Q _18202_/Q _18491_/Q _18194_/Q _09852_/A _09858_/A vssd1 vssd1 vccd1
+ vccd1 _16987_/X sky130_fd_sc_hd__mux4_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18726_ _18726_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15938_ _15938_/A _15938_/B vssd1 vssd1 vccd1 vccd1 _15940_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14442__609 _14442__609/A vssd1 vssd1 vccd1 vccd1 _18244_/CLK sky130_fd_sc_hd__inv_2
X_18657_ _18657_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17608_ _17611_/CLK _17608_/D vssd1 vssd1 vccd1 vccd1 _17608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _19069_/Q _08961_/X _09394_/S vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18588_ _18588_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17539_/CLK _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19209_ _19209_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301__495 _14302__496/A vssd1 vssd1 vccd1 vccd1 _18130_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15672__973 _15673__974/A vssd1 vssd1 vccd1 vccd1 _18690_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17294__71 _17296__73/A vssd1 vssd1 vccd1 vccd1 _19267_/CLK sky130_fd_sc_hd__inv_2
X_09726_ _10698_/A vssd1 vssd1 vccd1 vccd1 _09726_/X sky130_fd_sc_hd__buf_4
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09657_ _09672_/S vssd1 vssd1 vccd1 vccd1 _09666_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_167_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09588_/A vssd1 vssd1 vccd1 vccd1 _18940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14874__792 _14876__794/A vssd1 vssd1 vccd1 vccd1 _18437_/CLK sky130_fd_sc_hd__inv_2
XFILLER_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11550_ _11550_/A vssd1 vssd1 vccd1 vccd1 _17711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10501_ _10501_/A vssd1 vssd1 vccd1 vccd1 _18528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _09130_/X _18053_/Q _11485_/S vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13220_ input61/X _13650_/A vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10432_ _10432_/A _10436_/A vssd1 vssd1 vccd1 vccd1 _10433_/B sky130_fd_sc_hd__or2_1
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13151_ _14136_/B vssd1 vssd1 vccd1 vccd1 _14134_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15838__140 _15840__142/A vssd1 vssd1 vccd1 vccd1 _18815_/CLK sky130_fd_sc_hd__inv_2
XFILLER_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10363_ _10363_/A vssd1 vssd1 vccd1 vccd1 _18589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _12102_/A vssd1 vssd1 vccd1 vccd1 _12102_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ _17698_/Q _12835_/A _12834_/A _17688_/Q _13081_/X vssd1 vssd1 vccd1 vccd1
+ _13082_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10294_ _18616_/Q _10175_/X _10302_/S vssd1 vssd1 vccd1 vccd1 _10295_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12033_ _12031_/X _12032_/X _12037_/S vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16910_ _18214_/Q _18198_/Q _18487_/Q _18190_/Q _16834_/X _09875_/X vssd1 vssd1 vccd1
+ vccd1 _16910_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _19109_/CLK _17890_/D vssd1 vssd1 vccd1 vccd1 _17890_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_238_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16841_ _19137_/Q _16797_/X _16840_/X _15628_/X vssd1 vssd1 vccd1 vccd1 _19137_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16772_ _19133_/Q _19131_/Q _16787_/S vssd1 vssd1 vccd1 vccd1 _16773_/B sky130_fd_sc_hd__mux2_1
XFILLER_219_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13984_ _17974_/Q _13968_/X _13983_/Y vssd1 vssd1 vccd1 vccd1 _17974_/D sky130_fd_sc_hd__o21a_1
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03160_ _14337_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03160_/X sky130_fd_sc_hd__clkbuf_16
X_18511_ _18511_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _15754_/A vssd1 vssd1 vccd1 vccd1 _15723_/X sky130_fd_sc_hd__buf_1
XFILLER_206_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12935_ _17659_/Q _12924_/X _12920_/X _17661_/Q vssd1 vssd1 vccd1 vccd1 _12942_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03091_ _14151_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03091_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18442_ _18442_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12830_/X _12866_/B vssd1 vssd1 vccd1 vccd1 _12867_/A sky130_fd_sc_hd__and2b_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052__41 _17053__42/A vssd1 vssd1 vccd1 vccd1 _19190_/CLK sky130_fd_sc_hd__inv_2
XFILLER_222_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14597_/X _14603_/X _14673_/S vssd1 vssd1 vccd1 vccd1 _14605_/X sky130_fd_sc_hd__mux2_2
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11817_ _17911_/Q _11812_/X _11809_/Y input14/X _11796_/X vssd1 vssd1 vccd1 vccd1
+ _11817_/X sky130_fd_sc_hd__a221o_1
X_18373_ _18373_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _18651_/Q _15585_/B _15585_/C vssd1 vssd1 vccd1 vccd1 _15595_/C sky130_fd_sc_hd__and3_1
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12795_/X _12797_/B vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__and2b_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17763_/Q _19280_/Q _17333_/S vssd1 vssd1 vccd1 vccd1 _17325_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14536_ _14536_/A vssd1 vssd1 vccd1 vccd1 _14536_/X sky130_fd_sc_hd__buf_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11748_ _17771_/Q _17880_/Q vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__and2b_4
Xclkbuf_1_1__f__03962_ clkbuf_0__03962_/X vssd1 vssd1 vccd1 vccd1 _15651__956/A sky130_fd_sc_hd__clkbuf_16
XFILLER_239_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140__425 _14141__426/A vssd1 vssd1 vccd1 vccd1 _18033_/CLK sky130_fd_sc_hd__inv_2
XFILLER_230_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _19257_/Q vssd1 vssd1 vccd1 vccd1 _17262_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_187_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03993_ _15805_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03993_/X sky130_fd_sc_hd__clkbuf_16
X_11679_ _16584_/A vssd1 vssd1 vccd1 vccd1 _16578_/A sky130_fd_sc_hd__buf_6
X_16206_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16206_/X sky130_fd_sc_hd__clkbuf_2
X_13418_ _13274_/X _13395_/X _13408_/X vssd1 vssd1 vccd1 vccd1 _13418_/Y sky130_fd_sc_hd__a21oi_1
X_17186_ _19239_/Q _17186_/B _17186_/C _17186_/D vssd1 vssd1 vccd1 vccd1 _17203_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_128_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16137_ _16280_/A _16137_/B vssd1 vssd1 vccd1 vccd1 _16137_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ _19145_/Q vssd1 vssd1 vccd1 vccd1 _14243_/A sky130_fd_sc_hd__buf_2
XFILLER_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15747__1034 _15747__1034/A vssd1 vssd1 vccd1 vccd1 _18751_/CLK sky130_fd_sc_hd__inv_2
X_16068_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16068_/X sky130_fd_sc_hd__buf_1
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15019_ _18463_/Q _15020_/B vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__nor2_1
XFILLER_130_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08890_ _11637_/A vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__buf_4
XFILLER_190_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04376_ clkbuf_0__04376_/X vssd1 vssd1 vccd1 vccd1 _16352__244/A sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09511_ _09511_/A vssd1 vssd1 vccd1 vccd1 _19004_/D sky130_fd_sc_hd__clkbuf_1
X_18709_ _18709_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09442_ _09442_/A _09442_/B _08842_/Y vssd1 vssd1 vccd1 vccd1 _16559_/C sky130_fd_sc_hd__or3b_2
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03189_ clkbuf_0__03189_/X vssd1 vssd1 vccd1 vccd1 _14486__644/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09373_ _19076_/Q _09112_/X _09375_/S vssd1 vssd1 vccd1 vccd1 _09374_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15151__861 _15153__863/A vssd1 vssd1 vccd1 vccd1 _18537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16631__273 _16631__273/A vssd1 vssd1 vccd1 vccd1 _19047_/CLK sky130_fd_sc_hd__inv_2
X_14299__494 _14299__494/A vssd1 vssd1 vccd1 vccd1 _18129_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_1 _18064_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761__701 _14763__703/A vssd1 vssd1 vccd1 vccd1 _18344_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03982_ clkbuf_0__03982_/X vssd1 vssd1 vccd1 vccd1 _15779_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16673__307 _16674__308/A vssd1 vssd1 vccd1 vccd1 _19081_/CLK sky130_fd_sc_hd__inv_2
X_09709_ _09709_/A vssd1 vssd1 vccd1 vccd1 _18894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10981_ _18284_/Q _09764_/X hold11/X vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12720_ _12727_/D _12720_/B vssd1 vssd1 vccd1 vccd1 _17623_/D sky130_fd_sc_hd__nor2_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12651_ _17604_/Q _17603_/Q _17602_/Q _12651_/D vssd1 vssd1 vccd1 vccd1 _12666_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_215_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11602_ _11617_/S vssd1 vssd1 vccd1 vccd1 _11611_/S sky130_fd_sc_hd__clkbuf_2
X_12582_ _12840_/A vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__inv_2
X_15370_ _19004_/Q _18966_/Q _18958_/Q _17547_/Q _15209_/X _15212_/X vssd1 vssd1 vccd1
+ vccd1 _15370_/X sky130_fd_sc_hd__mux4_2
XFILLER_180_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03416_ clkbuf_0__03416_/X vssd1 vssd1 vccd1 vccd1 _14851__774/A sky130_fd_sc_hd__clkbuf_16
XFILLER_196_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11533_ _08868_/X _17718_/Q _11539_/S vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11464_ _11464_/A vssd1 vssd1 vccd1 vccd1 _18061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _17734_/Q _13208_/B vssd1 vssd1 vccd1 vccd1 _13203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10415_ _10406_/B _10417_/A _10414_/Y vssd1 vssd1 vccd1 vccd1 _18566_/D sky130_fd_sc_hd__o21a_1
X_15679__979 _15679__979/A vssd1 vssd1 vccd1 vccd1 _18696_/CLK sky130_fd_sc_hd__inv_2
XFILLER_152_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11395_ _11395_/A vssd1 vssd1 vccd1 vccd1 _18118_/D sky130_fd_sc_hd__clkbuf_1
X_14183_ input78/X input54/X _11865_/B vssd1 vssd1 vccd1 vccd1 _14249_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ _14053_/A _13169_/B vssd1 vssd1 vccd1 vccd1 _14136_/B sky130_fd_sc_hd__and2_1
XFILLER_124_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _18595_/Q _10345_/X _10352_/S vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18991_ _18996_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A vssd1 vssd1 vccd1 vccd1 _17698_/D sky130_fd_sc_hd__clkbuf_1
X_17942_ _17951_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10277_ _10277_/A vssd1 vssd1 vccd1 vccd1 _18624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12016_ _12103_/A _12104_/A _12016_/S vssd1 vssd1 vccd1 vccd1 _12016_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17873_ _17878_/CLK _17873_/D vssd1 vssd1 vccd1 vccd1 _17873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16824_ _18243_/Q _18235_/Q _18227_/Q _18219_/Q _16822_/X _16823_/X vssd1 vssd1 vccd1
+ vccd1 _16825_/B sky130_fd_sc_hd__mux4_1
XFILLER_226_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16755_ _19129_/Q _16771_/B _16754_/X vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13967_ _13973_/A vssd1 vssd1 vccd1 vccd1 _13967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ _12918_/A vssd1 vssd1 vccd1 vccd1 _16690_/A sky130_fd_sc_hd__clkbuf_4
X_16686_ _19091_/Q vssd1 vssd1 vccd1 vccd1 _16687_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _17942_/Q _13879_/X _13897_/Y vssd1 vssd1 vccd1 vccd1 _17942_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18425_ _18425_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15637_ _16057_/A _15638_/B vssd1 vssd1 vccd1 vccd1 _18664_/D sky130_fd_sc_hd__nor2_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12849_ _12849_/A _12849_/B _12849_/C _12849_/D vssd1 vssd1 vccd1 vccd1 _12860_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_62_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18356_ _18356_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
X_15568_ _15579_/A _15568_/B _15571_/B vssd1 vssd1 vccd1 vccd1 _15568_/X sky130_fd_sc_hd__or3_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17307_ _17768_/Q _19275_/Q _17381_/B vssd1 vssd1 vccd1 vccd1 _17308_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18287_ _18287_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_1
X_15499_ _18650_/Q _15499_/B vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__or2_1
X_17238_ _17250_/D vssd1 vssd1 vccd1 vccd1 _17246_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__03976_ _15723_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03976_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_162_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17169_ _17173_/B _17169_/B _17169_/C vssd1 vssd1 vccd1 vccd1 _17169_/X sky130_fd_sc_hd__and3_1
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09991_ _09991_/A vssd1 vssd1 vccd1 vccd1 _18768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _08941_/X _19292_/Q _08942_/S vssd1 vssd1 vccd1 vccd1 _08943_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14413__585 _14414__586/A vssd1 vssd1 vccd1 vccd1 _18220_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__04528_ _16549_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04528_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_215_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14825__753 _14826__754/A vssd1 vssd1 vccd1 vccd1 _18396_/CLK sky130_fd_sc_hd__inv_2
X_08873_ _08873_/A vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _09425_/A vssd1 vssd1 vccd1 vccd1 _19054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09356_ _19083_/Q _09280_/X _09356_/S vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__mux2_1
X_16336__232 _16338__234/A vssd1 vssd1 vccd1 vccd1 _18948_/CLK sky130_fd_sc_hd__inv_2
XFILLER_200_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09287_ _19118_/Q _08949_/X _09293_/S vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14455__619 _14455__619/A vssd1 vssd1 vccd1 vccd1 _18254_/CLK sky130_fd_sc_hd__inv_2
XFILLER_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10200_ _10200_/A vssd1 vssd1 vccd1 vccd1 _18687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11180_ _11159_/X _18205_/Q _11184_/S vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10131_ _10131_/A vssd1 vssd1 vccd1 vccd1 _18713_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10062_ _10062_/A vssd1 vssd1 vccd1 vccd1 _18739_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16343__236 _16344__237/A vssd1 vssd1 vccd1 vccd1 _18952_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03965_ clkbuf_0__03965_/X vssd1 vssd1 vccd1 vccd1 _15667__969/A sky130_fd_sc_hd__clkbuf_16
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15197__883 _15198__884/A vssd1 vssd1 vccd1 vccd1 _18562_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14870_ _14870_/A vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__buf_1
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13821_ _19147_/Q input64/X _13828_/B vssd1 vssd1 vccd1 vccd1 _13821_/X sky130_fd_sc_hd__and3_1
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12234__379 _12234__379/A vssd1 vssd1 vccd1 vccd1 _17543_/CLK sky130_fd_sc_hd__inv_2
XFILLER_141_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13752_ _14083_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13752_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_108 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_119 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10964_ _10964_/A vssd1 vssd1 vccd1 vccd1 _18292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_6_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_16638__279 _16638__279/A vssd1 vssd1 vccd1 vccd1 _19053_/CLK sky130_fd_sc_hd__inv_2
X_12703_ _12703_/A _12703_/B vssd1 vssd1 vccd1 vccd1 _17618_/D sky130_fd_sc_hd__nor2_1
XFILLER_243_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16471_ _16471_/A vssd1 vssd1 vccd1 vccd1 _16498_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13683_ _13688_/A vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15746__1033 _15746__1033/A vssd1 vssd1 vccd1 vccd1 _18750_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18210_ _18210_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
X_14280__479 _14280__479/A vssd1 vssd1 vccd1 vccd1 _18114_/CLK sky130_fd_sc_hd__inv_2
X_12634_ _12638_/B _12641_/D vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__and2_1
X_19190_ _19190_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388__891 _15389__892/A vssd1 vssd1 vccd1 vccd1 _18578_/CLK sky130_fd_sc_hd__inv_2
XFILLER_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18141_ _18141_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
X_15353_ _19003_/Q _18965_/Q _18957_/Q _17546_/Q _15273_/X _15212_/X vssd1 vssd1 vccd1
+ vccd1 _15353_/X sky130_fd_sc_hd__mux4_2
X_12565_ _17590_/Q _17591_/Q _12610_/B _12610_/A _12555_/X _12556_/X vssd1 vssd1 vccd1
+ vccd1 _12565_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__07167_ clkbuf_0__07167_/X vssd1 vssd1 vccd1 vccd1 _17390_/A sky130_fd_sc_hd__clkbuf_16
X_11516_ _11516_/A vssd1 vssd1 vccd1 vccd1 _18038_/D sky130_fd_sc_hd__clkbuf_1
X_18072_ _18072_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
X_15284_ _15284_/A vssd1 vssd1 vccd1 vccd1 _15284_/Y sky130_fd_sc_hd__inv_2
X_12496_ _17595_/Q _12622_/A _12626_/A _12631_/A _12366_/X _12368_/X vssd1 vssd1 vccd1
+ vccd1 _12496_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14235_ _14235_/A vssd1 vssd1 vccd1 vccd1 _18087_/D sky130_fd_sc_hd__clkbuf_1
X_14768__707 _14768__707/A vssd1 vssd1 vccd1 vccd1 _18350_/CLK sky130_fd_sc_hd__inv_2
XFILLER_236_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11447_ _11447_/A vssd1 vssd1 vccd1 vccd1 _18095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14166_ _14166_/A vssd1 vssd1 vccd1 vccd1 _14166_/X sky130_fd_sc_hd__buf_1
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11378_ _11378_/A vssd1 vssd1 vccd1 vccd1 _18125_/D sky130_fd_sc_hd__clkbuf_1
X_12321__385 _12322__386/A vssd1 vssd1 vccd1 vccd1 _17566_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03592_ clkbuf_0__03592_/X vssd1 vssd1 vccd1 vccd1 _15122__838/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10329_ _10620_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10352_/S sky130_fd_sc_hd__nor2_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _13719_/A _14092_/X _14096_/X vssd1 vssd1 vccd1 vccd1 _14097_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _19135_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13048_ _13048_/A vssd1 vssd1 vccd1 vccd1 _17693_/D sky130_fd_sc_hd__clkbuf_1
X_17925_ _19132_/CLK _17925_/D vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17856_ _17953_/CLK _17856_/D vssd1 vssd1 vccd1 vccd1 _17856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _16820_/A vssd1 vssd1 vccd1 vccd1 _16982_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17787_ _17922_/CLK _17787_/D vssd1 vssd1 vccd1 vccd1 _17787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14999_ _14999_/A _15005_/B vssd1 vssd1 vccd1 vccd1 _14999_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16738_ _16741_/S vssd1 vssd1 vccd1 vccd1 _16787_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09210_ _09210_/A vssd1 vssd1 vccd1 vccd1 _19154_/D sky130_fd_sc_hd__clkbuf_1
X_18408_ _18408_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19388_ input3/X vssd1 vssd1 vccd1 vccd1 _19388_/X sky130_fd_sc_hd__buf_8
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09141_ _09141_/A vssd1 vssd1 vccd1 vccd1 _19182_/D sky130_fd_sc_hd__clkbuf_1
X_18339_ _18339_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09072_ _09072_/A vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _10638_/B vssd1 vssd1 vccd1 vccd1 _10528_/B sky130_fd_sc_hd__buf_4
XFILLER_44_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08925_ _09685_/A vssd1 vssd1 vccd1 vccd1 _08925_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08856_ _09250_/A _08997_/C vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__nor2_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08787_ _19347_/Q _08786_/X _08796_/S vssd1 vssd1 vccd1 vccd1 _08788_/A sky130_fd_sc_hd__mux2_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _08933_/X _19061_/Q _09412_/S vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10680_ _18417_/Q _09729_/X _10682_/S vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _10456_/A vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__buf_4
XFILLER_178_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _18005_/Q vssd1 vssd1 vccd1 vccd1 _14067_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__04164_ clkbuf_0__04164_/X vssd1 vssd1 vccd1 vccd1 _16077__192/A sky130_fd_sc_hd__clkbuf_16
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ _18155_/Q _11282_/X _11301_/S vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__mux2_1
X_12281_ _17559_/Q _18018_/Q _12287_/S vssd1 vssd1 vccd1 vccd1 _12282_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14020_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11232_ _11232_/A vssd1 vssd1 vccd1 vccd1 _18183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15164__871 _15165__872/A vssd1 vssd1 vccd1 vccd1 _18547_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11163_ _11162_/X _18212_/Q _11166_/S vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16087__200 _16091__204/A vssd1 vssd1 vccd1 vccd1 _18905_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_36_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _18027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10114_ _10136_/S vssd1 vssd1 vccd1 vccd1 _10127_/S sky130_fd_sc_hd__buf_2
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _09035_/X _18240_/Q _11098_/S vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15971_ _15969_/X _15970_/X _16033_/A vssd1 vssd1 vccd1 vccd1 _18863_/D sky130_fd_sc_hd__a21oi_1
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _17710_/CLK _17710_/D vssd1 vssd1 vccd1 vccd1 _17710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ _18465_/Q _14922_/B vssd1 vssd1 vccd1 vccd1 _14936_/C sky130_fd_sc_hd__nand2_1
X_10045_ _10045_/A vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17086__69 _17086__69/A vssd1 vssd1 vccd1 vccd1 _19218_/CLK sky130_fd_sc_hd__inv_2
X_18690_ _18690_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _19247_/CLK _17641_/D vssd1 vssd1 vccd1 vccd1 _17641_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _17911_/Q _13796_/X _13803_/Y vssd1 vssd1 vccd1 vccd1 _17911_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17572_ _17572_/CLK _17572_/D vssd1 vssd1 vccd1 vccd1 _17572_/Q sky130_fd_sc_hd__dfxtp_1
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14784_/X sky130_fd_sc_hd__buf_1
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _19253_/Q _19254_/Q _17250_/B _17252_/A _11995_/X _11938_/A vssd1 vssd1 vccd1
+ vccd1 _11996_/X sky130_fd_sc_hd__mux4_2
XFILLER_205_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19311_ _19311_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16523_ _16523_/A vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__clkbuf_1
X_13735_ _13792_/A _13735_/B vssd1 vssd1 vccd1 vccd1 _13735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10947_ _18299_/Q _10910_/X hold16/X vssd1 vssd1 vccd1 vccd1 _10948_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19242_ _19247_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16454_ _16467_/A _16454_/B _16458_/B vssd1 vssd1 vccd1 vccd1 _16454_/X sky130_fd_sc_hd__or3_1
X_13666_ _13666_/A vssd1 vssd1 vccd1 vccd1 _13666_/X sky130_fd_sc_hd__clkbuf_2
X_10878_ _10878_/A vssd1 vssd1 vccd1 vccd1 _18335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12617_ _12695_/A vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__clkbuf_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19173_ _19173_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _17798_/Q _16389_/B vssd1 vssd1 vccd1 vccd1 _16386_/B sky130_fd_sc_hd__xor2_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _13596_/Y _13493_/A _13597_/S vssd1 vssd1 vccd1 vccd1 _13598_/B sky130_fd_sc_hd__mux2_1
XFILLER_223_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08199_ clkbuf_0__08199_/X vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__clkbuf_16
X_18124_ _18124_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_1
X_15336_ _19321_/Q _19305_/Q _19297_/Q _19272_/Q _15273_/X _15212_/X vssd1 vssd1 vccd1
+ vccd1 _15336_/X sky130_fd_sc_hd__mux4_2
X_12548_ _12548_/A vssd1 vssd1 vccd1 vccd1 _12548_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18055_ _18055_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
X_15267_ _15267_/A vssd1 vssd1 vccd1 vccd1 _15267_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12479_ _12390_/X _12376_/X _12547_/S vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17006_ _17006_/A vssd1 vssd1 vccd1 vccd1 _17006_/X sky130_fd_sc_hd__buf_1
XFILLER_160_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14218_ _13759_/A input38/X _14218_/S vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15438__932 _15439__933/A vssd1 vssd1 vccd1 vccd1 _18619_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18957_ _18957_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17908_ _17922_/CLK _17908_/D vssd1 vssd1 vccd1 vccd1 _17908_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09690_ _09690_/A vssd1 vssd1 vccd1 vccd1 _18901_/D sky130_fd_sc_hd__clkbuf_1
X_18888_ _18888_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17839_ _17840_/CLK _17839_/D vssd1 vssd1 vccd1 vccd1 _17839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14525__675 _14529__679/A vssd1 vssd1 vccd1 vccd1 _18310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_208_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ _09146_/S vssd1 vssd1 vccd1 vccd1 _09137_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09055_ _11344_/A vssd1 vssd1 vccd1 vccd1 _09055_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15745__1032 _15746__1033/A vssd1 vssd1 vccd1 vccd1 _18749_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832__135 _15833__136/A vssd1 vssd1 vccd1 vccd1 _18810_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _09957_/A vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__04851_ clkbuf_0__04851_/X vssd1 vssd1 vccd1 vccd1 _17080__64/A sky130_fd_sc_hd__clkbuf_16
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ _08908_/A vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09888_ _10987_/B _10985_/B vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__03802_ clkbuf_0__03802_/X vssd1 vssd1 vccd1 vccd1 _15434__929/A sky130_fd_sc_hd__clkbuf_16
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ hold7/A hold20/A hold21/A vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__and3_1
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11850_ _17921_/Q _11839_/X _11840_/X _17902_/Q vssd1 vssd1 vccd1 vccd1 _11851_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16082__196 _16085__199/A vssd1 vssd1 vccd1 vccd1 _18901_/CLK sky130_fd_sc_hd__inv_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10801_ _18367_/Q _10800_/X _10804_/S vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__mux2_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _18067_/Q vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__buf_2
X_14426__595 _14427__596/A vssd1 vssd1 vccd1 vccd1 _18230_/CLK sky130_fd_sc_hd__inv_2
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03595_ clkbuf_0__03595_/X vssd1 vssd1 vccd1 vccd1 _15136__849/A sky130_fd_sc_hd__clkbuf_16
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13520_ _13520_/A _13520_/B vssd1 vssd1 vccd1 vccd1 _16052_/A sky130_fd_sc_hd__nor2_2
XFILLER_242_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10732_ _18395_/Q _10713_/X _10732_/S vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13451_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10663_ _10663_/A vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12402_ _17599_/Q vssd1 vssd1 vccd1 vccd1 _12638_/B sky130_fd_sc_hd__clkbuf_1
X_16170_ _18595_/Q _18611_/Q _18737_/Q _18518_/Q _16106_/X _16138_/X vssd1 vssd1 vccd1
+ vccd1 _16171_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13382_ _17117_/A _13366_/S _13381_/Y vssd1 vssd1 vccd1 vccd1 _17782_/D sky130_fd_sc_hd__o21a_1
XFILLER_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10594_ _09043_/X _18487_/Q _10594_/S vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12333_ _12333_/A vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__buf_1
XFILLER_177_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15052_ _15052_/A vssd1 vssd1 vccd1 vccd1 _18468_/D sky130_fd_sc_hd__clkbuf_1
X_12264_ _17554_/Q _18023_/Q _12270_/S vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__mux2_1
XFILLER_177_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _17981_/Q _13989_/X _14002_/Y vssd1 vssd1 vccd1 vccd1 _17981_/D sky130_fd_sc_hd__o21a_1
X_11215_ _11215_/A vssd1 vssd1 vccd1 vccd1 _18190_/D sky130_fd_sc_hd__clkbuf_1
X_12195_ _12195_/A vssd1 vssd1 vccd1 vccd1 _17491_/B sky130_fd_sc_hd__buf_4
XFILLER_150_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18811_ _18811_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput83 _11774_/A vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__buf_2
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11146_ _11146_/A vssd1 vssd1 vccd1 vccd1 _18218_/D sky130_fd_sc_hd__clkbuf_1
Xoutput94 _11734_/X vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__buf_2
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17059__47 _17061__49/A vssd1 vssd1 vccd1 vccd1 _19196_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11077_ _09039_/X _18247_/Q _11079_/S vssd1 vssd1 vccd1 vccd1 _11078_/A sky130_fd_sc_hd__mux2_1
X_15954_ _15945_/X _15954_/B _15954_/C vssd1 vssd1 vccd1 vccd1 _16063_/B sky130_fd_sc_hd__and3b_1
X_18742_ _18742_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _17845_/Q _14913_/B vssd1 vssd1 vccd1 vccd1 _14906_/B sky130_fd_sc_hd__xor2_1
X_10028_ _18751_/Q _09967_/X _10028_/S vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18673_ _18673_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _16036_/A _18852_/Q _16010_/A vssd1 vssd1 vccd1 vccd1 _15886_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _17629_/CLK _17624_/D vssd1 vssd1 vccd1 vccd1 _17624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04012_ _15862_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04012_/X sky130_fd_sc_hd__clkbuf_16
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17555_ _17776_/CLK _17555_/D vssd1 vssd1 vccd1 vccd1 _17555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11979_ _19230_/Q vssd1 vssd1 vccd1 vccd1 _17158_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16506_ _16506_/A _18986_/Q _16511_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16507_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_232_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13718_ _17882_/Q _13715_/X _13717_/Y _13710_/X vssd1 vssd1 vccd1 vccd1 _17882_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_232_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17486_ _19327_/Q _12182_/A _12180_/A _19324_/Q vssd1 vssd1 vccd1 vccd1 _17494_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14698_ _14736_/A _14698_/B vssd1 vssd1 vccd1 vccd1 _14698_/Y sky130_fd_sc_hd__nor2_1
X_19225_ _19261_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ _18970_/Q _18969_/Q _16437_/C vssd1 vssd1 vccd1 vccd1 _16445_/B sky130_fd_sc_hd__and3_1
XFILLER_177_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13649_ _13649_/A vssd1 vssd1 vccd1 vccd1 _13649_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19156_ _19156_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16368_ _17804_/Q _17803_/Q _17802_/Q _16412_/B vssd1 vssd1 vccd1 vccd1 _16397_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_160_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18107_ _18107_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15319_ _19001_/Q _18963_/Q _18955_/Q _17544_/Q _15273_/X _15212_/X vssd1 vssd1 vccd1
+ vccd1 _15319_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_0__04845_ _17044_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04845_/X sky130_fd_sc_hd__clkbuf_16
X_19087_ _19087_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_1
X_16299_ _18996_/Q vssd1 vssd1 vccd1 vccd1 _16514_/A sky130_fd_sc_hd__inv_2
XFILLER_173_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18038_ _18038_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09811_ _09811_/A vssd1 vssd1 vccd1 vccd1 _18827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _18853_/Q _09741_/X _09742_/S vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03589_ _15100_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03589_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09673_ _09673_/A vssd1 vssd1 vccd1 vccd1 _18906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12334__395 _12335__396/A vssd1 vssd1 vccd1 vccd1 _17576_/CLK sky130_fd_sc_hd__inv_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115__832 _15117__834/A vssd1 vssd1 vccd1 vccd1 _18508_/CLK sky130_fd_sc_hd__inv_2
XFILLER_195_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09107_ _18989_/Q vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__buf_4
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ _18665_/Q vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11000_ _18277_/Q _09139_/X _11004_/S vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _17966_/Q _17671_/Q _13022_/B vssd1 vssd1 vccd1 vccd1 _12952_/B sky130_fd_sc_hd__mux2_1
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11902_ _17780_/Q vssd1 vssd1 vccd1 vccd1 _12036_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12882_ _17978_/Q _17658_/Q _12891_/S vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__mux2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _09433_/X _14605_/X _14620_/Y vssd1 vssd1 vccd1 vccd1 _14621_/X sky130_fd_sc_hd__a21o_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _17926_/Q _11815_/X _11848_/A _11832_/X vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17437_/A vssd1 vssd1 vccd1 vccd1 _17340_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14552_ _19047_/Q vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__buf_2
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _18002_/Q _17884_/Q vssd1 vssd1 vccd1 vccd1 _11765_/A sky130_fd_sc_hd__and2b_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _13285_/X _13500_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _13503_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17274_/C _17270_/C _17274_/B vssd1 vssd1 vccd1 vccd1 _17272_/C sky130_fd_sc_hd__a21o_1
XFILLER_158_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10715_ _10715_/A vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11695_ _12828_/A vssd1 vssd1 vccd1 vccd1 _12918_/A sky130_fd_sc_hd__buf_4
X_19010_ _19010_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16222_ _18441_/Q _18691_/Q _18699_/Q _18707_/Q _16198_/X _16172_/X vssd1 vssd1 vccd1
+ vccd1 _16223_/B sky130_fd_sc_hd__mux4_1
XFILLER_201_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13434_ _13434_/A vssd1 vssd1 vccd1 vccd1 _13434_/X sky130_fd_sc_hd__buf_6
XFILLER_139_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10646_ _09268_/X _18433_/Q _10648_/S vssd1 vssd1 vccd1 vccd1 _10647_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _16289_/S vssd1 vssd1 vccd1 vccd1 _16248_/S sky130_fd_sc_hd__clkbuf_2
X_13365_ _16689_/A _13365_/B _14076_/B vssd1 vssd1 vccd1 vccd1 _13366_/S sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_51_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19247_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10577_ _10577_/A vssd1 vssd1 vccd1 vccd1 _18494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12316_ _12316_/A _12316_/B _12316_/C _12316_/D vssd1 vssd1 vccd1 vccd1 _12316_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04530_ clkbuf_0__04530_/X vssd1 vssd1 vccd1 vccd1 _16626__269/A sky130_fd_sc_hd__clkbuf_16
XFILLER_127_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _13240_/X _13288_/X _13293_/X vssd1 vssd1 vccd1 vccd1 _13296_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15035_ _15035_/A vssd1 vssd1 vccd1 vccd1 _18465_/D sky130_fd_sc_hd__clkbuf_1
X_16724__339 _16724__339/A vssd1 vssd1 vccd1 vccd1 _19118_/CLK sky130_fd_sc_hd__inv_2
X_12247_ _12245_/X _12247_/B vssd1 vssd1 vccd1 vccd1 _12248_/A sky130_fd_sc_hd__and2b_1
XFILLER_64_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03412_ clkbuf_0__03412_/X vssd1 vssd1 vccd1 vccd1 _14829__756/A sky130_fd_sc_hd__clkbuf_16
XFILLER_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12178_ _12178_/A vssd1 vssd1 vccd1 vccd1 _17530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11129_ _11129_/A vssd1 vssd1 vccd1 vccd1 _18225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16986_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18725_ _18725_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _17817_/Q _15937_/B vssd1 vssd1 vccd1 vccd1 _15938_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18656_ _18657_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_1
X_15868_ _15890_/A vssd1 vssd1 vccd1 vccd1 _15868_/X sky130_fd_sc_hd__buf_1
XFILLER_188_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17607_ _17611_/CLK _17607_/D vssd1 vssd1 vccd1 vccd1 _17607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18587_ _18587_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_1
X_15799_ _15799_/A vssd1 vssd1 vccd1 vccd1 _15799_/X sky130_fd_sc_hd__buf_1
XFILLER_225_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17538_ _17538_/CLK _17538_/D vssd1 vssd1 vccd1 vccd1 _17538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15744__1031 _15746__1033/A vssd1 vssd1 vccd1 vccd1 _18748_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17469_ _17454_/X _17469_/B vssd1 vssd1 vccd1 vccd1 _17470_/A sky130_fd_sc_hd__and2b_1
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19208_ _19208_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19139_ _19144_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16330__227 _16332__229/A vssd1 vssd1 vccd1 vccd1 _18943_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ _09725_/A vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09656_ _10157_/A _10546_/B vssd1 vssd1 vccd1 vccd1 _09672_/S sky130_fd_sc_hd__nor2_2
XFILLER_167_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09587_ _18940_/Q _09489_/X _09591_/S vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__mux2_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10500_ _10123_/X _18528_/Q _10502_/S vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11480_ _11480_/A vssd1 vssd1 vccd1 vccd1 _18054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ _10424_/B _10424_/C _10430_/Y vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13150_ _13783_/A vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__buf_6
XFILLER_100_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10362_ _18589_/Q _09729_/X _10364_/S vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12101_ _12096_/X _12100_/X _12109_/S vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _17689_/Q _13081_/B vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__xor2_1
X_10293_ _10308_/S vssd1 vssd1 vccd1 vccd1 _10302_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_105_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _11910_/X _11913_/X _12032_/S vssd1 vssd1 vccd1 vccd1 _12032_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16840_ _09845_/X _16817_/X _16839_/Y vssd1 vssd1 vccd1 vccd1 _16840_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _19132_/Q _16771_/B vssd1 vssd1 vccd1 vccd1 _16771_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13983_ _13733_/A _13973_/X _13978_/X vssd1 vssd1 vccd1 vccd1 _13983_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18510_ _18510_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ _17666_/Q _13090_/B vssd1 vssd1 vccd1 vccd1 _12942_/A sky130_fd_sc_hd__xnor2_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03090_ _14145_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03090_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18441_ _18441_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _17983_/Q _17653_/Q _12944_/B vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__mux2_1
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14604_ _14604_/A vssd1 vssd1 vccd1 vccd1 _14673_/S sky130_fd_sc_hd__buf_2
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _16689_/A vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__buf_2
X_18372_ _18372_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15584_ _18651_/Q _15584_/B vssd1 vssd1 vccd1 vccd1 _15586_/B sky130_fd_sc_hd__nor2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _17641_/Q _17994_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12797_/B sky130_fd_sc_hd__mux2_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17323_ _17437_/A vssd1 vssd1 vccd1 vccd1 _17323_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11747_/A vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_230_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17254_ _17254_/A vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03992_ _15799_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03992_/X sky130_fd_sc_hd__clkbuf_16
X_11678_ _13428_/A vssd1 vssd1 vccd1 vccd1 _16584_/A sky130_fd_sc_hd__buf_4
X_16205_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16205_/X sky130_fd_sc_hd__clkbuf_4
X_13417_ _17790_/Q _13393_/X _13416_/Y vssd1 vssd1 vccd1 vccd1 _17790_/D sky130_fd_sc_hd__o21a_1
X_17185_ _17186_/B _17184_/B _17184_/Y _17164_/X vssd1 vssd1 vccd1 vccd1 _19238_/D
+ sky130_fd_sc_hd__o211a_1
X_10629_ _10629_/A vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _18525_/Q _18533_/Q _18541_/Q _18549_/Q _10404_/A _16102_/X vssd1 vssd1 vccd1
+ vccd1 _16137_/B sky130_fd_sc_hd__mux4_1
X_13348_ _17775_/Q vssd1 vssd1 vccd1 vccd1 _17101_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ _16308_/A vssd1 vssd1 vccd1 vccd1 _16067_/X sky130_fd_sc_hd__buf_1
X_13279_ _13279_/A _13365_/B _14031_/B vssd1 vssd1 vccd1 vccd1 _13288_/A sky130_fd_sc_hd__and3_2
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15018_ _15059_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__04375_ clkbuf_0__04375_/X vssd1 vssd1 vccd1 vccd1 _16344__237/A sky130_fd_sc_hd__clkbuf_16
XFILLER_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16969_ _09859_/A _16968_/X _16886_/X vssd1 vssd1 vccd1 vccd1 _16969_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _19004_/Q _09481_/X _09518_/S vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18708_ _18708_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09441_/A _09441_/B _09441_/C _09441_/D vssd1 vssd1 vccd1 vccd1 _09442_/B
+ sky130_fd_sc_hd__or4_1
X_18639_ _18639_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03188_ clkbuf_0__03188_/X vssd1 vssd1 vccd1 vccd1 _14487_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_18_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ _09372_/A vssd1 vssd1 vccd1 vccd1 _19077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03981_ clkbuf_0__03981_/X vssd1 vssd1 vccd1 vccd1 _15753__1039/A sky130_fd_sc_hd__clkbuf_16
XINSDIODE2_2 _18924_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _09685_/X _18894_/Q _09710_/S vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10980_/A vssd1 vssd1 vccd1 vccd1 _18285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09639_ _09639_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09640_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _12650_/A vssd1 vssd1 vccd1 vccd1 _17603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ _11601_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11617_/S sky130_fd_sc_hd__nor2_2
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12581_ _12469_/S _12578_/X _12580_/X vssd1 vssd1 vccd1 vccd1 _12840_/A sky130_fd_sc_hd__o21ai_2
XFILLER_212_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03415_ clkbuf_0__03415_/X vssd1 vssd1 vccd1 vccd1 _14843__767/A sky130_fd_sc_hd__clkbuf_16
XFILLER_211_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11532_ _11532_/A vssd1 vssd1 vccd1 vccd1 _17719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ input79/X _14186_/D _14249_/Y vssd1 vssd1 vccd1 vccd1 _18090_/D sky130_fd_sc_hd__a21boi_2
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _11329_/X _18061_/Q _11467_/S vssd1 vssd1 vccd1 vccd1 _11464_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319__510 _14320__511/A vssd1 vssd1 vccd1 vccd1 _18145_/CLK sky130_fd_sc_hd__inv_2
X_13202_ _14083_/A vssd1 vssd1 vccd1 vccd1 _16056_/A sky130_fd_sc_hd__buf_12
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _10406_/B _10417_/A _10407_/X vssd1 vssd1 vccd1 vccd1 _10414_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_104_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128__842 _15128__842/A vssd1 vssd1 vccd1 vccd1 _18518_/CLK sky130_fd_sc_hd__inv_2
X_14182_ _16690_/A vssd1 vssd1 vccd1 vccd1 _14184_/A sky130_fd_sc_hd__buf_6
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11394_ _11335_/X _18118_/Q _11394_/S vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13133_ _13354_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10345_ _18475_/Q vssd1 vssd1 vccd1 vccd1 _10345_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18990_ _18996_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13064_ _13049_/X _13064_/B vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__and2b_1
X_17941_ _17951_/CLK _17941_/D vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _18624_/Q _10175_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12015_ _11898_/X _11917_/X _12115_/S vssd1 vssd1 vccd1 vccd1 _12104_/A sky130_fd_sc_hd__mux2_1
X_15743__1030 _15747__1034/A vssd1 vssd1 vccd1 vccd1 _18747_/CLK sky130_fd_sc_hd__inv_2
X_17872_ _17878_/CLK _17872_/D vssd1 vssd1 vccd1 vccd1 _17872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16823_ _16894_/A vssd1 vssd1 vccd1 vccd1 _16823_/X sky130_fd_sc_hd__buf_2
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15432__927 _15433__928/A vssd1 vssd1 vccd1 vccd1 _18614_/CLK sky130_fd_sc_hd__inv_2
X_13966_ _14090_/A _13987_/B _14076_/C vssd1 vssd1 vccd1 vccd1 _13973_/A sky130_fd_sc_hd__and3_2
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16754_ _16767_/S _17783_/Q input14/X _16742_/X _16788_/A vssd1 vssd1 vccd1 vccd1
+ _16754_/X sky130_fd_sc_hd__a311o_1
XFILLER_235_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12917_ _12917_/A vssd1 vssd1 vccd1 vccd1 _17668_/D sky130_fd_sc_hd__clkbuf_1
X_15705_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__buf_1
XFILLER_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13897_ _13733_/A _13885_/X _13894_/X vssd1 vssd1 vccd1 vccd1 _13897_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18424_ _18424_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
X_12848_ _17646_/Q _13085_/B vssd1 vssd1 vccd1 vccd1 _12849_/D sky130_fd_sc_hd__xor2_1
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15636_ _16056_/A _15638_/B vssd1 vssd1 vccd1 vccd1 _18663_/D sky130_fd_sc_hd__nor2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _15572_/B _15572_/C vssd1 vssd1 vccd1 vccd1 _15571_/B sky130_fd_sc_hd__and2_1
X_18355_ _18355_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12779_ _17636_/Q _17999_/Q _12862_/B vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17306_ _17357_/S vssd1 vssd1 vccd1 vccd1 _17381_/B sky130_fd_sc_hd__clkbuf_2
X_14518_ _14524_/A vssd1 vssd1 vccd1 vccd1 _14518_/X sky130_fd_sc_hd__buf_1
XFILLER_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15498_ _15585_/B _15499_/B vssd1 vssd1 vccd1 vccd1 _15498_/Y sky130_fd_sc_hd__nand2_1
X_18286_ _18286_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17237_ _19253_/Q _17237_/B _17237_/C _17237_/D vssd1 vssd1 vccd1 vccd1 _17250_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03975_ _15717_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03975_/X sky130_fd_sc_hd__clkbuf_16
X_14449_ _14449_/A vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__buf_1
XFILLER_128_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179__455 _14252__456/A vssd1 vssd1 vccd1 vccd1 _18063_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17168_ _17169_/B _17169_/C _17167_/Y vssd1 vssd1 vccd1 vccd1 _19233_/D sky130_fd_sc_hd__a21oi_1
XFILLER_190_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16119_ _16290_/S vssd1 vssd1 vccd1 vccd1 _16119_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _17776_/Q _17775_/Q _17773_/Q _12095_/A vssd1 vssd1 vccd1 vccd1 _17099_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09990_ _18768_/Q _09963_/X _09992_/S vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08941_ _09697_/A vssd1 vssd1 vccd1 vccd1 _08941_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04527_ _16543_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04527_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08872_ _19313_/Q _08871_/X _08878_/S vssd1 vssd1 vccd1 vccd1 _08873_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03409_ _14809_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03409_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09424_ _08929_/X _19054_/Q _09424_/S vssd1 vssd1 vccd1 vccd1 _09425_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09355_ _09355_/A vssd1 vssd1 vccd1 vccd1 _19084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09286_ _09286_/A vssd1 vssd1 vccd1 vccd1 _19119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10130_ _10129_/X _18713_/Q _10136_/S vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__mux2_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _18739_/Q _10060_/X _10064_/S vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__mux2_1
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03964_ clkbuf_0__03964_/X vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__clkbuf_16
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _13820_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ _17894_/Q _13738_/X _13750_/Y _13741_/X vssd1 vssd1 vccd1 vccd1 _17894_/D
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_109 _19386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _08883_/X _18292_/Q hold9/X vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12702_ _12707_/A _12700_/A _12695_/X vssd1 vssd1 vccd1 vccd1 _12703_/B sky130_fd_sc_hd__o21ai_1
XFILLER_204_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16470_ _16467_/X _16468_/Y _16469_/X vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__a21oi_1
X_13682_ _13688_/A vssd1 vssd1 vccd1 vccd1 _13682_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_243_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10894_ _10894_/A vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15881__175 _15882__176/A vssd1 vssd1 vccd1 vccd1 _18850_/CLK sky130_fd_sc_hd__inv_2
X_15685__984 _15685__984/A vssd1 vssd1 vccd1 vccd1 _18701_/CLK sky130_fd_sc_hd__inv_2
XFILLER_204_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12633_ _12633_/A vssd1 vssd1 vccd1 vccd1 _17598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15352_ _19322_/Q _19306_/Q _19298_/Q _19273_/Q _15293_/X _15215_/X vssd1 vssd1 vccd1
+ vccd1 _15352_/X sky130_fd_sc_hd__mux4_2
X_18140_ _18140_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ _17592_/Q vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__04378_ clkbuf_0__04378_/X vssd1 vssd1 vccd1 vccd1 _16542__254/A sky130_fd_sc_hd__clkbuf_16
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ _18038_/Q _11326_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18071_ _18072_/CLK _18071_/D vssd1 vssd1 vccd1 vccd1 _18071_/Q sky130_fd_sc_hd__dfxtp_1
X_15283_ _19069_/Q _19061_/Q _19053_/Q _19007_/Q _15232_/X _15233_/X vssd1 vssd1 vccd1
+ vccd1 _15284_/A sky130_fd_sc_hd__mux4_1
X_12495_ _17591_/Q _17592_/Q _12610_/A _12394_/X _12396_/X _12397_/X vssd1 vssd1 vccd1
+ vccd1 _12495_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14234_ _18087_/Q input45/X _16997_/S vssd1 vssd1 vccd1 vccd1 _14235_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11446_ _18095_/Q _11270_/X _11448_/S vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ _11338_/X _18125_/Q _11381_/S vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03591_ clkbuf_0__03591_/X vssd1 vssd1 vccd1 vccd1 _15117__834/A sky130_fd_sc_hd__clkbuf_16
XFILLER_125_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__buf_1
XFILLER_180_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _18480_/Q vssd1 vssd1 vccd1 vccd1 _10328_/X sky130_fd_sc_hd__clkbuf_4
X_14096_ _16570_/A vssd1 vssd1 vccd1 vccd1 _14096_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _19133_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13032_/X _13047_/B vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__and2b_1
X_17924_ _19132_/CLK _17924_/D vssd1 vssd1 vccd1 vccd1 _17924_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10259_/A vssd1 vssd1 vccd1 vccd1 _18632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17855_ _18462_/CLK _17855_/D vssd1 vssd1 vccd1 vccd1 _17855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16806_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16820_/A sky130_fd_sc_hd__inv_2
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17786_ _19132_/CLK _17786_/D vssd1 vssd1 vccd1 vccd1 _17786_/Q sky130_fd_sc_hd__dfxtp_1
X_14998_ _18459_/Q _18458_/Q _14998_/C vssd1 vssd1 vccd1 vccd1 _15005_/B sky130_fd_sc_hd__and3_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16737_ _19091_/Q _16737_/B vssd1 vssd1 vccd1 vccd1 _16762_/A sky130_fd_sc_hd__nand2_2
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13949_ _13173_/X _13946_/X _13948_/Y _13937_/X vssd1 vssd1 vccd1 vccd1 _17960_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_235_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18407_ _18407_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _18670_/Q _18660_/Q _18659_/Q _18658_/Q vssd1 vssd1 vccd1 vccd1 _15619_/X
+ sky130_fd_sc_hd__and4_1
X_19387_ input6/X vssd1 vssd1 vccd1 vccd1 _19387_/X sky130_fd_sc_hd__buf_12
X_16599_ _19028_/Q _16596_/B _16598_/Y vssd1 vssd1 vccd1 vccd1 _19028_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09140_ _19182_/Q _09139_/X _09146_/S vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18338_ _18338_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_wb_clk_i _17819_/CLK vssd1 vssd1 vccd1 vccd1 _18876_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ _19199_/Q _08877_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__mux2_1
X_18269_ _18269_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09973_ _15174_/B _10424_/C vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__nand2_4
X_14153__436 _14155__438/A vssd1 vssd1 vccd1 vccd1 _18044_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ _18884_/Q vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__buf_4
XFILLER_170_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08855_ _18078_/Q _18079_/Q _08855_/C _18076_/Q vssd1 vssd1 vccd1 vccd1 _08997_/C
+ sky130_fd_sc_hd__or4b_2
XFILLER_245_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08786_ _18886_/Q vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__buf_2
XFILLER_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461__624 _14461__624/A vssd1 vssd1 vccd1 vccd1 _18259_/CLK sky130_fd_sc_hd__inv_2
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09407_ _09407_/A vssd1 vssd1 vccd1 vccd1 _19062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09338_ _09971_/A _09936_/C _10432_/A vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__or3b_4
XFILLER_200_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _19124_/Q _09268_/X _09272_/S vssd1 vssd1 vccd1 vccd1 _09270_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__04163_ clkbuf_0__04163_/X vssd1 vssd1 vccd1 vccd1 _16073__189/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11300_ _11300_/A vssd1 vssd1 vccd1 vccd1 _18156_/D sky130_fd_sc_hd__clkbuf_1
X_12280_ _12812_/A vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11231_ _11153_/X _18183_/Q _11233_/S vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11162_ _11341_/A vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__buf_2
XFILLER_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10113_ _10602_/B _10564_/B vssd1 vssd1 vccd1 vccd1 _10136_/S sky130_fd_sc_hd__or2_2
X_16644__284 _16644__284/A vssd1 vssd1 vccd1 vccd1 _19058_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ _11093_/A vssd1 vssd1 vccd1 vccd1 _18241_/D sky130_fd_sc_hd__clkbuf_1
X_15970_ _15970_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _15970_/X sky130_fd_sc_hd__or2_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14921_ _18465_/Q _17848_/Q vssd1 vssd1 vccd1 vccd1 _14936_/B sky130_fd_sc_hd__or2_1
X_10044_ _18744_/Q _09963_/X _10046_/S vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19016_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _19247_/CLK _17640_/D vssd1 vssd1 vccd1 vccd1 _17640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852_ _14852_/A vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__buf_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _13529_/X _13802_/X _13789_/X vssd1 vssd1 vccd1 vccd1 _13803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17571_ _17571_/CLK _17571_/D vssd1 vssd1 vccd1 vccd1 _17571_/Q sky130_fd_sc_hd__dfxtp_1
X_11995_ _12007_/S vssd1 vssd1 vccd1 vccd1 _11995_/X sky130_fd_sc_hd__buf_2
XFILLER_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _19310_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13734_ _17888_/Q _13719_/B _13733_/Y _13726_/X vssd1 vssd1 vccd1 vccd1 _17888_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16522_ _16522_/A _16530_/B vssd1 vssd1 vccd1 vccd1 _16523_/A sky130_fd_sc_hd__and2_1
XFILLER_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ _10946_/A vssd1 vssd1 vccd1 vccd1 _18300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14774__712 _14776__714/A vssd1 vssd1 vccd1 vccd1 _18355_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19241_ _19247_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _17864_/Q _13659_/X _13664_/Y vssd1 vssd1 vccd1 vccd1 _17864_/D sky130_fd_sc_hd__o21a_1
X_16453_ _18973_/Q _16453_/B _16453_/C vssd1 vssd1 vccd1 vccd1 _16458_/B sky130_fd_sc_hd__and3_1
XFILLER_220_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10877_ _18335_/Q _10800_/X _10879_/S vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12616_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__buf_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15404_/X sky130_fd_sc_hd__buf_1
X_19172_ _19172_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_1
X_16384_ _18979_/Q _16384_/B vssd1 vssd1 vccd1 vccd1 _16421_/B sky130_fd_sc_hd__xor2_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _17844_/Q vssd1 vssd1 vccd1 vccd1 _13596_/Y sky130_fd_sc_hd__inv_2
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__08198_ clkbuf_0__08198_/X vssd1 vssd1 vccd1 vccd1 _13108__414/A sky130_fd_sc_hd__clkbuf_16
X_15335_ _19002_/Q _18964_/Q _18956_/Q _17545_/Q _15293_/X _15215_/X vssd1 vssd1 vccd1
+ vccd1 _15335_/X sky130_fd_sc_hd__mux4_2
X_18123_ _18123_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_1
X_12547_ _12535_/X _12546_/X _12547_/S vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18054_ _18054_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
X_15266_ _15260_/X _15265_/X _09615_/A vssd1 vssd1 vccd1 vccd1 _15266_/X sky130_fd_sc_hd__o21a_1
X_12478_ _12478_/A vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14217_ _14217_/A vssd1 vssd1 vccd1 vccd1 _18079_/D sky130_fd_sc_hd__clkbuf_1
X_11429_ _11429_/A vssd1 vssd1 vccd1 vccd1 _18103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700__995 _15701__996/A vssd1 vssd1 vccd1 vccd1 _18712_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__08201_ _13116_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__08201_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_112_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _14079_/A _14083_/B vssd1 vssd1 vccd1 vccd1 _14079_/Y sky130_fd_sc_hd__nor2_2
X_18956_ _18956_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17907_ _19109_/CLK _17907_/D vssd1 vssd1 vccd1 vccd1 _17907_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18887_ _18996_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17838_ _17840_/CLK _17838_/D vssd1 vssd1 vccd1 vccd1 _17838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _17772_/CLK _17769_/D vssd1 vssd1 vccd1 vccd1 _17769_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ _11365_/A _11260_/A vssd1 vssd1 vccd1 vccd1 _09146_/S sky130_fd_sc_hd__nor2_1
XFILLER_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09054_ _18661_/Q vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _18778_/Q _09955_/X _09956_/S vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__04850_ clkbuf_0__04850_/X vssd1 vssd1 vccd1 vccd1 _17384_/A sky130_fd_sc_hd__clkbuf_16
X_08907_ _19300_/Q _08804_/X _08907_/S vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _11456_/B _11383_/B _09892_/B _09886_/X _09870_/X vssd1 vssd1 vccd1 vccd1
+ _18805_/D sky130_fd_sc_hd__o311a_1
Xclkbuf_1_0__f__03801_ clkbuf_0__03801_/X vssd1 vssd1 vccd1 vccd1 _15425__921/A sky130_fd_sc_hd__clkbuf_16
XFILLER_100_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08838_/A _09442_/A vssd1 vssd1 vccd1 vccd1 _08853_/A sky130_fd_sc_hd__nor2_1
XFILLER_246_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877__360 _11879__362/A vssd1 vssd1 vccd1 vccd1 _17507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08769_ hold14/A _08769_/B _09611_/A vssd1 vssd1 vccd1 vccd1 _08772_/A sky130_fd_sc_hd__and3_1
XFILLER_122_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11791_/B vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__buf_2
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03594_ clkbuf_0__03594_/X vssd1 vssd1 vccd1 vccd1 _15128__842/A sky130_fd_sc_hd__clkbuf_16
XFILLER_241_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10731_ _10731_/A vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14838__764 _14838__764/A vssd1 vssd1 vccd1 vccd1 _18407_/CLK sky130_fd_sc_hd__inv_2
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _17798_/Q _13457_/B vssd1 vssd1 vccd1 vccd1 _13450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10662_ _18425_/Q _09729_/X _10662_/S vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12401_ _17598_/Q vssd1 vssd1 vccd1 vccd1 _12631_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13381_ _13274_/X _13366_/S _13337_/X vssd1 vssd1 vccd1 vccd1 _13381_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10593_ _10593_/A vssd1 vssd1 vccd1 vccd1 _18488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _16216_/A _15051_/B vssd1 vssd1 vccd1 vccd1 _15052_/A sky130_fd_sc_hd__and2_1
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _12812_/A vssd1 vssd1 vccd1 vccd1 _12263_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ _13414_/A _13995_/X _13992_/X vssd1 vssd1 vccd1 vccd1 _14002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11214_ _18190_/Q _11056_/X _11214_/S vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__mux2_1
X_12194_ _17528_/Q _17489_/B vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__xor2_1
XFILLER_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18810_ _18810_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11145_ _11142_/X _18218_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__mux2_1
Xoutput84 _11772_/A vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__buf_2
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput95 _11730_/X vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _18741_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11076_ _11076_/A vssd1 vssd1 vccd1 vccd1 _18248_/D sky130_fd_sc_hd__clkbuf_1
X_15953_ _15951_/Y _15951_/B _15953_/S vssd1 vssd1 vccd1 vccd1 _15954_/C sky130_fd_sc_hd__mux2_1
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14904_ _14904_/A _14904_/B vssd1 vssd1 vccd1 vccd1 _14960_/B sky130_fd_sc_hd__xnor2_1
X_10027_ _10027_/A vssd1 vssd1 vccd1 vccd1 _18752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18672_ _18672_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _09253_/A _16052_/A _14244_/X _14095_/A vssd1 vssd1 vccd1 vccd1 _16010_/A
+ sky130_fd_sc_hd__a31o_4
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _17629_/CLK _17623_/D vssd1 vssd1 vccd1 vccd1 _17623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04011_ _15861_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04011_/X sky130_fd_sc_hd__clkbuf_16
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17554_ _17776_/CLK _17554_/D vssd1 vssd1 vccd1 vccd1 _17554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _19228_/Q vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _16514_/A _16534_/B _16298_/Y vssd1 vssd1 vccd1 vccd1 _16505_/X sky130_fd_sc_hd__o21a_1
X_13717_ _13717_/A _13719_/B vssd1 vssd1 vccd1 vccd1 _13717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _18307_/Q _10910_/X _10929_/S vssd1 vssd1 vccd1 vccd1 _10930_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17485_ _17485_/A _17485_/B _17485_/C _17485_/D vssd1 vssd1 vccd1 vccd1 _17485_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _17586_/Q _18384_/Q _18392_/Q _18426_/Q _14574_/X _14637_/X vssd1 vssd1 vccd1
+ vccd1 _14698_/B sky130_fd_sc_hd__mux4_2
XFILLER_205_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16356__247 _16358__249/A vssd1 vssd1 vccd1 vccd1 _18963_/CLK sky130_fd_sc_hd__inv_2
X_19224_ _19261_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16436_ _16471_/A vssd1 vssd1 vccd1 vccd1 _16467_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ _13761_/A _13681_/B vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__nor2_2
XFILLER_188_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19155_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_1
X_13579_ _13579_/A vssd1 vssd1 vccd1 vccd1 _17837_/D sky130_fd_sc_hd__clkbuf_1
X_16367_ _17805_/Q _16402_/B vssd1 vssd1 vccd1 vccd1 _16412_/B sky130_fd_sc_hd__or2_1
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18106_ _18106_/CLK _18106_/D vssd1 vssd1 vccd1 vccd1 _18106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04844_ _17043_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04844_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15318_ _19320_/Q _19304_/Q _19296_/Q _19271_/Q _15293_/X _15218_/X vssd1 vssd1 vccd1
+ vccd1 _15318_/X sky130_fd_sc_hd__mux4_2
X_19086_ _19086_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_1
X_16298_ _18995_/Q vssd1 vssd1 vccd1 vccd1 _16298_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15698__994 _15698__994/A vssd1 vssd1 vccd1 vccd1 _18711_/CLK sky130_fd_sc_hd__inv_2
X_18037_ _18037_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15249_ _15291_/A vssd1 vssd1 vccd1 vccd1 _15249_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14531__680 _14532__681/A vssd1 vssd1 vccd1 vccd1 _18315_/CLK sky130_fd_sc_hd__inv_2
X_09810_ _09674_/X _18827_/Q _09818_/S vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09741_ _10713_/A vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18939_ _18939_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03588_ _15094_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03588_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_246_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09672_ _18906_/Q _09280_/X _09672_/S vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15451__941 _15453__943/A vssd1 vssd1 vccd1 vccd1 _18628_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09106_ _09106_/A vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _09037_/A vssd1 vssd1 vccd1 vccd1 _19209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313__505 _14314__506/A vssd1 vssd1 vccd1 vccd1 _18140_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09939_ _09968_/S vssd1 vssd1 vccd1 vccd1 _09956_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_218_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _12950_/A vssd1 vssd1 vccd1 vccd1 _17670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ _19252_/Q _19253_/Q _11956_/S vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12881_/A vssd1 vssd1 vccd1 vccd1 _17657_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17064__51 _17066__53/A vssd1 vssd1 vccd1 vccd1 _19200_/CLK sky130_fd_sc_hd__inv_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _17907_/Q _11793_/X _11831_/X _11802_/X vssd1 vssd1 vccd1 vccd1 _11832_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14620_ _14664_/A _14618_/X _14619_/X vssd1 vssd1 vccd1 vccd1 _14620_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14551_ _14547_/X _14548_/X _14729_/S vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__mux2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11763_ _11763_/A vssd1 vssd1 vccd1 vccd1 _11763_/X sky130_fd_sc_hd__buf_2
XFILLER_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13502_ _17811_/Q _13499_/X _13501_/Y vssd1 vssd1 vccd1 vccd1 _17811_/D sky130_fd_sc_hd__o21a_1
X_10714_ _18403_/Q _10713_/X _10714_/S vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__mux2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17274_/B _17274_/C _17270_/C vssd1 vssd1 vccd1 vccd1 _17276_/B sky130_fd_sc_hd__and3_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _16578_/A _11694_/B _11694_/C vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__nor3_1
X_13433_ _14078_/A _13433_/B vssd1 vssd1 vccd1 vccd1 _17793_/D sky130_fd_sc_hd__nor2_1
X_16221_ _16278_/A _16221_/B vssd1 vssd1 vccd1 vccd1 _16221_/Y sky130_fd_sc_hd__nor2_1
X_10645_ _10645_/A vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16152_ _16152_/A vssd1 vssd1 vccd1 vccd1 _16289_/S sky130_fd_sc_hd__buf_2
X_13364_ _13361_/X _13355_/X _13363_/Y _13359_/X vssd1 vssd1 vccd1 vccd1 _17776_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10576_ _10129_/X _18494_/Q _10580_/S vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__mux2_1
X_14886__802 _14886__802/A vssd1 vssd1 vccd1 vccd1 _18447_/CLK sky130_fd_sc_hd__inv_2
XFILLER_155_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _12315_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12316_/D sky130_fd_sc_hd__nor2_1
XFILLER_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13295_ _17757_/Q _13280_/X _13294_/Y vssd1 vssd1 vccd1 vccd1 _17757_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15034_ _15034_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15035_/A sky130_fd_sc_hd__and2_1
XFILLER_154_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12246_ _17549_/Q _18028_/Q _12318_/B vssd1 vssd1 vccd1 vccd1 _12247_/B sky130_fd_sc_hd__mux2_1
XFILLER_177_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_91_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18477_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__03411_ clkbuf_0__03411_/X vssd1 vssd1 vccd1 vccd1 _14824__752/A sky130_fd_sc_hd__clkbuf_16
X_12177_ _12166_/X _12177_/B vssd1 vssd1 vccd1 vccd1 _12178_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_20_wb_clk_i _17526_/CLK vssd1 vssd1 vccd1 vccd1 _17881_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _18225_/Q _11047_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _11129_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16985_ _18186_/Q _18178_/Q _18170_/Q _18162_/Q _16827_/X _16828_/X vssd1 vssd1 vccd1
+ vccd1 _16986_/B sky130_fd_sc_hd__mux4_1
XFILLER_111_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18724_ _18724_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15936_ _15936_/A _15936_/B _15936_/C _15936_/D vssd1 vssd1 vccd1 vccd1 _15945_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11059_ _18663_/Q vssd1 vssd1 vccd1 vccd1 _11059_/X sky130_fd_sc_hd__buf_2
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__05012_ clkbuf_0__05012_/X vssd1 vssd1 vccd1 vccd1 _17383__79/A sky130_fd_sc_hd__clkbuf_16
X_18655_ _18655_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17606_ _17611_/CLK _17606_/D vssd1 vssd1 vccd1 vccd1 _17606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _18586_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16657__294 _16657__294/A vssd1 vssd1 vccd1 vccd1 _19068_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _17537_/CLK _17537_/D vssd1 vssd1 vccd1 vccd1 _17537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17468_ _17739_/Q _19337_/Q _17468_/S vssd1 vssd1 vccd1 vccd1 _17469_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19207_ _19207_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
X_16419_ _16419_/A _16419_/B _16419_/C _16419_/D vssd1 vssd1 vccd1 vccd1 _16420_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_220_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19138_ _19144_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15759__1043 _15760__1044/A vssd1 vssd1 vccd1 vccd1 _18760_/CLK sky130_fd_sc_hd__inv_2
XFILLER_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19069_ _19069_/CLK _19069_/D vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfxtp_1
X_14787__722 _14789__724/A vssd1 vssd1 vccd1 vccd1 _18365_/CLK sky130_fd_sc_hd__inv_2
XFILLER_218_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__04589_ clkbuf_0__04589_/X vssd1 vssd1 vccd1 vccd1 _17006_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09724_ _18859_/Q _09723_/X _09733_/S vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13104__410 _13106__412/A vssd1 vssd1 vccd1 vccd1 _17706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _09975_/C _10424_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10546_/B sky130_fd_sc_hd__nand3_4
XFILLER_216_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09586_/A vssd1 vssd1 vccd1 vccd1 _18941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ _10424_/B _10424_/C _10433_/C vssd1 vssd1 vccd1 vccd1 _10430_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14538__686 _14539__687/A vssd1 vssd1 vccd1 vccd1 _18321_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10361_ _10361_/A vssd1 vssd1 vccd1 vccd1 _18590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12100_ _19262_/Q _19263_/Q _19264_/Q _19265_/Q _11995_/X _11938_/A vssd1 vssd1 vccd1
+ vccd1 _12100_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _17695_/Q _12920_/X _12921_/A _17694_/Q vssd1 vssd1 vccd1 vccd1 _13087_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_174_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10292_ _10456_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10308_/S sky130_fd_sc_hd__nor2_2
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12031_ _11925_/X _11908_/X _12032_/S vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__mux2_1
X_15458__947 _15460__949/A vssd1 vssd1 vccd1 vccd1 _18634_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14881__798 _14881__798/A vssd1 vssd1 vccd1 vccd1 _18443_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16770_ _16775_/A _16770_/B vssd1 vssd1 vccd1 vccd1 _19131_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _17973_/Q _13968_/X _13981_/Y vssd1 vssd1 vccd1 vccd1 _17973_/D sky130_fd_sc_hd__o21a_1
XFILLER_120_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _17653_/Q _12850_/X _12932_/X _17656_/Q vssd1 vssd1 vccd1 vccd1 _12933_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18440_ _18440_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12915_/S vssd1 vssd1 vccd1 vccd1 _12944_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15845__146 _15846__147/A vssd1 vssd1 vccd1 vccd1 _18821_/CLK sky130_fd_sc_hd__inv_2
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14598_/X _14601_/X _14726_/S vssd1 vssd1 vccd1 vccd1 _14603_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11815_ _11815_/A vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__buf_2
X_18371_ _18371_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12812_/A vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15583_ _15583_/A vssd1 vssd1 vccd1 vccd1 _15611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17322_ _17322_/A vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11746_ _17860_/Q _17531_/Q _17770_/Q vssd1 vssd1 vccd1 vccd1 _11747_/A sky130_fd_sc_hd__mux2_8
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16730__344 _16730__344/A vssd1 vssd1 vccd1 vccd1 _19123_/CLK sky130_fd_sc_hd__inv_2
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17253_ _17258_/C _17265_/B _17253_/C vssd1 vssd1 vccd1 vccd1 _17254_/A sky130_fd_sc_hd__and3b_1
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11677_ _13892_/A vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__03991_ _15793_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03991_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ _18746_/Q _18754_/Q _18762_/Q _18770_/Q _16127_/X _16128_/X vssd1 vssd1 vccd1
+ vccd1 _16204_/X sky130_fd_sc_hd__mux4_1
X_13416_ _13271_/X _13395_/X _13408_/X vssd1 vssd1 vccd1 vccd1 _13416_/Y sky130_fd_sc_hd__a21oi_1
X_10628_ _18441_/Q _10123_/A _10630_/S vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__mux2_1
X_17184_ _17186_/B _17184_/B vssd1 vssd1 vccd1 vccd1 _17184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13347_ input72/X _16518_/B _13330_/X _13346_/X _13343_/X vssd1 vssd1 vccd1 vccd1
+ _17774_/D sky130_fd_sc_hd__a311o_1
XFILLER_155_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16135_ _18914_/Q _16098_/X _16134_/Y _14247_/X vssd1 vssd1 vccd1 vccd1 _18914_/D
+ sky130_fd_sc_hd__o211a_1
X_10559_ _10559_/A vssd1 vssd1 vccd1 vccd1 _18502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ _13645_/A _13278_/B vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__nor2_2
X_16066_ _16049_/A _16064_/C _15993_/B _16010_/A vssd1 vssd1 vccd1 vccd1 _18889_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15017_ _18462_/Q _14978_/X _15016_/X vssd1 vssd1 vccd1 vccd1 _15018_/B sky130_fd_sc_hd__a21oi_1
X_12229_ _12229_/A vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__buf_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__04374_ clkbuf_0__04374_/X vssd1 vssd1 vccd1 vccd1 _16543_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16968_ _18217_/Q _18201_/Q _18490_/Q _18193_/Q _09852_/A _09858_/A vssd1 vssd1 vccd1
+ vccd1 _16968_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18707_ _18707_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_1
X_15919_ _15927_/A _17824_/Q _17823_/Q vssd1 vssd1 vccd1 vccd1 _15929_/B sky130_fd_sc_hd__or3_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16899_ _18059_/Q _18051_/Q _18043_/Q _18035_/Q _16870_/X _16871_/X vssd1 vssd1 vccd1
+ vccd1 _16899_/X sky130_fd_sc_hd__mux4_2
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09440_ _09440_/A _09440_/B vssd1 vssd1 vccd1 vccd1 _09441_/D sky130_fd_sc_hd__nand2_1
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18638_ _18638_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03187_ clkbuf_0__03187_/X vssd1 vssd1 vccd1 vccd1 _14476__636/A sky130_fd_sc_hd__clkbuf_16
XFILLER_227_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ _19077_/Q _09108_/X _09375_/S vssd1 vssd1 vccd1 vccd1 _09372_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18569_ _18572_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03980_ clkbuf_0__03980_/X vssd1 vssd1 vccd1 vccd1 _15746__1033/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_3 _17112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09707_ _09707_/A vssd1 vssd1 vccd1 vccd1 _18895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09638_ _10219_/A _09636_/Y _09637_/Y vssd1 vssd1 vccd1 vccd1 _18929_/D sky130_fd_sc_hd__o21a_1
XFILLER_215_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09569_ _09569_/A vssd1 vssd1 vccd1 vccd1 _18948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11600_ _11600_/A vssd1 vssd1 vccd1 vccd1 _17573_/D sky130_fd_sc_hd__clkbuf_1
X_12580_ _12580_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__or2_1
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__03414_ clkbuf_0__03414_/X vssd1 vssd1 vccd1 vccd1 _14852_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_90_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11531_ _08830_/X _17719_/Q _11539_/S vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14250_ input79/X _11865_/B _14249_/Y vssd1 vssd1 vccd1 vccd1 _18089_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11462_ _11462_/A vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ _13374_/A vssd1 vssd1 vccd1 vccd1 _14083_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10413_ _10413_/A vssd1 vssd1 vccd1 vccd1 _18567_/D sky130_fd_sc_hd__clkbuf_1
X_14181_ _14186_/D _14249_/A vssd1 vssd1 vccd1 vccd1 _18064_/D sky130_fd_sc_hd__nor2_4
X_11393_ _11393_/A vssd1 vssd1 vccd1 vccd1 _18119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13132_ _13873_/D _13132_/B _13873_/B vssd1 vssd1 vccd1 vccd1 _13133_/B sky130_fd_sc_hd__or3b_4
X_10344_ _10344_/A vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17940_ _18024_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_1
X_13063_ _17940_/Q _17698_/Q _13070_/S vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__mux2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10275_ _10290_/S vssd1 vssd1 vccd1 vccd1 _10284_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12014_ _17779_/Q vssd1 vssd1 vccd1 vccd1 _12115_/S sky130_fd_sc_hd__inv_2
XFILLER_215_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17871_ _17878_/CLK _17871_/D vssd1 vssd1 vccd1 vccd1 _17871_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16822_ _16881_/A vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__buf_2
XFILLER_215_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16753_ _19110_/Q _17788_/Q _16744_/X vssd1 vssd1 vccd1 vccd1 _16788_/A sky130_fd_sc_hd__o21ai_2
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13965_ _16054_/A _13950_/B _13964_/Y _11697_/X vssd1 vssd1 vccd1 vccd1 _17967_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14326__515 _14330__519/A vssd1 vssd1 vccd1 vccd1 _18150_/CLK sky130_fd_sc_hd__inv_2
XFILLER_235_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12916_ _12911_/X _12916_/B vssd1 vssd1 vccd1 vccd1 _12917_/A sky130_fd_sc_hd__and2b_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758__1042 _15758__1042/A vssd1 vssd1 vccd1 vccd1 _18759_/CLK sky130_fd_sc_hd__inv_2
X_13896_ _17941_/Q _13879_/X _13895_/Y vssd1 vssd1 vccd1 vccd1 _17941_/D sky130_fd_sc_hd__o21a_1
XFILLER_111_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18423_ _18423_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15635_ _16055_/A _15638_/B vssd1 vssd1 vccd1 vccd1 _18662_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _17649_/Q _13090_/B vssd1 vssd1 vccd1 vccd1 _12849_/C sky130_fd_sc_hd__xor2_1
XFILLER_222_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18354_ _18354_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
X_15566_ _15572_/B _15572_/C vssd1 vssd1 vccd1 vccd1 _15568_/B sky130_fd_sc_hd__nor2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12778_ _12831_/S vssd1 vssd1 vccd1 vccd1 _12862_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17305_ _17772_/Q _17423_/B vssd1 vssd1 vccd1 vccd1 _17357_/S sky130_fd_sc_hd__and2_2
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11729_ _11717_/X _17932_/Q vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__and2b_4
X_18285_ _18285_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15497_ _17834_/Q _15501_/A vssd1 vssd1 vccd1 vccd1 _15499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ _17236_/A vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03974_ _15711_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03974_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_163_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17167_ _17169_/B _17169_/C _17126_/X vssd1 vssd1 vccd1 vccd1 _17167_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _18445_/Q _19083_/Q _19120_/Q _18429_/Q _16117_/X _10420_/X vssd1 vssd1 vccd1
+ vccd1 _16118_/X sky130_fd_sc_hd__mux4_2
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17098_ _17098_/A vssd1 vssd1 vccd1 vccd1 _17098_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08940_ _18880_/Q vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__buf_2
X_16049_ _16049_/A _18888_/Q _16049_/C _16049_/D vssd1 vssd1 vccd1 vccd1 _16050_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_233_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08871_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _08871_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_233_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__03408_ _14808_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03408_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_238_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _09423_/A vssd1 vssd1 vccd1 vccd1 _19055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09354_ _19084_/Q _09277_/X _09356_/S vssd1 vssd1 vccd1 vccd1 _09355_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09285_ _19119_/Q _08944_/X _09293_/S vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14832__759 _14832__759/A vssd1 vssd1 vccd1 vccd1 _18402_/CLK sky130_fd_sc_hd__inv_2
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15794__115 _15796__117/A vssd1 vssd1 vccd1 vccd1 _18787_/CLK sky130_fd_sc_hd__inv_2
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _10123_/A vssd1 vssd1 vccd1 vccd1 _10060_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03963_ clkbuf_0__03963_/X vssd1 vssd1 vccd1 vccd1 _15657__961/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_13_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_79_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13750_ _13750_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10962_ _10962_/A vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ _12707_/A _12707_/B _12707_/C vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__and3_1
XFILLER_141_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _13681_/A _13681_/B vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__nor2_1
X_10893_ _18321_/Q _10892_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _12641_/D _12759_/A _12632_/C vssd1 vssd1 vccd1 vccd1 _12633_/A sky130_fd_sc_hd__and3b_1
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12563_ _18013_/Q _12563_/B _12563_/C _12563_/D vssd1 vssd1 vccd1 vccd1 _12563_/X
+ sky130_fd_sc_hd__and4_1
X_13117__420 _13120__423/A vssd1 vssd1 vccd1 vccd1 _17716_/CLK sky130_fd_sc_hd__inv_2
X_15351_ _19118_/Q _18949_/Q _18607_/Q _19347_/Q _15251_/X _15291_/X vssd1 vssd1 vccd1
+ vccd1 _15351_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__04377_ clkbuf_0__04377_/X vssd1 vssd1 vccd1 vccd1 _16358__249/A sky130_fd_sc_hd__clkbuf_16
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11514_ _11514_/A vssd1 vssd1 vccd1 vccd1 _18039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18070_ _18072_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
X_12494_ _12437_/X _12439_/X _12556_/A vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__mux2_1
X_15282_ _19214_/Q _19102_/Q _18285_/Q _19094_/Q _15230_/X _09631_/X vssd1 vssd1 vccd1
+ vccd1 _15282_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14233_ _14233_/A vssd1 vssd1 vccd1 vccd1 _18086_/D sky130_fd_sc_hd__clkbuf_1
X_11445_ _11445_/A vssd1 vssd1 vccd1 vccd1 _18096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11376_ _11376_/A vssd1 vssd1 vccd1 vccd1 _18126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03590_ clkbuf_0__03590_/X vssd1 vssd1 vccd1 vccd1 _15109__827/A sky130_fd_sc_hd__clkbuf_16
X_10327_ _10327_/A vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__clkbuf_1
X_14095_ _14095_/A vssd1 vssd1 vccd1 vccd1 _16570_/A sky130_fd_sc_hd__buf_2
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18972_ _19133_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _17945_/Q _17693_/Q _13053_/S vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__mux2_1
X_17923_ _17923_/CLK _17923_/D vssd1 vssd1 vccd1 vccd1 _17923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _18632_/Q _10175_/X _10266_/S vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17854_ _17935_/CLK _17854_/D vssd1 vssd1 vccd1 vccd1 _17854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15395__897 _15395__897/A vssd1 vssd1 vccd1 vccd1 _18584_/CLK sky130_fd_sc_hd__inv_2
X_10189_ _18476_/Q vssd1 vssd1 vccd1 vccd1 _10189_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16805_ _18147_/Q _18139_/Q _18131_/Q _18275_/Q _16803_/X _16804_/X vssd1 vssd1 vccd1
+ vccd1 _16805_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17785_ _19128_/CLK _17785_/D vssd1 vssd1 vccd1 vccd1 _17785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14997_ _18458_/Q _14998_/C _18459_/Q vssd1 vssd1 vccd1 vccd1 _14999_/A sky130_fd_sc_hd__a21oi_1
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16736_ _16736_/A vssd1 vssd1 vccd1 vccd1 _16775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ _17960_/Q _13950_/B vssd1 vssd1 vccd1 vccd1 _13948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13879_ _13885_/A vssd1 vssd1 vccd1 vccd1 _13879_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18406_ _18406_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15618_ _18670_/Q vssd1 vssd1 vccd1 vccd1 _15618_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19386_ input1/X vssd1 vssd1 vccd1 vccd1 _19386_/X sky130_fd_sc_hd__buf_8
X_16598_ _19028_/Q _16596_/B _16564_/X vssd1 vssd1 vccd1 vccd1 _16598_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18337_ _18337_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ _15557_/B _15557_/C vssd1 vssd1 vccd1 vccd1 _15551_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09070_ _09070_/A vssd1 vssd1 vccd1 vccd1 _19200_/D sky130_fd_sc_hd__clkbuf_1
X_18268_ _18268_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
X_17219_ _17219_/A vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18199_ _18199_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09972_ _09972_/A _10436_/A vssd1 vssd1 vccd1 vccd1 _10424_/C sky130_fd_sc_hd__and2_2
X_16704__327 _16704__327/A vssd1 vssd1 vccd1 vccd1 _19102_/CLK sky130_fd_sc_hd__inv_2
XFILLER_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08923_ _08923_/A vssd1 vssd1 vccd1 vccd1 _19297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08854_ _19014_/Q _09084_/C vssd1 vssd1 vccd1 vccd1 _08860_/A sky130_fd_sc_hd__and2_1
XFILLER_112_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08785_ _08785_/A vssd1 vssd1 vccd1 vccd1 _19348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09406_ _08929_/X _19062_/Q _09406_/S vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09337_ _09337_/A vssd1 vssd1 vccd1 vccd1 _19092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15802__122 _15804__124/A vssd1 vssd1 vccd1 vccd1 _18794_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09268_ _18477_/Q vssd1 vssd1 vccd1 vccd1 _09268_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__04162_ clkbuf_0__04162_/X vssd1 vssd1 vccd1 vccd1 _16086_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09199_ _09199_/A vssd1 vssd1 vccd1 vccd1 _19158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11230_/A vssd1 vssd1 vccd1 vccd1 _18184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757__1041 _15758__1042/A vssd1 vssd1 vccd1 vccd1 _18758_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11161_ _11161_/A vssd1 vssd1 vccd1 vccd1 _18213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10112_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _09031_/X _18241_/Q _11098_/S vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__mux2_1
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _18463_/Q _14920_/B vssd1 vssd1 vccd1 vccd1 _14960_/C sky130_fd_sc_hd__xnor2_1
X_10043_ _10043_/A vssd1 vssd1 vccd1 vccd1 _18745_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13802_ _13802_/A vssd1 vssd1 vccd1 vccd1 _13802_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _17570_/CLK _17570_/D vssd1 vssd1 vccd1 vccd1 _17570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11994_ _11956_/X _11993_/X _12036_/S vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16521_ _16521_/A vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__clkbuf_1
X_13733_ _13733_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13733_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10945_ _18300_/Q _10907_/X hold16/A vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19248_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19240_ _19240_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15171__877 _15172__878/A vssd1 vssd1 vccd1 vccd1 _18553_/CLK sky130_fd_sc_hd__inv_2
XFILLER_204_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16452_ _16453_/B _16453_/C _18973_/Q vssd1 vssd1 vccd1 vccd1 _16454_/B sky130_fd_sc_hd__a21oi_1
XFILLER_177_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13664_ _13285_/X _13660_/X _13661_/X vssd1 vssd1 vccd1 vccd1 _13664_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10876_ _10876_/A vssd1 vssd1 vccd1 vccd1 _18336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12615_ _12630_/C vssd1 vssd1 vccd1 vccd1 _12622_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _19171_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_1
X_16094__206 _16307__209/A vssd1 vssd1 vccd1 vccd1 _18911_/CLK sky130_fd_sc_hd__inv_2
XFILLER_223_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _16383_/A _16383_/B vssd1 vssd1 vccd1 vccd1 _16384_/B sky130_fd_sc_hd__nand2_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13595_ _14078_/A _13595_/B vssd1 vssd1 vccd1 vccd1 _17843_/D sky130_fd_sc_hd__nor2_1
X_16651__289 _16651__289/A vssd1 vssd1 vccd1 vccd1 _19063_/CLK sky130_fd_sc_hd__inv_2
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14438__605 _14440__607/A vssd1 vssd1 vccd1 vccd1 _18240_/CLK sky130_fd_sc_hd__inv_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18122_ _18122_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15334_ _19117_/Q _18948_/Q _18606_/Q _19346_/Q _15245_/X _15291_/X vssd1 vssd1 vccd1
+ vccd1 _15334_/X sky130_fd_sc_hd__mux4_1
X_12546_ _12746_/A _17633_/Q _17634_/Q _17635_/Q _12396_/X _12397_/X vssd1 vssd1 vccd1
+ vccd1 _12546_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18053_ _18053_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
X_15265_ _15220_/X _15261_/X _15264_/X _15222_/X vssd1 vssd1 vccd1 vccd1 _15265_/X
+ sky130_fd_sc_hd__o211a_1
X_12477_ _12379_/X _12360_/X _12547_/S vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14216_ _18079_/Q input37/X _14218_/S vssd1 vssd1 vccd1 vccd1 _14217_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11428_ _18103_/Q _11270_/X _11430_/S vssd1 vssd1 vccd1 vccd1 _11429_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11359_ _18133_/Q _11276_/X _11363_/S vssd1 vssd1 vccd1 vccd1 _11360_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__08200_ _13110_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__08200_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14781__717 _14782__718/A vssd1 vssd1 vccd1 vccd1 _18360_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14078_ _14078_/A _14078_/B vssd1 vssd1 vccd1 vccd1 _18008_/D sky130_fd_sc_hd__nor2_1
X_18955_ _18955_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13029_ _17950_/Q _17688_/Q _13099_/B vssd1 vssd1 vccd1 vccd1 _13030_/B sky130_fd_sc_hd__mux2_1
X_17906_ _17922_/CLK _17906_/D vssd1 vssd1 vccd1 vccd1 _17906_/Q sky130_fd_sc_hd__dfxtp_4
X_18886_ _18886_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ _18462_/CLK _17837_/D vssd1 vssd1 vccd1 vccd1 _17837_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17768_ _19340_/CLK _17768_/D vssd1 vssd1 vccd1 vccd1 _17768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16719_ _17000_/A vssd1 vssd1 vccd1 vccd1 _16719_/X sky130_fd_sc_hd__buf_1
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17699_ _17951_/CLK _17699_/D vssd1 vssd1 vccd1 vccd1 _17699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17388__83 _17389__84/A vssd1 vssd1 vccd1 vccd1 _19296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _11493_/A vssd1 vssd1 vccd1 vccd1 _11260_/A sky130_fd_sc_hd__buf_4
XFILLER_37_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15445__938 _15446__939/A vssd1 vssd1 vccd1 vccd1 _18625_/CLK sky130_fd_sc_hd__inv_2
XFILLER_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09053_ _09053_/A vssd1 vssd1 vccd1 vccd1 _19205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _10126_/A vssd1 vssd1 vccd1 vccd1 _09955_/X sky130_fd_sc_hd__clkbuf_2
X_08906_ _08906_/A vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03800_ clkbuf_0__03800_/X vssd1 vssd1 vccd1 vccd1 _15422__919/A sky130_fd_sc_hd__clkbuf_16
XFILLER_246_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09011_/A _09894_/B _11383_/A vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__a21o_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _19048_/Q hold7/A vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__xor2_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17076__60 _17078__62/A vssd1 vssd1 vccd1 vccd1 _19209_/CLK sky130_fd_sc_hd__inv_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _18932_/Q hold4/A vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__xnor2_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03593_ clkbuf_0__03593_/X vssd1 vssd1 vccd1 vccd1 _15149_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_202_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10730_ _18396_/Q _10710_/X _10732_/S vssd1 vssd1 vccd1 vccd1 _10731_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12346__405 _12348__407/A vssd1 vssd1 vccd1 vccd1 _17586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_159_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10661_ _10661_/A vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ _17597_/Q vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13380_ _17782_/Q vssd1 vssd1 vccd1 vccd1 _17117_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10592_ _09039_/X _18488_/Q _10594_/S vssd1 vssd1 vccd1 vccd1 _10593_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ _12918_/A vssd1 vssd1 vccd1 vccd1 _12812_/A sky130_fd_sc_hd__clkbuf_4
X_15050_ _15026_/X _15048_/Y _15049_/X _14978_/X _18468_/Q vssd1 vssd1 vccd1 vccd1
+ _15051_/B sky130_fd_sc_hd__a32o_1
X_11884__365 _12222__369/A vssd1 vssd1 vccd1 vccd1 _17512_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14001_ _17980_/Q _13988_/X _14000_/Y vssd1 vssd1 vccd1 vccd1 _17980_/D sky130_fd_sc_hd__o21a_1
X_11213_ _11213_/A vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ _17527_/Q _17492_/B vssd1 vssd1 vccd1 vccd1 _12198_/A sky130_fd_sc_hd__xor2_1
XFILLER_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11144_ _11166_/S vssd1 vssd1 vccd1 vccd1 _11157_/S sky130_fd_sc_hd__clkbuf_2
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 _11769_/X vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__buf_2
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 _11726_/X vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__buf_2
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14845__769 _14845__769/A vssd1 vssd1 vccd1 vccd1 _18414_/CLK sky130_fd_sc_hd__inv_2
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _18740_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11075_ _09035_/X _18248_/Q _11079_/S vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__mux2_1
X_15952_ _15949_/Y _17811_/Q _15951_/A _18876_/Q vssd1 vssd1 vccd1 vccd1 _15953_/S
+ sky130_fd_sc_hd__o22a_1
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14903_ _17845_/Q _14913_/B vssd1 vssd1 vccd1 vccd1 _14904_/B sky130_fd_sc_hd__nor2_1
X_10026_ _18752_/Q _09963_/X _10028_/S vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _18671_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15883_ _15955_/A vssd1 vssd1 vccd1 vccd1 _16036_/A sky130_fd_sc_hd__inv_2
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17622_ _17629_/CLK _17622_/D vssd1 vssd1 vccd1 vccd1 _17622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04010_ _15855_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04010_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17553_ _17772_/CLK _17553_/D vssd1 vssd1 vccd1 vccd1 _17553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _14771_/A vssd1 vssd1 vccd1 vccd1 _14765_/X sky130_fd_sc_hd__buf_1
X_11977_ _11975_/X _11976_/X _11977_/S vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ _18984_/Q vssd1 vssd1 vccd1 vccd1 _16511_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_232_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13716_ _13735_/B vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17484_ _19330_/Q _12202_/A _12204_/X _19331_/Q _17483_/X vssd1 vssd1 vccd1 vccd1
+ _17485_/D sky130_fd_sc_hd__o221a_1
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10928_ _10928_/A vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ _14696_/A _14696_/B vssd1 vssd1 vccd1 vccd1 _14696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19223_ _19252_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16435_ _16464_/A _16435_/B vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__nor2_1
X_13647_ _16688_/B _13704_/B vssd1 vssd1 vccd1 vccd1 _13681_/B sky130_fd_sc_hd__nand2_2
XFILLER_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10859_ _18343_/Q _10800_/X _10861_/S vssd1 vssd1 vccd1 vccd1 _10860_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19154_ _19154_/CLK _19154_/D vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _17808_/Q _17807_/Q _17806_/Q vssd1 vssd1 vccd1 vccd1 _16402_/B sky130_fd_sc_hd__or3_1
XFILLER_160_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13578_ _13629_/A _13578_/B vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__or2_1
X_18105_ _18105_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__04843_ _17037_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__04843_/X sky130_fd_sc_hd__clkbuf_16
X_15317_ _19116_/Q _18947_/Q _18605_/Q _19345_/Q _15245_/X _15291_/X vssd1 vssd1 vccd1
+ vccd1 _15317_/X sky130_fd_sc_hd__mux4_1
X_12529_ _12529_/A vssd1 vssd1 vccd1 vccd1 _12529_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19085_ _19085_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16297_ _18996_/Q vssd1 vssd1 vccd1 vccd1 _16506_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18036_ _18036_/CLK _18036_/D vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
X_15248_ _15273_/A vssd1 vssd1 vccd1 vccd1 _15248_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15179_ _18669_/Q vssd1 vssd1 vccd1 vccd1 _15642_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09740_ _09740_/A vssd1 vssd1 vccd1 vccd1 _18854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18938_ _18938_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03587_ _15093_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__03587_/X sky130_fd_sc_hd__clkbuf_16
.ends

