VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Blink
  CLASS BLOCK ;
  FOREIGN Blink ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 200.000 150.240 ;
    END
  END blink[0]
  PIN blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.680 200.000 50.280 ;
    END
  END blink[1]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 6.990 10.640 190.350 187.920 ;
      LAYER met3 ;
        RECT 4.000 150.640 196.000 187.845 ;
        RECT 4.400 149.240 195.600 150.640 ;
        RECT 4.000 50.680 196.000 149.240 ;
        RECT 4.400 49.280 195.600 50.680 ;
        RECT 4.000 10.715 196.000 49.280 ;
      LAYER met4 ;
        RECT 95.975 49.815 97.440 115.425 ;
        RECT 99.840 49.815 115.625 115.425 ;
  END
END Blink
END LIBRARY

