VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Art
  CLASS BLOCK ;
  FOREIGN Art ;
  ORIGIN -0.200 0.000 ;
  SIZE 302.920 BY 750.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.20000 0.00000 1.80000 750.00000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 298.20000 0.00000 299.80000 750.00000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.000 30.000 105.000 70.000 ;
        RECT 5.000 5.000 25.000 25.000 ;
      LAYER met1 ;
        RECT 85.000 60.000 105.000 70.120 ;
        RECT 65.000 50.000 105.000 60.000 ;
        RECT 45.000 40.000 105.000 50.000 ;
        RECT 25.000 30.120 105.000 40.000 ;
        RECT 25.000 30.000 85.000 30.120 ;
        RECT 25.000 5.000 45.000 25.000 ;
      LAYER met2 ;
        POLYGON 155.010 191.730 155.010 191.305 140.290 191.305 ;
        POLYGON 155.010 191.730 169.730 191.305 155.010 191.305 ;
        POLYGON 250.010 191.730 250.010 191.305 235.290 191.305 ;
        POLYGON 250.010 191.730 264.730 191.305 250.010 191.305 ;
        POLYGON 140.290 191.305 140.290 190.380 133.705 190.380 ;
        RECT 140.290 190.380 169.730 191.305 ;
        POLYGON 169.730 191.305 176.315 190.380 169.730 190.380 ;
        POLYGON 235.290 191.305 235.290 190.380 228.705 190.380 ;
        RECT 235.290 190.380 264.730 191.305 ;
        POLYGON 264.730 191.305 271.315 190.380 264.730 190.380 ;
        POLYGON 133.705 190.380 133.705 189.240 127.370 189.240 ;
        RECT 133.705 189.240 176.315 190.380 ;
        POLYGON 176.315 190.380 182.645 189.240 176.315 189.240 ;
        POLYGON 228.705 190.380 228.705 189.240 222.370 189.240 ;
        RECT 228.705 189.240 271.315 190.380 ;
        POLYGON 271.315 190.380 277.645 189.240 271.315 189.240 ;
        POLYGON 127.370 189.240 127.370 187.890 121.255 187.890 ;
        RECT 127.370 187.890 182.645 189.240 ;
        POLYGON 182.645 189.240 188.765 187.890 182.645 187.890 ;
        POLYGON 222.370 189.240 222.370 187.890 216.255 187.890 ;
        RECT 222.370 187.890 277.645 189.240 ;
        POLYGON 277.645 189.240 283.765 187.890 277.645 187.890 ;
        POLYGON 121.255 187.890 121.255 186.305 115.315 186.305 ;
        RECT 121.255 186.305 188.765 187.890 ;
        POLYGON 188.765 187.890 194.705 186.305 188.765 186.305 ;
        POLYGON 216.255 187.890 216.255 186.305 210.315 186.305 ;
        RECT 216.255 186.305 283.765 187.890 ;
        POLYGON 283.765 187.890 289.705 186.305 283.765 186.305 ;
        POLYGON 115.315 186.305 115.315 184.485 109.510 184.485 ;
        RECT 115.315 184.485 194.705 186.305 ;
        POLYGON 194.705 186.305 200.505 184.485 194.705 184.485 ;
        POLYGON 210.315 186.305 210.315 184.485 204.510 184.485 ;
        RECT 210.315 184.485 289.705 186.305 ;
        POLYGON 289.705 186.305 295.505 184.485 289.705 184.485 ;
        POLYGON 109.510 184.485 109.510 182.410 103.815 182.410 ;
        RECT 109.510 183.755 200.505 184.485 ;
        POLYGON 200.505 184.485 202.505 183.755 200.505 183.755 ;
        POLYGON 204.510 184.485 204.510 183.755 202.510 183.755 ;
        RECT 204.510 183.755 295.505 184.485 ;
        RECT 109.510 182.410 295.505 183.755 ;
        POLYGON 295.505 184.485 301.205 182.410 295.505 182.410 ;
        POLYGON 103.815 182.410 103.815 180.080 98.180 180.080 ;
        RECT 103.815 181.620 301.205 182.410 ;
        POLYGON 301.205 182.410 303.120 181.620 301.205 181.620 ;
        RECT 103.815 180.080 303.120 181.620 ;
        POLYGON 98.180 180.080 98.180 177.475 92.570 177.475 ;
        RECT 98.180 177.475 303.120 180.080 ;
        POLYGON 92.570 177.475 92.570 173.390 84.855 173.390 ;
        RECT 92.570 173.390 303.120 177.475 ;
        POLYGON 84.855 173.390 84.855 168.870 77.450 168.870 ;
        RECT 84.855 168.870 303.120 173.390 ;
        POLYGON 77.450 168.870 77.450 163.925 70.370 163.925 ;
        RECT 77.450 163.925 303.120 168.870 ;
        POLYGON 70.370 163.925 70.370 158.575 63.630 158.575 ;
        RECT 70.370 158.575 303.120 163.925 ;
        POLYGON 63.630 158.575 63.630 152.845 57.250 152.845 ;
        RECT 63.630 152.845 303.120 158.575 ;
        POLYGON 57.250 152.845 57.250 146.750 51.235 146.750 ;
        RECT 57.250 146.750 303.120 152.845 ;
        POLYGON 51.235 146.750 51.235 140.310 45.605 140.310 ;
        RECT 51.235 140.310 303.120 146.750 ;
        POLYGON 45.605 140.310 45.605 133.550 40.375 133.550 ;
        RECT 45.605 133.550 303.120 140.310 ;
        POLYGON 40.375 133.550 40.375 126.490 35.560 126.490 ;
        RECT 40.375 126.490 303.120 133.550 ;
        POLYGON 35.560 126.490 35.560 119.145 31.170 119.145 ;
        RECT 35.560 119.145 303.120 126.490 ;
        POLYGON 31.170 119.145 31.170 111.535 27.225 111.535 ;
        RECT 31.170 111.535 303.120 119.145 ;
        POLYGON 27.225 111.535 27.225 103.685 23.730 103.685 ;
        RECT 27.225 103.685 303.120 111.535 ;
        POLYGON 23.730 103.685 23.730 95.610 20.715 95.610 ;
        RECT 23.730 95.610 303.120 103.685 ;
        POLYGON 20.715 95.610 20.715 87.330 18.180 87.330 ;
        RECT 20.715 87.330 303.120 95.610 ;
        POLYGON 18.180 87.330 18.180 78.870 16.145 78.870 ;
        RECT 18.180 78.870 303.120 87.330 ;
        POLYGON 16.145 78.870 16.145 70.245 14.625 70.245 ;
        RECT 16.145 70.245 303.120 78.870 ;
        POLYGON 14.625 70.245 14.625 65.420 14.030 65.420 ;
        RECT 14.625 65.420 303.120 70.245 ;
        POLYGON 14.030 65.420 14.030 60.390 13.610 60.390 ;
        RECT 14.030 60.390 303.120 65.420 ;
        POLYGON 13.610 60.390 13.610 55.230 13.355 55.230 ;
        RECT 13.610 55.230 303.120 60.390 ;
        POLYGON 13.355 55.230 13.355 50.000 13.270 50.000 ;
        RECT 13.355 50.000 303.120 55.230 ;
        RECT 5.000 40.000 303.120 50.000 ;
        POLYGON 13.590 40.000 13.610 40.000 13.610 39.610 ;
        RECT 13.610 39.610 303.120 40.000 ;
        POLYGON 13.610 39.610 14.030 39.610 14.030 34.580 ;
        RECT 14.030 34.580 303.120 39.610 ;
        POLYGON 14.030 34.580 14.625 34.580 14.625 29.755 ;
        RECT 14.625 29.755 303.120 34.580 ;
        POLYGON 14.625 29.755 16.145 29.755 16.145 21.130 ;
        RECT 16.145 21.130 303.120 29.755 ;
        POLYGON 16.145 21.130 18.180 21.130 18.180 12.670 ;
        RECT 18.180 12.670 303.120 21.130 ;
        POLYGON 18.180 12.670 20.715 12.670 20.715 4.390 ;
        RECT 20.715 4.390 303.120 12.670 ;
        POLYGON 20.715 4.390 22.355 4.390 22.355 0.000 ;
        RECT 22.355 0.000 303.120 4.390 ;
      LAYER met3 ;
        POLYGON 155.010 191.730 155.010 191.355 142.020 191.355 ;
        POLYGON 155.010 191.730 156.360 191.695 155.010 191.695 ;
        RECT 155.010 191.530 156.370 191.695 ;
        POLYGON 156.370 191.695 161.935 191.530 156.370 191.530 ;
        RECT 155.010 191.430 161.965 191.530 ;
        POLYGON 161.965 191.530 165.400 191.430 161.965 191.430 ;
        RECT 155.010 191.355 165.410 191.430 ;
        POLYGON 142.005 191.355 142.005 191.305 140.290 191.305 ;
        RECT 142.005 191.335 165.410 191.355 ;
        POLYGON 165.410 191.430 168.760 191.335 165.410 191.335 ;
        RECT 142.005 191.305 168.775 191.335 ;
        POLYGON 168.775 191.335 169.730 191.305 168.775 191.305 ;
        POLYGON 140.290 191.305 140.290 190.760 136.405 190.760 ;
        RECT 140.290 190.980 169.730 191.305 ;
        POLYGON 169.730 191.305 172.055 190.980 169.730 190.980 ;
        RECT 140.290 190.760 172.055 190.980 ;
        POLYGON 136.405 190.760 136.405 190.380 133.705 190.380 ;
        RECT 136.405 190.530 172.055 190.760 ;
        POLYGON 172.055 190.980 175.250 190.530 172.055 190.530 ;
        RECT 136.405 190.380 175.255 190.530 ;
        POLYGON 175.255 190.530 176.315 190.380 175.255 190.380 ;
        POLYGON 133.705 190.380 133.705 190.090 132.095 190.090 ;
        RECT 133.705 190.090 176.315 190.380 ;
        POLYGON 132.095 190.090 132.095 189.335 127.900 189.335 ;
        RECT 132.095 190.010 176.315 190.090 ;
        POLYGON 176.315 190.380 178.370 190.010 176.315 190.010 ;
        RECT 132.095 189.465 178.370 190.010 ;
        POLYGON 178.370 190.010 181.400 189.465 178.370 189.465 ;
        RECT 132.095 189.335 181.400 189.465 ;
        POLYGON 127.900 189.335 127.900 189.240 127.370 189.240 ;
        RECT 127.900 189.240 181.400 189.335 ;
        POLYGON 181.400 189.465 182.645 189.240 181.400 189.240 ;
        POLYGON 127.370 189.240 127.370 188.455 123.815 188.455 ;
        RECT 127.370 188.870 182.645 189.240 ;
        POLYGON 182.645 189.240 184.335 188.870 182.645 188.870 ;
        RECT 127.370 188.455 184.335 188.870 ;
        POLYGON 123.810 188.455 123.810 187.890 121.255 187.890 ;
        RECT 123.810 188.240 184.335 188.455 ;
        POLYGON 184.335 188.870 187.175 188.240 184.335 188.240 ;
        RECT 123.810 187.890 187.180 188.240 ;
        POLYGON 187.180 188.240 188.765 187.890 187.180 187.890 ;
        POLYGON 121.255 187.890 121.255 187.505 119.810 187.505 ;
        RECT 121.255 187.580 188.765 187.890 ;
        POLYGON 188.765 187.890 189.930 187.580 188.765 187.580 ;
        RECT 121.255 187.505 189.930 187.580 ;
        POLYGON 119.810 187.505 119.810 186.460 115.885 186.460 ;
        RECT 119.810 186.875 189.930 187.505 ;
        POLYGON 189.930 187.580 192.580 186.875 189.930 186.875 ;
        RECT 119.810 186.460 192.580 186.875 ;
        POLYGON 115.885 186.460 115.885 186.305 115.315 186.305 ;
        RECT 115.885 186.305 192.580 186.460 ;
        POLYGON 192.580 186.875 194.705 186.305 192.580 186.305 ;
        POLYGON 115.315 186.305 115.315 185.270 112.015 185.270 ;
        RECT 115.315 186.175 194.705 186.305 ;
        POLYGON 194.705 186.305 195.130 186.175 194.705 186.175 ;
        RECT 115.315 185.405 195.130 186.175 ;
        POLYGON 195.130 186.175 197.580 185.405 195.130 185.405 ;
        RECT 115.315 185.270 197.580 185.405 ;
        POLYGON 112.015 185.270 112.015 184.485 109.510 184.485 ;
        RECT 112.015 184.665 197.580 185.270 ;
        POLYGON 197.580 185.405 199.925 184.665 197.580 184.665 ;
        RECT 112.015 184.485 199.925 184.665 ;
        POLYGON 199.925 184.665 200.505 184.485 199.925 184.485 ;
        POLYGON 109.510 184.485 109.510 182.625 104.395 182.625 ;
        RECT 109.510 183.880 200.505 184.485 ;
        POLYGON 200.505 184.485 202.165 183.880 200.505 183.880 ;
        RECT 109.510 183.230 202.165 183.880 ;
        RECT 109.510 183.010 147.225 183.230 ;
        POLYGON 147.225 183.230 154.005 183.230 147.225 183.010 ;
        POLYGON 154.005 183.230 156.355 183.230 156.355 183.185 ;
        RECT 156.355 183.185 202.165 183.230 ;
        POLYGON 156.370 183.185 160.840 183.185 160.840 183.105 ;
        RECT 160.840 183.110 202.165 183.185 ;
        POLYGON 202.165 183.880 204.290 183.110 202.165 183.110 ;
        RECT 160.840 183.105 204.295 183.110 ;
        POLYGON 160.840 183.105 161.960 183.105 161.960 183.020 ;
        RECT 161.960 183.020 204.295 183.105 ;
        POLYGON 161.965 183.020 162.100 183.020 162.100 183.010 ;
        RECT 162.100 183.010 204.295 183.020 ;
        RECT 109.510 182.625 142.005 183.010 ;
        POLYGON 104.395 182.625 104.395 182.410 103.815 182.410 ;
        RECT 104.395 182.580 142.005 182.625 ;
        POLYGON 142.005 183.010 147.225 183.010 142.005 182.580 ;
        POLYGON 162.100 183.010 165.400 183.010 165.400 182.770 ;
        RECT 165.400 182.770 204.295 183.010 ;
        POLYGON 165.410 182.770 168.005 182.770 168.005 182.580 ;
        RECT 168.005 182.580 204.295 182.770 ;
        RECT 104.395 182.455 140.500 182.580 ;
        POLYGON 140.500 182.580 142.000 182.580 140.500 182.455 ;
        POLYGON 168.005 182.580 168.760 182.580 168.760 182.525 ;
        RECT 168.760 182.525 204.295 182.580 ;
        POLYGON 168.775 182.525 168.790 182.525 168.790 182.520 ;
        RECT 168.790 182.520 204.295 182.525 ;
        POLYGON 168.790 182.520 169.275 182.520 169.275 182.455 ;
        RECT 169.275 182.455 204.295 182.520 ;
        RECT 104.395 182.425 140.290 182.455 ;
        POLYGON 140.290 182.455 140.500 182.455 140.290 182.425 ;
        POLYGON 169.275 182.455 169.500 182.455 169.500 182.425 ;
        RECT 169.500 182.425 204.295 182.455 ;
        RECT 104.395 182.410 136.405 182.425 ;
        POLYGON 103.815 182.410 103.815 180.935 100.250 180.935 ;
        RECT 103.815 181.905 136.405 182.410 ;
        POLYGON 136.405 182.425 140.290 182.425 136.405 181.905 ;
        POLYGON 169.500 182.425 169.725 182.425 169.725 182.395 ;
        RECT 169.725 182.410 204.295 182.425 ;
        POLYGON 204.295 183.110 206.205 182.410 204.295 182.410 ;
        POLYGON 250.935 183.080 250.935 183.025 246.055 183.025 ;
        POLYGON 246.055 183.025 246.055 182.790 241.205 182.790 ;
        RECT 246.055 182.960 250.935 183.025 ;
        POLYGON 250.935 183.080 255.845 182.960 250.935 182.960 ;
        RECT 246.055 182.790 255.845 182.960 ;
        POLYGON 241.205 182.790 241.205 182.410 236.685 182.410 ;
        RECT 241.205 182.410 255.845 182.790 ;
        RECT 169.725 182.395 206.205 182.410 ;
        POLYGON 169.730 182.395 172.050 182.395 172.050 182.085 ;
        RECT 172.050 182.370 206.205 182.395 ;
        POLYGON 206.205 182.410 206.310 182.370 206.205 182.370 ;
        POLYGON 236.685 182.410 236.685 182.385 236.385 182.385 ;
        RECT 236.685 182.385 255.845 182.410 ;
        POLYGON 236.385 182.385 236.385 182.370 236.260 182.370 ;
        RECT 236.385 182.375 255.845 182.385 ;
        POLYGON 255.845 182.960 263.785 182.375 255.845 182.375 ;
        RECT 236.385 182.370 263.785 182.375 ;
        RECT 172.050 182.085 206.310 182.370 ;
        POLYGON 172.055 182.085 173.410 182.085 173.410 181.905 ;
        RECT 173.410 181.905 206.310 182.085 ;
        RECT 103.815 181.565 133.840 181.905 ;
        POLYGON 133.840 181.905 136.405 181.905 133.840 181.565 ;
        POLYGON 173.410 181.905 175.255 181.905 175.255 181.660 ;
        RECT 175.255 181.660 206.310 181.905 ;
        POLYGON 175.255 181.660 175.945 181.660 175.945 181.565 ;
        RECT 175.945 181.645 206.310 181.660 ;
        POLYGON 206.310 182.370 208.060 181.645 206.310 181.645 ;
        POLYGON 236.260 182.370 236.260 181.805 231.605 181.805 ;
        RECT 236.260 181.805 263.785 182.370 ;
        POLYGON 231.605 181.805 231.605 181.645 230.595 181.645 ;
        RECT 231.605 181.645 263.785 181.805 ;
        RECT 175.945 181.565 208.060 181.645 ;
        RECT 103.815 181.540 133.705 181.565 ;
        POLYGON 133.705 181.565 133.840 181.565 133.705 181.540 ;
        POLYGON 175.945 181.565 176.125 181.565 176.125 181.540 ;
        RECT 176.125 181.540 208.060 181.565 ;
        RECT 103.815 181.240 132.095 181.540 ;
        POLYGON 132.095 181.540 133.705 181.540 132.095 181.240 ;
        POLYGON 176.125 181.540 176.310 181.540 176.310 181.515 ;
        RECT 176.310 181.515 208.060 181.540 ;
        POLYGON 176.315 181.515 176.640 181.515 176.640 181.475 ;
        RECT 176.640 181.475 208.060 181.515 ;
        POLYGON 176.640 181.475 177.835 181.475 177.835 181.240 ;
        RECT 177.835 181.240 208.060 181.475 ;
        RECT 103.815 180.935 127.900 181.240 ;
        POLYGON 100.250 180.935 100.250 180.080 98.180 180.080 ;
        RECT 100.250 180.460 127.900 180.935 ;
        POLYGON 127.900 181.240 132.095 181.240 127.900 180.460 ;
        POLYGON 177.835 181.240 178.370 181.240 178.370 181.135 ;
        RECT 178.370 181.135 208.060 181.240 ;
        POLYGON 178.370 181.135 181.395 181.135 181.395 180.545 ;
        RECT 181.395 181.020 208.060 181.135 ;
        POLYGON 208.060 181.645 209.570 181.020 208.060 181.020 ;
        POLYGON 230.595 181.645 230.595 181.055 226.865 181.055 ;
        RECT 230.595 181.330 263.785 181.645 ;
        POLYGON 263.785 182.375 271.630 181.330 263.785 181.330 ;
        RECT 230.595 181.055 271.630 181.330 ;
        POLYGON 226.865 181.055 226.865 181.020 226.685 181.020 ;
        RECT 226.865 181.020 271.630 181.055 ;
        RECT 181.395 180.545 209.570 181.020 ;
        POLYGON 181.400 180.545 181.840 180.545 181.840 180.460 ;
        RECT 181.840 180.485 209.570 180.545 ;
        POLYGON 209.570 181.020 210.860 180.485 209.570 180.485 ;
        POLYGON 226.685 181.020 226.685 180.485 223.940 180.485 ;
        RECT 226.685 180.485 271.630 181.020 ;
        RECT 181.840 180.460 210.865 180.485 ;
        RECT 100.250 180.365 127.375 180.460 ;
        POLYGON 127.375 180.460 127.900 180.460 127.375 180.365 ;
        POLYGON 181.840 180.460 182.330 180.460 182.330 180.365 ;
        RECT 182.330 180.365 210.865 180.460 ;
        RECT 100.250 180.340 127.260 180.365 ;
        POLYGON 127.260 180.365 127.370 180.365 127.260 180.340 ;
        POLYGON 182.330 180.365 182.460 180.365 182.460 180.340 ;
        RECT 182.460 180.340 210.865 180.365 ;
        RECT 100.250 180.080 123.810 180.340 ;
        POLYGON 98.180 180.080 98.180 179.160 96.205 179.160 ;
        RECT 98.180 179.520 123.810 180.080 ;
        POLYGON 123.810 180.340 127.260 180.340 123.810 179.520 ;
        POLYGON 182.460 180.340 182.645 180.340 182.645 180.305 ;
        RECT 182.645 180.305 210.865 180.340 ;
        POLYGON 182.645 180.305 184.335 180.305 184.335 179.975 ;
        RECT 184.335 180.080 210.865 180.305 ;
        POLYGON 210.865 180.485 211.840 180.080 210.865 180.080 ;
        POLYGON 223.940 180.485 223.940 180.140 222.170 180.140 ;
        RECT 223.940 180.140 271.630 180.485 ;
        POLYGON 222.170 180.140 222.170 180.080 221.915 180.080 ;
        RECT 222.170 180.080 271.630 180.140 ;
        RECT 184.335 180.020 211.840 180.080 ;
        POLYGON 211.840 180.080 211.965 180.020 211.840 180.020 ;
        POLYGON 221.915 180.080 221.915 180.020 221.655 180.020 ;
        RECT 221.915 180.020 271.630 180.080 ;
        RECT 184.335 179.975 211.970 180.020 ;
        POLYGON 184.335 179.975 184.370 179.975 184.370 179.970 ;
        RECT 184.370 179.970 211.970 179.975 ;
        POLYGON 184.370 179.970 186.110 179.970 186.110 179.520 ;
        RECT 186.110 179.790 211.970 179.970 ;
        POLYGON 211.970 180.020 212.460 179.790 211.970 179.790 ;
        POLYGON 221.655 180.020 221.655 179.790 220.670 179.790 ;
        RECT 221.655 179.825 271.630 180.020 ;
        POLYGON 271.630 181.330 279.355 179.825 271.630 179.825 ;
        RECT 221.655 179.790 279.355 179.825 ;
        RECT 186.110 179.580 212.460 179.790 ;
        POLYGON 212.460 179.790 212.915 179.580 212.460 179.580 ;
        POLYGON 220.670 179.790 220.670 179.580 219.775 179.580 ;
        RECT 220.670 179.580 279.355 179.790 ;
        RECT 186.110 179.520 212.915 179.580 ;
        RECT 98.180 179.160 121.255 179.520 ;
        POLYGON 96.205 179.160 96.205 177.475 92.570 177.475 ;
        RECT 96.205 178.910 121.255 179.160 ;
        POLYGON 121.255 179.520 123.810 179.520 121.255 178.910 ;
        POLYGON 186.110 179.520 187.180 179.520 187.180 179.245 ;
        RECT 187.180 179.385 212.915 179.520 ;
        POLYGON 212.915 179.580 213.335 179.385 212.915 179.385 ;
        POLYGON 219.775 179.580 219.775 179.385 218.940 179.385 ;
        RECT 219.775 179.385 279.355 179.580 ;
        RECT 187.180 179.245 213.335 179.385 ;
        POLYGON 187.180 179.245 188.490 179.245 188.490 178.910 ;
        RECT 188.490 179.200 213.335 179.245 ;
        POLYGON 213.335 179.385 213.725 179.200 213.335 179.200 ;
        POLYGON 218.940 179.385 218.940 179.200 218.145 179.200 ;
        RECT 218.940 179.200 279.355 179.385 ;
        RECT 188.490 179.055 213.730 179.200 ;
        POLYGON 213.730 179.200 214.040 179.055 213.730 179.055 ;
        POLYGON 218.145 179.200 218.145 179.055 217.525 179.055 ;
        RECT 218.145 179.055 279.355 179.200 ;
        RECT 188.490 178.910 214.040 179.055 ;
        RECT 96.205 178.795 120.770 178.910 ;
        POLYGON 120.770 178.910 121.255 178.910 120.770 178.795 ;
        POLYGON 188.490 178.910 188.765 178.910 188.765 178.840 ;
        RECT 188.765 178.870 214.040 178.910 ;
        POLYGON 214.040 179.055 214.435 178.870 214.040 178.870 ;
        POLYGON 217.525 179.055 217.525 178.870 216.840 178.870 ;
        RECT 217.525 178.870 279.355 179.055 ;
        RECT 188.765 178.840 214.440 178.870 ;
        POLYGON 188.765 178.840 188.935 178.840 188.935 178.795 ;
        RECT 188.935 178.795 214.440 178.840 ;
        RECT 96.205 178.515 119.810 178.795 ;
        POLYGON 119.810 178.795 120.770 178.795 119.810 178.515 ;
        POLYGON 188.935 178.795 189.925 178.795 189.925 178.540 ;
        RECT 189.925 178.575 214.440 178.795 ;
        POLYGON 214.440 178.870 215.070 178.575 214.440 178.575 ;
        POLYGON 216.840 178.870 216.840 178.575 215.755 178.575 ;
        RECT 216.840 178.575 279.355 178.870 ;
        RECT 189.925 178.540 215.070 178.575 ;
        POLYGON 189.930 178.540 190.025 178.540 190.025 178.515 ;
        RECT 190.025 178.515 215.070 178.540 ;
        RECT 96.205 177.475 115.885 178.515 ;
        POLYGON 92.570 177.475 92.570 177.315 92.270 177.315 ;
        RECT 92.570 177.365 115.885 177.475 ;
        POLYGON 115.885 178.515 119.810 178.515 115.885 177.365 ;
        POLYGON 190.025 178.515 191.965 178.515 191.965 178.015 ;
        RECT 191.965 178.505 215.070 178.515 ;
        POLYGON 215.070 178.575 215.225 178.505 215.070 178.505 ;
        POLYGON 215.755 178.575 215.755 178.505 215.495 178.505 ;
        RECT 215.755 178.505 279.355 178.575 ;
        RECT 191.965 178.465 215.225 178.505 ;
        POLYGON 215.225 178.505 215.310 178.465 215.225 178.465 ;
        POLYGON 215.495 178.505 215.495 178.465 215.345 178.465 ;
        RECT 215.495 178.465 279.355 178.505 ;
        RECT 191.965 178.460 215.310 178.465 ;
        POLYGON 215.310 178.465 215.320 178.460 215.310 178.460 ;
        POLYGON 215.345 178.465 215.345 178.460 215.335 178.460 ;
        RECT 215.345 178.460 279.355 178.465 ;
        RECT 191.965 178.015 279.355 178.460 ;
        POLYGON 191.965 178.015 192.580 178.015 192.580 177.820 ;
        RECT 192.580 177.875 279.355 178.015 ;
        POLYGON 279.355 179.825 286.945 177.875 279.355 177.875 ;
        RECT 192.580 177.820 286.945 177.875 ;
        POLYGON 192.580 177.820 194.000 177.820 194.000 177.365 ;
        RECT 194.000 177.365 286.945 177.820 ;
        RECT 92.570 177.315 115.315 177.365 ;
        POLYGON 92.270 177.315 92.270 175.295 88.450 175.295 ;
        RECT 92.270 177.195 115.315 177.315 ;
        POLYGON 115.315 177.365 115.885 177.365 115.315 177.195 ;
        POLYGON 194.000 177.365 194.530 177.365 194.530 177.195 ;
        RECT 194.530 177.195 286.945 177.365 ;
        RECT 92.270 176.920 114.370 177.195 ;
        POLYGON 114.370 177.195 115.315 177.195 114.370 176.920 ;
        POLYGON 194.530 177.195 194.705 177.195 194.705 177.140 ;
        RECT 194.705 177.140 286.945 177.195 ;
        POLYGON 194.705 177.140 195.130 177.140 195.130 177.005 ;
        RECT 195.130 177.005 286.945 177.140 ;
        POLYGON 195.130 177.005 195.390 177.005 195.390 176.920 ;
        RECT 195.390 176.920 286.945 177.005 ;
        RECT 92.270 176.100 112.015 176.920 ;
        POLYGON 112.015 176.920 114.370 176.920 112.015 176.100 ;
        POLYGON 195.390 176.920 197.580 176.920 197.580 176.215 ;
        RECT 197.580 176.215 286.945 176.920 ;
        POLYGON 197.580 176.215 197.935 176.215 197.935 176.100 ;
        RECT 197.935 176.100 286.945 176.215 ;
        RECT 92.270 175.295 109.510 176.100 ;
        POLYGON 88.450 175.295 88.450 173.390 84.855 173.390 ;
        RECT 88.450 175.225 109.510 175.295 ;
        POLYGON 109.510 176.100 112.015 176.100 109.510 175.225 ;
        POLYGON 197.935 176.100 199.410 176.100 199.410 175.630 ;
        RECT 199.410 175.630 286.945 176.100 ;
        POLYGON 199.410 175.630 199.925 175.630 199.925 175.430 ;
        RECT 199.925 175.495 286.945 175.630 ;
        POLYGON 286.945 177.875 294.380 175.495 286.945 175.495 ;
        RECT 199.925 175.430 294.380 175.495 ;
        POLYGON 199.925 175.430 200.450 175.430 200.450 175.225 ;
        RECT 200.450 175.225 294.380 175.430 ;
        RECT 88.450 174.765 108.190 175.225 ;
        POLYGON 108.190 175.225 109.510 175.225 108.190 174.765 ;
        POLYGON 200.450 175.225 200.505 175.225 200.505 175.205 ;
        RECT 200.505 175.205 294.380 175.225 ;
        POLYGON 200.505 175.205 201.440 175.205 201.440 174.845 ;
        RECT 201.440 174.845 294.380 175.205 ;
        POLYGON 201.440 174.845 201.645 174.845 201.645 174.765 ;
        RECT 201.645 174.765 294.380 174.845 ;
        RECT 88.450 174.725 108.080 174.765 ;
        POLYGON 108.080 174.765 108.190 174.765 108.080 174.725 ;
        POLYGON 201.645 174.765 201.750 174.765 201.750 174.725 ;
        RECT 201.750 174.725 294.380 174.765 ;
        RECT 88.450 173.390 104.395 174.725 ;
        POLYGON 84.855 173.390 84.855 173.335 84.765 173.335 ;
        RECT 84.855 173.335 104.395 173.390 ;
        POLYGON 84.765 173.335 84.765 171.170 81.220 171.170 ;
        RECT 84.765 173.225 104.395 173.335 ;
        POLYGON 104.395 174.725 108.080 174.725 104.395 173.225 ;
        POLYGON 201.750 174.725 202.165 174.725 202.165 174.565 ;
        RECT 202.165 174.565 294.380 174.725 ;
        POLYGON 202.165 174.565 202.765 174.565 202.765 174.365 ;
        POLYGON 202.765 174.360 202.765 174.160 202.165 174.160 ;
        RECT 202.765 174.160 294.380 174.565 ;
        POLYGON 202.165 174.160 202.165 173.885 201.460 173.885 ;
        RECT 202.165 173.885 294.380 174.160 ;
        POLYGON 201.460 173.885 201.460 173.740 201.085 173.740 ;
        RECT 201.460 173.740 294.380 173.885 ;
        POLYGON 201.085 173.740 201.085 173.225 199.765 173.225 ;
        RECT 201.085 173.225 294.380 173.740 ;
        RECT 84.765 172.990 103.815 173.225 ;
        POLYGON 103.815 173.225 104.390 173.225 103.815 172.990 ;
        POLYGON 199.765 173.225 199.765 173.125 199.510 173.125 ;
        RECT 199.765 173.125 294.380 173.225 ;
        POLYGON 199.510 173.125 199.510 172.990 199.195 172.990 ;
        RECT 199.510 172.990 294.380 173.125 ;
        RECT 84.765 172.215 101.910 172.990 ;
        POLYGON 101.910 172.990 103.815 172.990 101.910 172.215 ;
        POLYGON 199.195 172.990 199.195 172.960 199.125 172.960 ;
        RECT 199.195 172.960 294.380 172.990 ;
        POLYGON 199.125 172.960 199.125 172.820 198.800 172.820 ;
        RECT 199.125 172.820 294.380 172.960 ;
        POLYGON 198.800 172.820 198.800 172.215 197.400 172.215 ;
        RECT 198.800 172.685 294.380 172.820 ;
        POLYGON 294.380 175.495 301.645 172.685 294.380 172.685 ;
        RECT 198.800 172.215 301.645 172.685 ;
        RECT 84.765 171.445 100.250 172.215 ;
        POLYGON 100.250 172.215 101.910 172.215 100.250 171.445 ;
        POLYGON 197.400 172.215 197.400 172.190 197.340 172.190 ;
        RECT 197.400 172.190 301.645 172.215 ;
        POLYGON 197.340 172.190 197.340 171.505 195.750 171.505 ;
        RECT 197.340 172.015 301.645 172.190 ;
        POLYGON 301.645 172.685 303.120 172.015 301.645 172.015 ;
        RECT 197.340 171.505 303.120 172.015 ;
        POLYGON 195.750 171.505 195.750 171.445 195.610 171.445 ;
        RECT 195.750 171.445 303.120 171.505 ;
        RECT 84.765 171.170 98.180 171.445 ;
        POLYGON 81.220 171.170 81.220 169.100 77.825 169.100 ;
        RECT 81.220 170.475 98.180 171.170 ;
        POLYGON 98.180 171.445 100.250 171.445 98.180 170.475 ;
        POLYGON 195.610 171.445 195.610 171.255 195.170 171.255 ;
        RECT 195.610 171.255 303.120 171.445 ;
        POLYGON 195.170 171.255 195.170 170.915 194.455 170.915 ;
        RECT 195.170 170.915 303.120 171.255 ;
        POLYGON 194.455 170.915 194.455 170.475 193.525 170.475 ;
        RECT 194.455 170.475 303.120 170.915 ;
        RECT 81.220 169.555 96.205 170.475 ;
        POLYGON 96.205 170.475 98.180 170.475 96.205 169.555 ;
        POLYGON 193.525 170.475 193.525 170.470 193.515 170.470 ;
        RECT 193.525 170.470 303.120 170.475 ;
        POLYGON 193.515 170.470 193.515 170.410 193.390 170.410 ;
        RECT 193.515 170.410 303.120 170.470 ;
        POLYGON 193.390 170.410 193.390 170.350 193.260 170.350 ;
        RECT 193.390 170.350 303.120 170.410 ;
        POLYGON 149.190 170.350 149.190 170.310 147.245 170.310 ;
        POLYGON 147.225 170.310 147.225 170.205 142.005 170.205 ;
        RECT 147.225 170.250 149.190 170.310 ;
        POLYGON 149.190 170.350 153.980 170.250 149.190 170.250 ;
        POLYGON 193.260 170.350 193.260 170.250 193.050 170.250 ;
        RECT 193.260 170.250 303.120 170.350 ;
        RECT 147.225 170.205 154.005 170.250 ;
        POLYGON 142.000 170.205 142.000 170.085 140.500 170.085 ;
        RECT 142.000 170.200 154.005 170.205 ;
        POLYGON 154.005 170.250 156.370 170.200 154.005 170.200 ;
        POLYGON 193.050 170.250 193.050 170.200 192.945 170.200 ;
        RECT 193.050 170.220 303.120 170.250 ;
        RECT 193.050 170.200 241.225 170.220 ;
        RECT 142.000 170.085 156.370 170.200 ;
        POLYGON 140.500 170.085 140.500 170.065 140.290 170.065 ;
        RECT 140.500 170.065 156.370 170.085 ;
        POLYGON 140.290 170.065 140.290 169.755 136.405 169.755 ;
        RECT 140.290 169.835 156.370 170.065 ;
        POLYGON 156.370 170.200 160.830 169.835 156.370 169.835 ;
        POLYGON 192.945 170.200 192.945 170.185 192.915 170.185 ;
        RECT 192.945 170.185 241.225 170.200 ;
        POLYGON 192.915 170.185 192.915 169.980 192.480 169.980 ;
        RECT 192.915 170.160 241.225 170.185 ;
        POLYGON 241.225 170.220 244.205 170.220 241.225 170.160 ;
        POLYGON 244.205 170.220 246.035 170.220 246.035 170.180 ;
        RECT 246.035 170.180 303.120 170.220 ;
        POLYGON 246.055 170.180 246.975 170.180 246.975 170.160 ;
        RECT 246.975 170.160 303.120 170.180 ;
        RECT 192.915 170.075 237.025 170.160 ;
        POLYGON 237.025 170.160 241.205 170.160 237.025 170.075 ;
        POLYGON 246.975 170.160 250.910 170.160 250.910 170.075 ;
        RECT 250.910 170.075 303.120 170.160 ;
        RECT 192.915 170.020 236.390 170.075 ;
        POLYGON 236.390 170.075 237.025 170.075 236.390 170.020 ;
        POLYGON 250.935 170.075 251.380 170.075 251.380 170.065 ;
        RECT 251.380 170.065 303.120 170.075 ;
        POLYGON 251.380 170.065 251.935 170.065 251.935 170.020 ;
        RECT 251.935 170.020 303.120 170.065 ;
        RECT 192.915 169.980 231.610 170.020 ;
        POLYGON 192.480 169.980 192.480 169.835 192.175 169.835 ;
        RECT 192.480 169.835 231.610 169.980 ;
        RECT 140.290 169.755 160.840 169.835 ;
        POLYGON 136.405 169.755 136.405 169.555 135.140 169.555 ;
        RECT 136.405 169.745 160.840 169.755 ;
        POLYGON 160.840 169.835 161.965 169.745 160.840 169.745 ;
        POLYGON 192.175 169.835 192.175 169.785 192.070 169.785 ;
        RECT 192.175 169.785 231.610 169.835 ;
        POLYGON 192.070 169.785 192.070 169.745 191.985 169.745 ;
        RECT 192.070 169.745 231.610 169.785 ;
        RECT 136.405 169.555 161.965 169.745 ;
        RECT 81.220 169.395 95.860 169.555 ;
        POLYGON 95.860 169.555 96.205 169.555 95.860 169.395 ;
        POLYGON 135.140 169.555 135.140 169.395 134.130 169.395 ;
        RECT 135.140 169.395 161.965 169.555 ;
        RECT 81.220 169.100 92.570 169.395 ;
        POLYGON 77.825 169.100 77.825 168.870 77.450 168.870 ;
        RECT 77.825 168.870 92.570 169.100 ;
        POLYGON 77.450 168.870 77.450 166.875 74.595 166.875 ;
        RECT 77.450 167.650 92.570 168.870 ;
        POLYGON 92.570 169.395 95.860 169.395 92.570 167.650 ;
        POLYGON 134.130 169.395 134.130 169.350 133.845 169.350 ;
        RECT 134.130 169.350 161.965 169.395 ;
        POLYGON 133.840 169.350 133.840 169.325 133.705 169.325 ;
        RECT 133.840 169.325 161.965 169.350 ;
        POLYGON 133.705 169.325 133.705 169.075 132.095 169.075 ;
        RECT 133.705 169.205 161.965 169.325 ;
        POLYGON 161.965 169.745 165.410 169.205 161.965 169.205 ;
        POLYGON 191.985 169.745 191.985 169.610 191.700 169.610 ;
        RECT 191.985 169.640 231.610 169.745 ;
        POLYGON 231.610 170.020 236.385 170.020 231.610 169.640 ;
        POLYGON 251.935 170.020 255.835 170.020 255.835 169.705 ;
        RECT 255.835 169.705 303.120 170.020 ;
        POLYGON 255.845 169.705 256.655 169.705 256.655 169.640 ;
        RECT 256.655 169.640 303.120 169.705 ;
        RECT 191.985 169.625 231.435 169.640 ;
        POLYGON 231.435 169.640 231.605 169.640 231.435 169.625 ;
        POLYGON 256.655 169.640 256.845 169.640 256.845 169.625 ;
        RECT 256.845 169.625 303.120 169.640 ;
        RECT 191.985 169.620 231.405 169.625 ;
        POLYGON 231.405 169.625 231.435 169.625 231.405 169.620 ;
        POLYGON 256.845 169.625 256.905 169.625 256.905 169.620 ;
        RECT 256.905 169.620 303.120 169.625 ;
        RECT 191.985 169.615 231.370 169.620 ;
        POLYGON 231.370 169.620 231.405 169.620 231.370 169.615 ;
        POLYGON 256.905 169.620 256.970 169.620 256.970 169.615 ;
        RECT 256.970 169.615 303.120 169.620 ;
        RECT 191.985 169.610 231.350 169.615 ;
        POLYGON 231.350 169.615 231.360 169.610 231.350 169.610 ;
        POLYGON 256.970 169.615 257.000 169.615 257.000 169.610 ;
        RECT 257.000 169.610 303.120 169.615 ;
        POLYGON 191.700 169.610 191.700 169.590 191.660 169.590 ;
        RECT 191.700 169.590 231.360 169.610 ;
        POLYGON 191.660 169.590 191.660 169.235 190.910 169.235 ;
        RECT 191.660 169.565 231.360 169.590 ;
        POLYGON 231.360 169.610 231.435 169.565 231.360 169.565 ;
        POLYGON 257.000 169.610 257.285 169.610 257.285 169.565 ;
        RECT 257.285 169.565 303.120 169.610 ;
        RECT 191.660 169.235 231.435 169.565 ;
        POLYGON 190.910 169.235 190.910 169.205 190.850 169.205 ;
        RECT 190.910 169.205 231.435 169.235 ;
        RECT 133.705 169.075 165.410 169.205 ;
        POLYGON 132.095 169.075 132.095 168.255 127.900 168.255 ;
        RECT 132.095 168.560 165.410 169.075 ;
        POLYGON 165.410 169.205 168.775 168.560 165.410 168.560 ;
        POLYGON 190.850 169.205 190.850 168.900 190.265 168.900 ;
        RECT 190.850 168.945 231.435 169.205 ;
        POLYGON 231.435 169.565 232.450 168.945 231.435 168.945 ;
        POLYGON 257.285 169.565 260.410 169.565 260.410 169.075 ;
        RECT 260.410 169.075 303.120 169.565 ;
        POLYGON 260.410 169.075 261.090 169.075 261.090 168.945 ;
        RECT 261.090 168.945 303.120 169.075 ;
        RECT 190.850 168.900 232.450 168.945 ;
        POLYGON 190.265 168.900 190.265 168.820 190.110 168.820 ;
        RECT 190.265 168.895 232.450 168.900 ;
        POLYGON 232.450 168.945 232.530 168.895 232.450 168.895 ;
        POLYGON 261.090 168.945 261.355 168.945 261.355 168.895 ;
        RECT 261.355 168.895 303.120 168.945 ;
        RECT 190.265 168.870 232.530 168.895 ;
        POLYGON 232.530 168.895 232.570 168.870 232.530 168.870 ;
        POLYGON 261.355 168.895 261.485 168.895 261.485 168.870 ;
        RECT 261.485 168.870 303.120 168.895 ;
        RECT 190.265 168.820 232.570 168.870 ;
        POLYGON 190.110 168.820 190.110 168.755 189.985 168.755 ;
        RECT 190.110 168.755 232.570 168.820 ;
        POLYGON 189.985 168.755 189.985 168.705 189.885 168.705 ;
        RECT 189.985 168.705 232.570 168.755 ;
        POLYGON 189.885 168.705 189.885 168.665 189.810 168.665 ;
        RECT 189.885 168.665 232.570 168.705 ;
        POLYGON 189.810 168.665 189.810 168.630 189.740 168.630 ;
        RECT 189.810 168.630 232.570 168.665 ;
        POLYGON 189.740 168.630 189.740 168.560 189.605 168.560 ;
        RECT 189.740 168.560 232.570 168.630 ;
        RECT 132.095 168.345 168.790 168.560 ;
        POLYGON 168.790 168.560 169.730 168.345 168.790 168.345 ;
        POLYGON 189.605 168.560 189.605 168.345 189.190 168.345 ;
        RECT 189.605 168.345 232.570 168.560 ;
        RECT 132.095 168.255 169.730 168.345 ;
        POLYGON 127.900 168.255 127.900 168.130 127.370 168.130 ;
        RECT 127.900 168.130 169.730 168.255 ;
        POLYGON 127.370 168.130 127.370 168.105 127.260 168.105 ;
        RECT 127.370 168.105 169.730 168.130 ;
        POLYGON 127.260 168.105 127.260 167.650 125.310 167.650 ;
        RECT 127.260 167.825 169.730 168.105 ;
        POLYGON 169.730 168.345 172.055 167.825 169.730 167.825 ;
        POLYGON 189.190 168.345 189.190 167.825 188.185 167.825 ;
        RECT 189.190 167.825 232.570 168.345 ;
        RECT 127.260 167.650 172.055 167.825 ;
        RECT 77.450 167.490 92.270 167.650 ;
        POLYGON 92.270 167.650 92.570 167.650 92.270 167.490 ;
        POLYGON 125.310 167.650 125.310 167.490 124.625 167.490 ;
        RECT 125.310 167.490 172.055 167.650 ;
        RECT 77.450 166.875 89.950 167.490 ;
        POLYGON 74.595 166.875 74.595 164.630 71.385 164.630 ;
        RECT 74.595 166.260 89.950 166.875 ;
        POLYGON 89.950 167.490 92.270 167.490 89.950 166.260 ;
        POLYGON 124.625 167.490 124.625 167.300 123.810 167.300 ;
        RECT 124.625 167.300 172.055 167.490 ;
        POLYGON 123.810 167.300 123.810 166.595 121.255 166.595 ;
        RECT 123.810 166.990 172.055 167.300 ;
        POLYGON 172.055 167.825 175.255 166.990 172.055 166.990 ;
        POLYGON 188.185 167.825 188.185 167.645 187.840 167.645 ;
        RECT 188.185 167.645 232.570 167.825 ;
        POLYGON 187.840 167.645 187.840 167.060 186.710 167.060 ;
        RECT 187.840 167.075 232.570 167.645 ;
        RECT 187.840 167.065 218.470 167.075 ;
        POLYGON 218.470 167.075 218.505 167.075 218.470 167.065 ;
        POLYGON 218.520 167.075 218.540 167.075 218.540 167.065 ;
        RECT 218.540 167.065 232.570 167.075 ;
        RECT 187.840 167.060 218.345 167.065 ;
        POLYGON 186.710 167.060 186.710 166.990 186.585 166.990 ;
        RECT 186.710 167.030 218.345 167.060 ;
        POLYGON 218.345 167.065 218.470 167.065 218.345 167.030 ;
        POLYGON 218.545 167.065 218.610 167.065 218.610 167.030 ;
        RECT 218.610 167.030 232.570 167.065 ;
        RECT 186.710 166.990 217.890 167.030 ;
        RECT 123.810 166.675 175.255 166.990 ;
        POLYGON 175.255 166.990 176.310 166.675 175.255 166.675 ;
        POLYGON 186.585 166.990 186.585 166.675 186.025 166.675 ;
        RECT 186.585 166.905 217.890 166.990 ;
        POLYGON 217.890 167.030 218.340 167.030 217.890 166.905 ;
        POLYGON 218.610 167.030 218.850 167.030 218.850 166.905 ;
        RECT 218.850 166.905 232.570 167.030 ;
        RECT 186.585 166.805 217.525 166.905 ;
        POLYGON 217.525 166.905 217.890 166.905 217.525 166.805 ;
        POLYGON 218.850 166.905 219.035 166.905 219.035 166.805 ;
        RECT 219.035 166.805 232.570 166.905 ;
        RECT 186.585 166.675 217.050 166.805 ;
        POLYGON 217.050 166.805 217.525 166.805 217.050 166.675 ;
        POLYGON 219.035 166.805 219.280 166.805 219.280 166.675 ;
        RECT 219.280 166.675 232.570 166.805 ;
        RECT 123.810 166.595 176.315 166.675 ;
        POLYGON 121.255 166.595 121.255 166.460 120.770 166.460 ;
        RECT 121.255 166.575 176.315 166.595 ;
        POLYGON 176.315 166.675 176.640 166.575 176.315 166.575 ;
        POLYGON 186.025 166.675 186.025 166.575 185.850 166.575 ;
        RECT 186.025 166.575 216.690 166.675 ;
        POLYGON 216.690 166.675 217.050 166.675 216.690 166.575 ;
        POLYGON 219.280 166.675 219.470 166.675 219.470 166.575 ;
        RECT 219.470 166.575 232.570 166.675 ;
        RECT 121.255 166.460 176.640 166.575 ;
        POLYGON 120.770 166.460 120.770 166.260 120.030 166.260 ;
        RECT 120.770 166.260 176.640 166.460 ;
        RECT 74.595 165.370 88.455 166.260 ;
        POLYGON 88.455 166.260 89.950 166.260 88.455 165.370 ;
        POLYGON 120.030 166.260 120.030 166.200 119.810 166.200 ;
        RECT 120.030 166.200 176.640 166.260 ;
        POLYGON 119.810 166.200 119.810 165.370 117.215 165.370 ;
        RECT 119.810 166.055 176.640 166.200 ;
        POLYGON 176.640 166.575 178.370 166.055 176.640 166.055 ;
        POLYGON 185.850 166.575 185.850 166.055 184.925 166.055 ;
        RECT 185.850 166.070 214.850 166.575 ;
        POLYGON 214.850 166.575 216.690 166.575 214.850 166.070 ;
        POLYGON 219.470 166.575 220.425 166.575 220.425 166.070 ;
        RECT 220.425 166.070 232.570 166.575 ;
        RECT 185.850 166.055 214.805 166.070 ;
        POLYGON 214.805 166.070 214.850 166.070 214.805 166.055 ;
        POLYGON 220.425 166.070 220.455 166.070 220.455 166.055 ;
        RECT 220.455 166.055 232.570 166.070 ;
        RECT 119.810 165.370 178.370 166.055 ;
        RECT 74.595 164.630 84.855 165.370 ;
        POLYGON 71.385 164.630 71.385 163.925 70.370 163.925 ;
        RECT 71.385 163.925 84.855 164.630 ;
        POLYGON 70.370 163.925 70.370 162.570 68.665 162.570 ;
        RECT 70.370 163.230 84.855 163.925 ;
        POLYGON 84.855 165.370 88.450 165.370 84.855 163.230 ;
        POLYGON 117.215 165.370 117.215 164.945 115.885 164.945 ;
        RECT 117.215 165.030 178.370 165.370 ;
        POLYGON 178.370 166.055 181.400 165.030 178.370 165.030 ;
        POLYGON 184.925 166.055 184.925 165.960 184.755 165.960 ;
        RECT 184.925 165.960 214.505 166.055 ;
        POLYGON 214.505 166.055 214.805 166.055 214.505 165.960 ;
        POLYGON 220.455 166.055 220.635 166.055 220.635 165.960 ;
        RECT 220.635 165.960 232.570 166.055 ;
        POLYGON 184.755 165.960 184.755 165.030 183.105 165.030 ;
        RECT 184.755 165.460 212.930 165.960 ;
        POLYGON 212.930 165.960 214.505 165.960 212.930 165.460 ;
        POLYGON 220.635 165.960 221.455 165.960 221.455 165.460 ;
        RECT 221.455 165.460 232.570 165.960 ;
        RECT 184.755 165.030 211.575 165.460 ;
        POLYGON 211.575 165.460 212.930 165.460 211.575 165.030 ;
        POLYGON 221.455 165.460 222.165 165.460 222.165 165.030 ;
        RECT 222.165 165.030 232.570 165.460 ;
        RECT 117.215 164.945 181.400 165.030 ;
        POLYGON 115.885 164.945 115.885 164.740 115.315 164.740 ;
        RECT 115.885 164.745 181.400 164.945 ;
        POLYGON 181.400 165.030 182.145 164.745 181.400 164.745 ;
        POLYGON 183.105 165.030 183.105 164.745 182.600 164.745 ;
        RECT 183.105 164.825 210.930 165.030 ;
        POLYGON 210.930 165.030 211.575 165.030 210.930 164.825 ;
        POLYGON 222.165 165.030 222.500 165.030 222.500 164.825 ;
        RECT 222.500 164.825 232.570 165.030 ;
        RECT 183.105 164.745 210.185 164.825 ;
        RECT 115.885 164.740 182.145 164.745 ;
        POLYGON 115.315 164.740 115.315 164.400 114.370 164.400 ;
        RECT 115.315 164.680 182.145 164.740 ;
        POLYGON 182.145 164.745 182.315 164.680 182.145 164.680 ;
        POLYGON 182.600 164.745 182.600 164.680 182.495 164.680 ;
        RECT 182.600 164.680 210.185 164.745 ;
        RECT 115.315 164.655 182.315 164.680 ;
        POLYGON 182.315 164.680 182.380 164.655 182.315 164.655 ;
        POLYGON 182.495 164.680 182.495 164.655 182.455 164.655 ;
        RECT 182.495 164.655 210.185 164.680 ;
        RECT 115.315 164.645 182.380 164.655 ;
        POLYGON 182.380 164.655 182.405 164.645 182.380 164.645 ;
        POLYGON 182.455 164.655 182.455 164.645 182.440 164.645 ;
        RECT 182.455 164.645 210.185 164.655 ;
        RECT 115.315 164.635 182.405 164.645 ;
        POLYGON 182.405 164.645 182.425 164.635 182.405 164.635 ;
        POLYGON 182.440 164.645 182.440 164.640 182.430 164.640 ;
        RECT 182.440 164.640 210.185 164.645 ;
        POLYGON 182.430 164.640 182.430 164.635 182.425 164.635 ;
        RECT 182.430 164.635 210.185 164.640 ;
        RECT 115.315 164.555 210.185 164.635 ;
        POLYGON 210.185 164.825 210.930 164.825 210.185 164.555 ;
        POLYGON 222.500 164.825 222.950 164.825 222.950 164.555 ;
        RECT 222.950 164.555 232.570 164.825 ;
        RECT 115.315 164.400 208.410 164.555 ;
        POLYGON 114.370 164.400 114.370 163.545 112.015 163.545 ;
        RECT 114.370 163.910 208.410 164.400 ;
        POLYGON 208.410 164.555 210.185 164.555 208.410 163.910 ;
        POLYGON 222.950 164.555 224.015 164.555 224.015 163.910 ;
        RECT 224.015 163.925 232.570 164.555 ;
        POLYGON 232.570 168.870 239.645 163.925 232.570 163.925 ;
        POLYGON 261.485 168.870 263.770 168.870 263.770 168.435 ;
        RECT 263.770 168.435 303.120 168.870 ;
        POLYGON 263.770 168.435 263.785 168.435 263.785 168.430 ;
        RECT 263.785 168.430 303.120 168.435 ;
        POLYGON 263.785 168.430 267.050 168.430 267.050 167.695 ;
        RECT 267.050 167.695 303.120 168.430 ;
        POLYGON 267.050 167.695 270.250 167.695 270.250 166.860 ;
        RECT 270.250 166.860 303.120 167.695 ;
        POLYGON 270.250 166.860 271.625 166.860 271.625 166.450 ;
        RECT 271.625 166.450 303.120 166.860 ;
        POLYGON 271.630 166.450 273.360 166.450 273.360 165.930 ;
        RECT 273.360 165.930 303.120 166.450 ;
        POLYGON 273.360 165.930 276.385 165.930 276.385 164.905 ;
        RECT 276.385 164.905 303.120 165.930 ;
        POLYGON 276.385 164.905 278.950 164.905 278.950 163.925 ;
        RECT 278.950 163.925 303.120 164.905 ;
        RECT 224.015 163.910 239.645 163.925 ;
        RECT 114.370 163.905 208.395 163.910 ;
        POLYGON 208.395 163.910 208.410 163.910 208.395 163.905 ;
        POLYGON 224.015 163.910 224.020 163.910 224.020 163.905 ;
        RECT 224.020 163.905 239.645 163.910 ;
        RECT 114.370 163.895 208.370 163.905 ;
        POLYGON 208.370 163.905 208.395 163.905 208.370 163.895 ;
        POLYGON 224.020 163.905 224.040 163.905 224.040 163.895 ;
        RECT 224.040 163.895 239.645 163.905 ;
        RECT 114.370 163.545 207.065 163.895 ;
        POLYGON 112.015 163.545 112.015 163.230 111.245 163.230 ;
        RECT 112.015 163.420 207.065 163.545 ;
        POLYGON 207.065 163.895 208.370 163.895 207.065 163.420 ;
        POLYGON 224.040 163.895 224.825 163.895 224.825 163.420 ;
        RECT 224.825 163.420 239.645 163.895 ;
        RECT 112.015 163.230 206.565 163.420 ;
        RECT 70.370 163.175 84.765 163.230 ;
        POLYGON 84.765 163.230 84.855 163.230 84.765 163.175 ;
        POLYGON 111.245 163.230 111.245 163.175 111.110 163.175 ;
        RECT 111.245 163.215 206.565 163.230 ;
        POLYGON 206.565 163.420 207.065 163.420 206.565 163.215 ;
        POLYGON 224.825 163.420 225.165 163.420 225.165 163.215 ;
        RECT 225.165 163.215 239.645 163.420 ;
        RECT 111.245 163.175 205.290 163.215 ;
        RECT 70.370 162.825 84.180 163.175 ;
        POLYGON 84.180 163.175 84.765 163.175 84.180 162.825 ;
        POLYGON 111.110 163.175 111.110 162.825 110.255 162.825 ;
        RECT 111.110 162.825 205.290 163.175 ;
        RECT 70.370 162.570 81.220 162.825 ;
        POLYGON 68.665 162.570 68.665 160.555 66.125 160.555 ;
        RECT 68.665 160.850 81.220 162.570 ;
        POLYGON 81.220 162.825 84.180 162.825 81.220 160.850 ;
        POLYGON 110.255 162.825 110.255 162.520 109.510 162.520 ;
        RECT 110.255 162.695 205.290 162.825 ;
        POLYGON 205.290 163.215 206.565 163.215 205.290 162.695 ;
        POLYGON 225.165 163.215 226.020 163.215 226.020 162.695 ;
        RECT 226.020 162.695 239.645 163.215 ;
        RECT 110.255 162.520 203.920 162.695 ;
        POLYGON 109.510 162.520 109.510 161.980 108.190 161.980 ;
        RECT 109.510 162.135 203.920 162.520 ;
        POLYGON 203.920 162.695 205.290 162.695 203.920 162.135 ;
        POLYGON 226.020 162.695 226.945 162.695 226.945 162.135 ;
        RECT 226.945 162.135 239.645 162.695 ;
        RECT 109.510 161.980 203.450 162.135 ;
        POLYGON 108.190 161.980 108.190 161.930 108.080 161.930 ;
        RECT 108.190 161.945 203.450 161.980 ;
        POLYGON 203.450 162.135 203.920 162.135 203.450 161.945 ;
        POLYGON 226.945 162.135 227.260 162.135 227.260 161.945 ;
        RECT 227.260 161.945 239.645 162.135 ;
        RECT 108.190 161.935 203.425 161.945 ;
        POLYGON 203.425 161.945 203.450 161.945 203.425 161.935 ;
        POLYGON 227.260 161.945 227.280 161.945 227.280 161.935 ;
        RECT 227.280 161.935 239.645 161.945 ;
        RECT 108.190 161.930 203.240 161.935 ;
        POLYGON 108.080 161.930 108.080 160.850 105.705 160.850 ;
        RECT 108.080 161.860 203.240 161.930 ;
        POLYGON 203.240 161.935 203.425 161.935 203.240 161.860 ;
        POLYGON 227.280 161.935 227.385 161.935 227.385 161.860 ;
        RECT 227.385 161.860 239.645 161.935 ;
        RECT 108.080 161.395 202.215 161.860 ;
        POLYGON 202.215 161.860 203.240 161.860 202.215 161.395 ;
        POLYGON 227.385 161.860 228.060 161.860 228.060 161.395 ;
        RECT 228.060 161.395 239.645 161.860 ;
        RECT 108.080 160.850 199.850 161.395 ;
        RECT 68.665 160.555 78.570 160.850 ;
        POLYGON 66.125 160.555 66.125 158.575 63.630 158.575 ;
        RECT 66.125 159.085 78.570 160.555 ;
        POLYGON 78.570 160.850 81.220 160.850 78.570 159.085 ;
        POLYGON 105.705 160.850 105.705 160.255 104.395 160.255 ;
        RECT 105.705 160.320 199.850 160.850 ;
        POLYGON 199.850 161.395 202.215 161.395 199.850 160.320 ;
        POLYGON 228.060 161.395 229.620 161.395 229.620 160.320 ;
        RECT 229.620 160.320 239.645 161.395 ;
        RECT 105.705 160.255 199.510 160.320 ;
        POLYGON 104.390 160.255 104.390 159.965 103.815 159.965 ;
        RECT 104.390 160.165 199.510 160.255 ;
        POLYGON 199.510 160.320 199.850 160.320 199.510 160.165 ;
        POLYGON 229.620 160.320 229.845 160.320 229.845 160.165 ;
        RECT 229.845 160.165 239.645 160.320 ;
        RECT 104.390 160.135 199.450 160.165 ;
        POLYGON 199.450 160.165 199.510 160.165 199.450 160.135 ;
        POLYGON 229.845 160.165 229.885 160.165 229.885 160.135 ;
        RECT 229.885 160.135 239.645 160.165 ;
        RECT 104.390 160.000 199.185 160.135 ;
        POLYGON 199.185 160.135 199.450 160.135 199.185 160.000 ;
        POLYGON 229.885 160.135 230.085 160.135 230.085 160.000 ;
        RECT 230.085 160.000 239.645 160.135 ;
        RECT 104.390 159.965 196.725 160.000 ;
        POLYGON 103.815 159.965 103.815 159.085 102.080 159.085 ;
        RECT 103.815 159.085 196.725 159.965 ;
        RECT 66.125 158.575 77.825 159.085 ;
        POLYGON 63.630 158.575 63.630 158.410 63.450 158.410 ;
        RECT 63.630 158.535 77.825 158.575 ;
        POLYGON 77.825 159.085 78.570 159.085 77.825 158.535 ;
        POLYGON 102.080 159.085 102.080 159.000 101.910 159.000 ;
        RECT 102.080 159.000 196.725 159.085 ;
        POLYGON 101.910 159.000 101.910 158.535 100.985 158.535 ;
        RECT 101.910 158.760 196.725 159.000 ;
        POLYGON 196.725 160.000 199.185 160.000 196.725 158.760 ;
        POLYGON 230.085 160.000 231.885 160.000 231.885 158.760 ;
        RECT 231.885 158.760 239.645 160.000 ;
        RECT 101.910 158.535 196.240 158.760 ;
        RECT 63.630 158.410 77.450 158.535 ;
        POLYGON 63.450 158.410 63.450 156.200 60.990 156.200 ;
        RECT 63.450 158.255 77.450 158.410 ;
        POLYGON 77.450 158.535 77.825 158.535 77.450 158.255 ;
        POLYGON 100.985 158.535 100.985 158.255 100.430 158.255 ;
        RECT 100.985 158.515 196.240 158.535 ;
        POLYGON 196.240 158.760 196.725 158.760 196.240 158.515 ;
        POLYGON 231.885 158.760 232.240 158.760 232.240 158.515 ;
        RECT 232.240 158.580 239.645 158.760 ;
        POLYGON 239.645 163.925 246.385 158.580 239.645 158.580 ;
        POLYGON 278.950 163.925 279.320 163.925 279.320 163.785 ;
        RECT 279.320 163.785 303.120 163.925 ;
        POLYGON 279.320 163.785 279.355 163.785 279.355 163.770 ;
        RECT 279.355 163.770 303.120 163.785 ;
        POLYGON 279.355 163.770 282.160 163.770 282.160 162.575 ;
        RECT 282.160 162.575 303.120 163.770 ;
        POLYGON 282.160 162.575 284.905 162.575 284.905 161.270 ;
        RECT 284.905 161.270 303.120 162.575 ;
        POLYGON 284.905 161.270 286.945 161.270 286.945 160.200 ;
        RECT 286.945 160.200 303.120 161.270 ;
        POLYGON 286.945 160.200 287.555 160.200 287.555 159.880 ;
        RECT 287.555 159.880 303.120 160.200 ;
        POLYGON 287.555 159.880 289.785 159.880 289.785 158.580 ;
        RECT 289.785 158.580 303.120 159.880 ;
        RECT 232.240 158.515 246.385 158.580 ;
        RECT 100.985 158.400 196.015 158.515 ;
        POLYGON 196.015 158.515 196.240 158.515 196.015 158.400 ;
        POLYGON 232.240 158.515 232.405 158.515 232.405 158.400 ;
        RECT 232.405 158.400 246.385 158.515 ;
        RECT 100.985 158.325 195.865 158.400 ;
        POLYGON 195.865 158.400 196.015 158.400 195.865 158.325 ;
        POLYGON 232.405 158.400 232.515 158.400 232.515 158.325 ;
        RECT 232.515 158.325 246.385 158.400 ;
        RECT 100.985 158.290 195.790 158.325 ;
        POLYGON 195.790 158.325 195.860 158.325 195.790 158.290 ;
        POLYGON 232.515 158.325 232.570 158.325 232.570 158.290 ;
        RECT 232.570 158.290 246.385 158.325 ;
        RECT 100.985 158.275 195.765 158.290 ;
        POLYGON 195.765 158.290 195.790 158.290 195.765 158.275 ;
        POLYGON 232.570 158.290 232.590 158.290 232.590 158.275 ;
        RECT 232.590 158.275 246.385 158.290 ;
        RECT 100.985 158.255 195.715 158.275 ;
        RECT 63.450 156.200 74.595 158.255 ;
        POLYGON 60.990 156.200 60.990 154.185 58.745 154.185 ;
        RECT 60.990 156.140 74.595 156.200 ;
        POLYGON 74.595 158.255 77.450 158.255 74.595 156.140 ;
        POLYGON 100.430 158.255 100.430 158.165 100.250 158.165 ;
        RECT 100.430 158.250 195.715 158.255 ;
        POLYGON 195.715 158.275 195.760 158.275 195.715 158.250 ;
        POLYGON 232.590 158.275 232.625 158.275 232.625 158.250 ;
        RECT 232.625 158.250 246.385 158.275 ;
        RECT 100.430 158.235 195.685 158.250 ;
        POLYGON 195.685 158.250 195.710 158.250 195.685 158.235 ;
        POLYGON 232.625 158.250 232.645 158.250 232.645 158.235 ;
        RECT 232.645 158.235 246.385 158.250 ;
        RECT 100.430 158.230 195.670 158.235 ;
        POLYGON 195.670 158.235 195.680 158.235 195.670 158.230 ;
        POLYGON 232.645 158.235 232.655 158.235 232.655 158.230 ;
        RECT 232.655 158.230 246.385 158.235 ;
        RECT 100.430 158.225 195.665 158.230 ;
        POLYGON 195.665 158.230 195.670 158.230 195.665 158.225 ;
        POLYGON 232.655 158.230 232.660 158.230 232.660 158.225 ;
        RECT 232.660 158.225 246.385 158.230 ;
        RECT 100.430 158.205 195.625 158.225 ;
        POLYGON 195.625 158.225 195.660 158.225 195.625 158.205 ;
        POLYGON 232.660 158.225 232.690 158.225 232.690 158.205 ;
        RECT 232.690 158.205 246.385 158.225 ;
        RECT 100.430 158.180 195.620 158.205 ;
        POLYGON 232.690 158.205 232.700 158.205 232.700 158.200 ;
        RECT 232.700 158.200 246.385 158.205 ;
        POLYGON 195.620 158.200 195.660 158.180 195.620 158.180 ;
        POLYGON 232.700 158.200 232.725 158.200 232.725 158.180 ;
        RECT 232.725 158.180 246.385 158.200 ;
        RECT 100.430 158.175 195.660 158.180 ;
        POLYGON 195.660 158.180 195.665 158.175 195.660 158.175 ;
        POLYGON 232.725 158.180 232.735 158.180 232.735 158.175 ;
        RECT 232.735 158.175 246.385 158.180 ;
        RECT 100.430 158.165 195.665 158.175 ;
        POLYGON 195.665 158.175 195.680 158.165 195.665 158.165 ;
        POLYGON 232.735 158.175 232.750 158.175 232.750 158.165 ;
        RECT 232.750 158.165 246.385 158.175 ;
        POLYGON 100.250 158.165 100.250 157.000 98.180 157.000 ;
        RECT 100.250 158.160 195.680 158.165 ;
        POLYGON 195.680 158.165 195.685 158.160 195.680 158.160 ;
        POLYGON 232.750 158.165 232.755 158.165 232.755 158.160 ;
        RECT 232.755 158.160 246.385 158.165 ;
        RECT 100.250 158.145 195.685 158.160 ;
        POLYGON 195.685 158.160 195.710 158.145 195.685 158.145 ;
        POLYGON 232.755 158.160 232.780 158.160 232.780 158.145 ;
        RECT 232.780 158.145 246.385 158.160 ;
        RECT 100.250 158.140 195.710 158.145 ;
        POLYGON 195.710 158.145 195.715 158.140 195.710 158.140 ;
        POLYGON 232.780 158.145 232.785 158.145 232.785 158.140 ;
        RECT 232.785 158.140 246.385 158.145 ;
        RECT 100.250 158.110 195.715 158.140 ;
        POLYGON 195.715 158.140 195.760 158.110 195.715 158.110 ;
        POLYGON 232.785 158.140 232.830 158.140 232.830 158.110 ;
        RECT 232.830 158.110 246.385 158.140 ;
        RECT 100.250 158.105 195.760 158.110 ;
        POLYGON 195.760 158.110 195.765 158.105 195.760 158.105 ;
        POLYGON 232.830 158.110 232.835 158.110 232.835 158.105 ;
        RECT 232.835 158.105 246.385 158.110 ;
        RECT 100.250 158.045 195.765 158.105 ;
        POLYGON 195.765 158.105 195.860 158.045 195.765 158.045 ;
        POLYGON 232.835 158.105 232.925 158.105 232.925 158.045 ;
        RECT 232.925 158.045 246.385 158.105 ;
        RECT 100.250 157.965 195.860 158.045 ;
        POLYGON 195.860 158.045 195.985 157.965 195.860 157.965 ;
        POLYGON 232.925 158.045 233.040 158.045 233.040 157.965 ;
        RECT 233.040 157.965 246.385 158.045 ;
        RECT 100.250 157.000 195.985 157.965 ;
        POLYGON 98.180 157.000 98.180 156.140 96.650 156.140 ;
        RECT 98.180 156.940 195.985 157.000 ;
        POLYGON 195.985 157.965 197.580 156.940 195.985 156.940 ;
        POLYGON 233.040 157.965 233.680 157.965 233.680 157.525 ;
        RECT 233.680 157.525 246.385 157.965 ;
        POLYGON 233.680 157.525 234.430 157.525 234.430 156.940 ;
        RECT 234.430 156.940 246.385 157.525 ;
        RECT 98.180 156.140 197.580 156.940 ;
        RECT 60.990 155.050 73.125 156.140 ;
        POLYGON 73.125 156.140 74.595 156.140 73.125 155.050 ;
        POLYGON 96.650 156.140 96.650 155.890 96.205 155.890 ;
        RECT 96.650 155.890 197.580 156.140 ;
        POLYGON 96.205 155.890 96.205 155.675 95.860 155.675 ;
        RECT 96.205 155.675 197.580 155.890 ;
        POLYGON 95.860 155.675 95.860 155.050 94.855 155.050 ;
        RECT 95.860 155.645 197.580 155.675 ;
        POLYGON 197.580 156.940 199.410 155.645 197.580 155.645 ;
        POLYGON 234.430 156.940 236.090 156.940 236.090 155.645 ;
        RECT 236.090 155.645 246.385 156.940 ;
        RECT 95.860 155.280 199.410 155.645 ;
        POLYGON 199.410 155.645 199.925 155.280 199.410 155.280 ;
        POLYGON 236.090 155.645 236.555 155.645 236.555 155.280 ;
        RECT 236.555 155.280 246.385 155.645 ;
        RECT 95.860 155.050 199.925 155.280 ;
        RECT 60.990 154.185 71.385 155.050 ;
        POLYGON 58.745 154.185 58.745 152.845 57.250 152.845 ;
        RECT 58.745 153.625 71.385 154.185 ;
        POLYGON 71.385 155.050 73.125 155.050 71.385 153.625 ;
        POLYGON 94.855 155.050 94.855 153.630 92.570 153.630 ;
        RECT 94.855 154.830 199.925 155.050 ;
        POLYGON 199.925 155.280 200.505 154.830 199.925 154.830 ;
        POLYGON 236.555 155.280 237.135 155.280 237.135 154.830 ;
        RECT 237.135 154.830 246.385 155.280 ;
        RECT 94.855 153.630 200.505 154.830 ;
        POLYGON 92.570 153.630 92.570 153.625 92.560 153.625 ;
        RECT 92.570 153.625 200.505 153.630 ;
        RECT 58.745 152.845 70.370 153.625 ;
        POLYGON 57.250 152.845 57.250 152.305 56.720 152.305 ;
        RECT 57.250 152.790 70.370 152.845 ;
        POLYGON 70.370 153.625 71.385 153.625 70.370 152.790 ;
        POLYGON 92.560 153.625 92.560 153.440 92.270 153.440 ;
        RECT 92.560 153.535 200.505 153.625 ;
        POLYGON 200.505 154.830 202.165 153.535 200.505 153.535 ;
        POLYGON 237.135 154.830 238.795 154.830 238.795 153.535 ;
        RECT 238.795 153.535 246.385 154.830 ;
        RECT 92.560 153.440 202.165 153.535 ;
        POLYGON 92.270 153.440 92.270 152.790 91.320 152.790 ;
        RECT 92.270 152.790 202.165 153.440 ;
        RECT 57.250 152.305 68.665 152.790 ;
        POLYGON 56.720 152.305 56.720 150.475 54.910 150.475 ;
        RECT 56.720 151.390 68.665 152.305 ;
        POLYGON 68.665 152.790 70.370 152.790 68.665 151.390 ;
        POLYGON 91.320 152.790 91.320 151.850 89.950 151.850 ;
        RECT 91.320 151.850 202.165 152.790 ;
        POLYGON 89.950 151.850 89.950 151.390 89.275 151.390 ;
        RECT 89.950 151.705 202.165 151.850 ;
        POLYGON 202.165 153.535 204.295 151.705 202.165 151.705 ;
        POLYGON 238.795 153.535 239.645 153.535 239.645 152.875 ;
        RECT 239.645 152.875 246.385 153.535 ;
        POLYGON 239.645 152.875 239.820 152.875 239.820 152.740 ;
        RECT 239.820 152.850 246.385 152.875 ;
        POLYGON 246.385 158.580 252.765 152.850 246.385 152.850 ;
        POLYGON 289.785 158.580 290.105 158.580 290.105 158.395 ;
        RECT 290.105 158.395 303.120 158.580 ;
        POLYGON 290.105 158.395 292.555 158.395 292.555 156.825 ;
        RECT 292.555 156.825 303.120 158.395 ;
        POLYGON 292.555 156.825 294.380 156.825 294.380 155.530 ;
        RECT 294.380 155.530 303.120 156.825 ;
        POLYGON 294.380 155.530 294.895 155.530 294.895 155.165 ;
        RECT 294.895 155.165 303.120 155.530 ;
        POLYGON 294.895 155.165 297.130 155.165 297.130 153.420 ;
        RECT 297.130 153.420 303.120 155.165 ;
        POLYGON 297.130 153.420 297.790 153.420 297.790 152.850 ;
        RECT 297.790 152.850 303.120 153.420 ;
        RECT 239.820 152.740 252.765 152.850 ;
        POLYGON 239.820 152.740 240.995 152.740 240.995 151.705 ;
        RECT 240.995 151.705 252.765 152.740 ;
        RECT 89.950 151.390 204.295 151.705 ;
        RECT 56.720 150.720 67.850 151.390 ;
        POLYGON 67.850 151.390 68.665 151.390 67.850 150.720 ;
        POLYGON 89.275 151.390 89.275 150.825 88.450 150.825 ;
        RECT 89.275 150.825 204.295 151.390 ;
        POLYGON 88.450 150.825 88.450 150.720 88.310 150.720 ;
        RECT 88.450 150.720 204.295 150.825 ;
        RECT 56.720 150.475 66.125 150.720 ;
        POLYGON 54.910 150.475 54.910 148.865 53.325 148.865 ;
        RECT 54.910 149.150 66.125 150.475 ;
        POLYGON 66.125 150.720 67.850 150.720 66.125 149.150 ;
        POLYGON 88.310 150.720 88.310 149.150 86.225 149.150 ;
        RECT 88.310 149.890 204.295 150.720 ;
        POLYGON 204.295 151.705 206.205 149.890 204.295 149.890 ;
        POLYGON 240.995 151.705 243.060 151.705 243.060 149.890 ;
        RECT 243.060 149.890 252.765 151.705 ;
        RECT 88.310 149.790 206.205 149.890 ;
        POLYGON 206.205 149.890 206.310 149.790 206.205 149.790 ;
        POLYGON 243.060 149.890 243.175 149.890 243.175 149.790 ;
        RECT 243.175 149.790 252.765 149.890 ;
        RECT 88.310 149.410 206.310 149.790 ;
        POLYGON 206.310 149.790 206.680 149.410 206.310 149.410 ;
        POLYGON 243.175 149.790 243.605 149.790 243.605 149.410 ;
        RECT 243.605 149.410 252.765 149.790 ;
        RECT 88.310 149.150 206.680 149.410 ;
        RECT 54.910 148.865 63.630 149.150 ;
        POLYGON 53.325 148.865 53.325 147.480 51.955 147.480 ;
        RECT 53.325 147.480 63.630 148.865 ;
        POLYGON 51.955 147.480 51.955 146.750 51.235 146.750 ;
        RECT 51.955 146.885 63.630 147.480 ;
        POLYGON 63.630 149.150 66.125 149.150 63.630 146.885 ;
        POLYGON 86.225 149.150 86.225 148.120 84.855 148.120 ;
        RECT 86.225 148.120 206.680 149.150 ;
        POLYGON 84.855 148.120 84.855 148.050 84.765 148.050 ;
        RECT 84.855 148.050 206.680 148.120 ;
        POLYGON 84.765 148.050 84.765 147.570 84.180 147.570 ;
        RECT 84.765 147.990 206.680 148.050 ;
        POLYGON 206.680 149.410 208.060 147.990 206.680 147.990 ;
        POLYGON 243.605 149.410 245.220 149.410 245.220 147.990 ;
        RECT 245.220 147.990 252.765 149.410 ;
        RECT 84.765 147.570 208.060 147.990 ;
        POLYGON 84.180 147.570 84.180 146.885 83.350 146.885 ;
        RECT 84.180 146.885 208.060 147.570 ;
        RECT 51.955 146.750 63.450 146.885 ;
        POLYGON 51.235 146.750 51.235 146.265 50.815 146.265 ;
        RECT 51.235 146.720 63.450 146.750 ;
        POLYGON 63.450 146.885 63.630 146.885 63.450 146.720 ;
        POLYGON 83.350 146.885 83.350 146.720 83.150 146.720 ;
        RECT 83.350 146.720 208.060 146.885 ;
        RECT 51.235 146.265 62.765 146.720 ;
        POLYGON 50.815 146.265 50.815 145.210 49.890 145.210 ;
        RECT 50.815 146.100 62.765 146.265 ;
        POLYGON 62.765 146.720 63.450 146.720 62.765 146.100 ;
        POLYGON 83.150 146.720 83.150 146.100 82.400 146.100 ;
        RECT 83.150 146.325 208.060 146.720 ;
        POLYGON 208.060 147.990 209.570 146.325 208.060 146.325 ;
        POLYGON 245.220 147.990 245.680 147.990 245.680 147.590 ;
        RECT 245.680 147.590 252.765 147.990 ;
        POLYGON 245.680 147.590 246.385 147.590 246.385 146.895 ;
        RECT 246.385 146.895 252.765 147.590 ;
        POLYGON 246.385 146.895 246.960 146.895 246.960 146.325 ;
        RECT 246.960 146.760 252.765 146.895 ;
        POLYGON 252.765 152.850 258.775 146.760 252.765 146.760 ;
        POLYGON 297.790 152.850 299.260 152.850 299.260 151.590 ;
        RECT 299.260 151.590 303.120 152.850 ;
        POLYGON 299.260 151.590 301.275 151.590 301.275 149.680 ;
        RECT 301.275 149.680 303.120 151.590 ;
        POLYGON 301.275 149.680 301.645 149.680 301.645 149.300 ;
        RECT 301.645 149.300 303.120 149.680 ;
        POLYGON 301.645 149.300 303.025 149.300 303.025 147.885 ;
        RECT 303.025 147.885 303.120 149.300 ;
        POLYGON 303.025 147.885 303.120 147.885 303.120 147.780 ;
        RECT 246.960 146.325 258.775 146.760 ;
        RECT 83.150 146.100 209.570 146.325 ;
        RECT 50.815 145.210 60.990 146.100 ;
        POLYGON 49.890 145.210 49.890 144.415 49.195 144.415 ;
        RECT 49.890 144.415 60.990 145.210 ;
        POLYGON 49.195 144.415 49.195 143.880 48.725 143.880 ;
        RECT 49.195 144.320 60.990 144.415 ;
        POLYGON 60.990 146.100 62.765 146.100 60.990 144.320 ;
        POLYGON 82.400 146.100 82.400 145.125 81.220 145.125 ;
        RECT 82.400 145.125 209.570 146.100 ;
        POLYGON 81.220 145.125 81.220 144.320 80.330 144.320 ;
        RECT 81.220 144.750 209.570 145.125 ;
        POLYGON 209.570 146.325 210.865 144.750 209.570 144.750 ;
        POLYGON 246.960 146.325 248.550 146.325 248.550 144.750 ;
        RECT 248.550 144.750 258.775 146.325 ;
        RECT 81.220 144.320 210.865 144.750 ;
        RECT 49.195 143.880 58.870 144.320 ;
        POLYGON 48.725 143.880 48.725 143.600 48.485 143.600 ;
        RECT 48.725 143.600 58.870 143.880 ;
        POLYGON 48.485 143.600 48.485 143.585 48.470 143.585 ;
        RECT 48.485 143.585 58.870 143.600 ;
        POLYGON 48.470 143.585 48.470 140.310 45.605 140.310 ;
        RECT 48.470 142.200 58.870 143.585 ;
        POLYGON 58.870 144.320 60.990 144.320 58.870 142.200 ;
        POLYGON 80.330 144.320 80.330 142.730 78.570 142.730 ;
        RECT 80.330 143.405 210.865 144.320 ;
        POLYGON 210.865 144.750 211.840 143.405 210.865 143.405 ;
        POLYGON 248.550 144.750 249.910 144.750 249.910 143.405 ;
        RECT 249.910 143.405 258.775 144.750 ;
        RECT 80.330 143.230 211.840 143.405 ;
        POLYGON 211.840 143.405 211.970 143.230 211.840 143.230 ;
        POLYGON 249.910 143.405 250.085 143.405 250.085 143.230 ;
        RECT 250.085 143.230 258.775 143.405 ;
        RECT 80.330 142.730 211.970 143.230 ;
        POLYGON 78.570 142.730 78.570 142.200 77.985 142.200 ;
        RECT 78.570 142.475 211.970 142.730 ;
        POLYGON 211.970 143.230 212.460 142.475 211.970 142.475 ;
        POLYGON 250.085 143.230 250.850 143.230 250.850 142.475 ;
        RECT 250.850 142.475 258.775 143.230 ;
        RECT 78.570 142.200 212.460 142.475 ;
        RECT 48.470 142.060 58.745 142.200 ;
        POLYGON 58.745 142.200 58.870 142.200 58.745 142.060 ;
        POLYGON 77.985 142.200 77.985 142.060 77.830 142.060 ;
        RECT 77.985 142.060 212.460 142.200 ;
        RECT 48.470 140.420 57.250 142.060 ;
        POLYGON 57.250 142.060 58.745 142.060 57.250 140.420 ;
        POLYGON 77.830 142.060 77.830 142.055 77.825 142.055 ;
        RECT 77.830 142.055 212.460 142.060 ;
        POLYGON 77.825 142.055 77.825 141.685 77.450 141.685 ;
        RECT 77.825 141.715 212.460 142.055 ;
        POLYGON 212.460 142.475 212.915 141.715 212.460 141.715 ;
        POLYGON 250.850 142.475 251.240 142.475 251.240 142.090 ;
        RECT 251.240 142.090 258.775 142.475 ;
        POLYGON 251.240 142.090 251.575 142.090 251.575 141.715 ;
        RECT 251.575 141.715 258.775 142.090 ;
        RECT 77.825 141.685 212.915 141.715 ;
        POLYGON 77.450 141.685 77.450 140.420 76.175 140.420 ;
        RECT 77.450 140.950 212.915 141.685 ;
        POLYGON 212.915 141.715 213.335 140.950 212.915 140.950 ;
        POLYGON 251.575 141.715 252.260 141.715 252.260 140.950 ;
        RECT 252.260 140.950 258.775 141.715 ;
        RECT 77.450 140.420 213.335 140.950 ;
        RECT 48.470 140.310 56.720 140.420 ;
        POLYGON 45.605 140.310 45.605 133.550 40.375 133.550 ;
        RECT 45.605 139.840 56.720 140.310 ;
        POLYGON 56.720 140.420 57.250 140.420 56.720 139.840 ;
        POLYGON 76.175 140.420 76.175 139.840 75.590 139.840 ;
        RECT 76.175 140.170 213.335 140.420 ;
        POLYGON 213.335 140.950 213.730 140.170 213.335 140.170 ;
        POLYGON 252.260 140.950 252.765 140.950 252.765 140.390 ;
        RECT 252.765 140.390 258.775 140.950 ;
        POLYGON 252.765 140.390 252.960 140.390 252.960 140.170 ;
        RECT 252.960 140.325 258.775 140.390 ;
        POLYGON 258.775 146.760 264.405 140.325 258.775 140.325 ;
        RECT 252.960 140.170 264.405 140.325 ;
        RECT 76.175 140.095 213.730 140.170 ;
        POLYGON 213.730 140.170 213.760 140.095 213.730 140.095 ;
        POLYGON 252.960 140.170 253.025 140.170 253.025 140.100 ;
        RECT 253.025 140.095 264.405 140.170 ;
        RECT 76.175 139.840 213.760 140.095 ;
        RECT 45.605 138.050 55.085 139.840 ;
        POLYGON 55.085 139.840 56.720 139.840 55.085 138.050 ;
        POLYGON 75.590 139.840 75.590 138.855 74.595 138.855 ;
        RECT 75.590 138.855 213.760 139.840 ;
        POLYGON 74.595 138.850 74.595 138.050 73.850 138.050 ;
        RECT 74.595 138.550 213.760 138.855 ;
        POLYGON 213.760 140.095 214.440 138.550 213.760 138.550 ;
        POLYGON 253.025 140.095 254.415 140.095 254.415 138.550 ;
        RECT 254.415 138.550 264.405 140.095 ;
        RECT 74.595 138.050 214.440 138.550 ;
        RECT 45.605 137.840 54.910 138.050 ;
        POLYGON 54.910 138.050 55.085 138.050 54.910 137.840 ;
        POLYGON 73.850 138.050 73.850 137.840 73.650 137.840 ;
        RECT 73.850 137.840 214.440 138.050 ;
        RECT 45.605 135.945 53.325 137.840 ;
        POLYGON 53.325 137.840 54.910 137.840 53.325 135.945 ;
        POLYGON 73.650 137.840 73.650 137.275 73.125 137.275 ;
        RECT 73.650 137.275 214.440 137.840 ;
        POLYGON 73.125 137.275 73.125 135.945 71.885 135.945 ;
        RECT 73.125 136.815 214.440 137.275 ;
        POLYGON 214.440 138.550 215.070 136.815 214.440 136.815 ;
        POLYGON 254.415 138.550 255.970 138.550 255.970 136.815 ;
        RECT 255.970 136.815 264.405 138.550 ;
        RECT 73.125 136.325 215.070 136.815 ;
        POLYGON 215.070 136.815 215.225 136.325 215.070 136.325 ;
        POLYGON 255.970 136.815 256.410 136.815 256.410 136.325 ;
        RECT 256.410 136.325 264.405 136.815 ;
        RECT 73.125 135.945 215.225 136.325 ;
        RECT 45.605 134.310 51.955 135.945 ;
        POLYGON 51.955 135.945 53.325 135.945 51.955 134.310 ;
        POLYGON 71.885 135.940 71.885 135.405 71.385 135.405 ;
        RECT 71.885 135.835 215.225 135.945 ;
        POLYGON 215.225 136.325 215.345 135.835 215.225 135.835 ;
        POLYGON 256.410 136.325 256.485 136.325 256.485 136.245 ;
        RECT 256.485 136.245 264.405 136.325 ;
        POLYGON 256.485 136.245 256.810 136.245 256.810 135.835 ;
        RECT 256.810 135.835 264.405 136.245 ;
        RECT 71.885 135.405 215.345 135.835 ;
        POLYGON 71.385 135.405 71.385 134.310 70.455 134.310 ;
        RECT 71.385 135.340 215.345 135.405 ;
        POLYGON 215.345 135.835 215.445 135.340 215.345 135.340 ;
        POLYGON 256.810 135.835 257.200 135.835 257.200 135.340 ;
        RECT 257.200 135.340 264.405 135.835 ;
        RECT 71.385 134.820 215.445 135.340 ;
        POLYGON 215.445 135.340 215.515 134.820 215.445 134.820 ;
        POLYGON 257.200 135.340 257.615 135.340 257.615 134.820 ;
        RECT 257.615 134.820 264.405 135.340 ;
        RECT 71.385 134.310 215.515 134.820 ;
        RECT 45.605 133.685 51.435 134.310 ;
        POLYGON 51.435 134.310 51.955 134.310 51.435 133.685 ;
        POLYGON 70.455 134.310 70.455 134.210 70.370 134.210 ;
        RECT 70.455 134.265 215.515 134.310 ;
        POLYGON 215.515 134.820 215.560 134.265 215.515 134.265 ;
        POLYGON 257.615 134.820 258.055 134.820 258.055 134.265 ;
        RECT 258.055 134.265 264.405 134.820 ;
        RECT 70.455 134.210 215.560 134.265 ;
        POLYGON 70.370 134.210 70.370 133.685 69.925 133.685 ;
        RECT 70.370 133.685 215.560 134.210 ;
        RECT 45.605 133.550 51.235 133.685 ;
        POLYGON 40.375 133.550 40.375 126.490 35.560 126.490 ;
        RECT 40.375 133.425 51.235 133.550 ;
        POLYGON 51.235 133.685 51.435 133.685 51.235 133.425 ;
        POLYGON 69.925 133.685 69.925 133.425 69.700 133.425 ;
        RECT 69.925 133.665 215.560 133.685 ;
        POLYGON 215.560 134.265 215.585 133.665 215.560 133.665 ;
        RECT 69.925 133.425 215.585 133.665 ;
        RECT 40.375 132.875 50.815 133.425 ;
        POLYGON 50.815 133.425 51.235 133.425 50.815 132.875 ;
        POLYGON 69.700 133.420 69.700 132.875 69.235 132.875 ;
        RECT 69.700 132.970 215.585 133.425 ;
        POLYGON 258.055 134.265 258.775 134.265 258.775 133.360 ;
        RECT 258.775 133.570 264.405 134.265 ;
        POLYGON 264.405 140.325 269.630 133.570 264.405 133.570 ;
        RECT 258.775 133.360 269.630 133.570 ;
        RECT 69.700 132.875 215.565 132.970 ;
        RECT 40.375 131.675 49.890 132.875 ;
        POLYGON 49.890 132.875 50.815 132.875 49.890 131.675 ;
        POLYGON 69.235 132.875 69.235 132.205 68.665 132.205 ;
        RECT 69.235 132.280 215.565 132.875 ;
        POLYGON 215.565 132.970 215.585 132.970 215.565 132.280 ;
        POLYGON 258.775 133.360 259.630 133.360 259.630 132.280 ;
        RECT 259.630 132.280 269.630 133.360 ;
        RECT 69.235 132.205 215.560 132.280 ;
        POLYGON 68.665 132.205 68.665 131.675 68.260 131.675 ;
        RECT 68.665 132.180 215.560 132.205 ;
        POLYGON 215.560 132.280 215.565 132.280 215.560 132.180 ;
        POLYGON 259.630 132.280 259.710 132.280 259.710 132.180 ;
        RECT 259.710 132.180 269.630 132.280 ;
        RECT 68.665 131.690 215.535 132.180 ;
        POLYGON 215.535 132.180 215.560 132.180 215.535 131.690 ;
        POLYGON 259.710 132.180 260.100 132.180 260.100 131.690 ;
        RECT 260.100 131.690 269.630 132.180 ;
        RECT 68.665 131.675 215.515 131.690 ;
        RECT 40.375 130.770 49.195 131.675 ;
        POLYGON 49.195 131.675 49.890 131.675 49.195 130.770 ;
        POLYGON 68.260 131.675 68.260 131.135 67.850 131.135 ;
        RECT 68.260 131.420 215.515 131.675 ;
        POLYGON 215.515 131.690 215.535 131.690 215.515 131.420 ;
        POLYGON 260.100 131.690 260.310 131.690 260.310 131.425 ;
        RECT 260.310 131.420 269.630 131.690 ;
        RECT 68.260 131.135 215.490 131.420 ;
        POLYGON 215.490 131.420 215.515 131.420 215.490 131.135 ;
        POLYGON 260.310 131.420 260.540 131.420 260.540 131.135 ;
        RECT 260.540 131.135 269.630 131.420 ;
        POLYGON 67.850 131.135 67.850 130.775 67.575 130.775 ;
        RECT 67.850 130.775 215.445 131.135 ;
        RECT 40.375 130.160 48.725 130.770 ;
        POLYGON 48.725 130.770 49.195 130.770 48.725 130.160 ;
        POLYGON 67.575 130.770 67.575 130.160 67.110 130.160 ;
        RECT 67.575 130.690 215.445 130.775 ;
        POLYGON 215.445 131.135 215.490 131.135 215.445 130.690 ;
        POLYGON 260.540 131.135 260.890 131.135 260.890 130.695 ;
        RECT 260.890 130.690 269.630 131.135 ;
        RECT 67.575 130.615 215.435 130.690 ;
        POLYGON 215.435 130.690 215.445 130.690 215.435 130.615 ;
        POLYGON 260.890 130.690 260.950 130.690 260.950 130.615 ;
        RECT 260.950 130.615 269.630 130.690 ;
        RECT 67.575 130.160 215.360 130.615 ;
        RECT 40.375 129.820 48.470 130.160 ;
        POLYGON 48.470 130.160 48.725 130.160 48.470 129.820 ;
        POLYGON 67.110 130.160 67.110 129.820 66.850 129.820 ;
        RECT 67.110 130.130 215.360 130.160 ;
        POLYGON 215.360 130.615 215.435 130.615 215.360 130.130 ;
        POLYGON 260.950 130.615 261.335 130.615 261.335 130.130 ;
        RECT 261.335 130.130 269.630 130.615 ;
        RECT 67.110 130.060 215.345 130.130 ;
        POLYGON 215.345 130.130 215.360 130.130 215.345 130.060 ;
        POLYGON 261.335 130.130 261.390 130.130 261.390 130.065 ;
        RECT 261.390 130.060 269.630 130.130 ;
        RECT 67.110 129.820 215.270 130.060 ;
        RECT 40.375 129.135 47.940 129.820 ;
        POLYGON 47.940 129.820 48.470 129.820 47.940 129.135 ;
        POLYGON 66.850 129.820 66.850 129.135 66.330 129.135 ;
        RECT 66.850 129.675 215.270 129.820 ;
        POLYGON 215.270 130.060 215.345 130.060 215.270 129.675 ;
        POLYGON 261.390 130.060 261.660 130.060 261.660 129.680 ;
        RECT 261.660 129.675 269.630 130.060 ;
        RECT 66.850 129.500 215.225 129.675 ;
        POLYGON 215.225 129.675 215.270 129.675 215.225 129.500 ;
        POLYGON 261.660 129.675 261.785 129.675 261.785 129.500 ;
        RECT 261.785 129.500 269.630 129.675 ;
        RECT 66.850 129.245 215.155 129.500 ;
        POLYGON 215.155 129.500 215.225 129.500 215.155 129.245 ;
        POLYGON 261.785 129.500 261.965 129.500 261.965 129.245 ;
        RECT 261.965 129.245 269.630 129.500 ;
        RECT 66.850 129.135 215.095 129.245 ;
        RECT 40.375 126.490 45.605 129.135 ;
        POLYGON 35.560 126.490 35.560 119.145 31.170 119.145 ;
        RECT 35.560 125.825 45.605 126.490 ;
        POLYGON 45.605 129.135 47.940 129.135 45.605 125.825 ;
        POLYGON 66.330 129.135 66.330 128.865 66.125 128.865 ;
        RECT 66.330 129.035 215.095 129.135 ;
        POLYGON 215.095 129.245 215.155 129.245 215.095 129.035 ;
        POLYGON 261.965 129.245 262.110 129.245 262.110 129.035 ;
        RECT 262.110 129.035 269.630 129.245 ;
        RECT 66.330 128.975 215.070 129.035 ;
        POLYGON 215.070 129.035 215.095 129.035 215.070 128.975 ;
        POLYGON 262.110 129.035 262.155 129.035 262.155 128.975 ;
        RECT 262.155 128.975 269.630 129.035 ;
        RECT 66.330 128.865 215.025 128.975 ;
        POLYGON 66.125 128.865 66.125 125.825 64.025 125.825 ;
        RECT 66.125 128.835 215.025 128.865 ;
        POLYGON 215.025 128.975 215.070 128.975 215.025 128.835 ;
        POLYGON 262.155 128.975 262.250 128.975 262.250 128.835 ;
        RECT 262.250 128.835 269.630 128.975 ;
        RECT 66.125 128.635 214.950 128.835 ;
        POLYGON 214.950 128.835 215.025 128.835 214.950 128.635 ;
        POLYGON 262.250 128.835 262.390 128.835 262.390 128.640 ;
        RECT 262.390 128.635 269.630 128.835 ;
        RECT 66.125 128.445 214.870 128.635 ;
        POLYGON 214.870 128.635 214.950 128.635 214.870 128.445 ;
        POLYGON 262.390 128.635 262.525 128.635 262.525 128.445 ;
        RECT 262.525 128.445 269.630 128.635 ;
        RECT 66.125 128.255 214.785 128.445 ;
        POLYGON 214.785 128.445 214.870 128.445 214.785 128.255 ;
        POLYGON 262.525 128.445 262.660 128.445 262.660 128.255 ;
        RECT 262.660 128.255 269.630 128.445 ;
        RECT 66.125 127.885 214.595 128.255 ;
        POLYGON 214.595 128.255 214.785 128.255 214.595 127.885 ;
        POLYGON 262.660 128.255 262.920 128.255 262.920 127.885 ;
        RECT 262.920 127.885 269.630 128.255 ;
        RECT 66.125 127.705 214.490 127.885 ;
        POLYGON 214.490 127.885 214.595 127.885 214.490 127.705 ;
        POLYGON 262.920 127.885 263.045 127.885 263.045 127.705 ;
        RECT 263.045 127.705 269.630 127.885 ;
        RECT 66.125 127.625 214.440 127.705 ;
        POLYGON 214.440 127.705 214.490 127.705 214.440 127.625 ;
        POLYGON 263.045 127.705 263.100 127.705 263.100 127.625 ;
        RECT 263.100 127.625 269.630 127.705 ;
        RECT 66.125 127.345 214.260 127.625 ;
        POLYGON 214.260 127.625 214.440 127.625 214.260 127.345 ;
        POLYGON 263.100 127.625 263.295 127.625 263.295 127.350 ;
        RECT 263.295 127.345 269.630 127.625 ;
        RECT 66.125 126.995 214.000 127.345 ;
        POLYGON 214.000 127.345 214.260 127.345 214.000 126.995 ;
        POLYGON 263.295 127.345 263.545 127.345 263.545 126.995 ;
        RECT 263.545 126.995 269.630 127.345 ;
        RECT 66.125 126.665 213.730 126.995 ;
        POLYGON 213.730 126.995 214.000 126.995 213.730 126.665 ;
        POLYGON 263.545 126.995 263.775 126.995 263.775 126.665 ;
        RECT 263.775 126.665 269.630 126.995 ;
        RECT 66.125 126.645 213.710 126.665 ;
        POLYGON 213.710 126.665 213.730 126.665 213.710 126.645 ;
        POLYGON 263.775 126.665 263.790 126.665 263.790 126.645 ;
        RECT 263.790 126.645 269.630 126.665 ;
        RECT 66.125 126.290 213.390 126.645 ;
        POLYGON 213.390 126.645 213.710 126.645 213.390 126.290 ;
        POLYGON 263.790 126.645 264.035 126.645 264.035 126.295 ;
        RECT 264.035 126.505 269.630 126.645 ;
        POLYGON 269.630 133.570 274.450 126.505 269.630 126.505 ;
        RECT 264.035 126.290 274.450 126.505 ;
        RECT 66.125 126.235 213.335 126.290 ;
        POLYGON 213.335 126.290 213.390 126.290 213.335 126.235 ;
        POLYGON 264.035 126.290 264.075 126.290 264.075 126.240 ;
        RECT 264.075 126.235 274.450 126.290 ;
        RECT 66.125 125.935 213.040 126.235 ;
        POLYGON 213.040 126.235 213.335 126.235 213.040 125.935 ;
        POLYGON 264.075 126.235 264.285 126.235 264.285 125.940 ;
        RECT 264.285 125.935 274.450 126.235 ;
        RECT 66.125 125.825 212.915 125.935 ;
        RECT 35.560 124.435 44.630 125.825 ;
        POLYGON 44.630 125.825 45.605 125.825 44.630 124.435 ;
        POLYGON 64.025 125.825 64.025 125.255 63.630 125.255 ;
        RECT 64.025 125.815 212.915 125.825 ;
        POLYGON 212.915 125.935 213.040 125.935 212.915 125.815 ;
        POLYGON 264.285 125.935 264.370 125.935 264.370 125.815 ;
        RECT 264.370 125.815 274.450 125.935 ;
        RECT 64.025 125.565 212.650 125.815 ;
        POLYGON 212.650 125.815 212.915 125.815 212.650 125.565 ;
        POLYGON 264.370 125.815 264.405 125.815 264.405 125.770 ;
        RECT 264.405 125.770 274.450 125.815 ;
        POLYGON 264.405 125.770 264.545 125.770 264.545 125.570 ;
        RECT 264.545 125.565 274.450 125.770 ;
        RECT 64.025 125.395 212.460 125.565 ;
        POLYGON 212.460 125.565 212.650 125.565 212.460 125.395 ;
        POLYGON 264.545 125.565 264.665 125.565 264.665 125.395 ;
        RECT 264.665 125.395 274.450 125.565 ;
        RECT 64.025 125.255 212.300 125.395 ;
        POLYGON 63.630 125.255 63.630 124.990 63.450 124.990 ;
        RECT 63.630 125.250 212.300 125.255 ;
        POLYGON 212.300 125.395 212.460 125.395 212.300 125.250 ;
        POLYGON 264.665 125.395 264.765 125.395 264.765 125.255 ;
        RECT 264.765 125.250 274.450 125.395 ;
        RECT 63.630 124.990 211.970 125.250 ;
        POLYGON 63.450 124.990 63.450 124.440 63.100 124.440 ;
        RECT 63.450 124.970 211.970 124.990 ;
        POLYGON 211.970 125.250 212.300 125.250 211.970 124.970 ;
        POLYGON 264.765 125.250 264.965 125.250 264.965 124.970 ;
        RECT 264.965 124.970 274.450 125.250 ;
        RECT 63.450 124.955 211.945 124.970 ;
        POLYGON 211.945 124.970 211.970 124.970 211.945 124.955 ;
        POLYGON 264.965 124.970 264.975 124.970 264.975 124.955 ;
        RECT 264.975 124.955 274.450 124.970 ;
        RECT 63.450 124.665 211.585 124.955 ;
        POLYGON 211.585 124.955 211.945 124.955 211.585 124.665 ;
        POLYGON 264.975 124.955 265.175 124.955 265.175 124.670 ;
        RECT 265.175 124.665 274.450 124.955 ;
        RECT 63.450 124.440 211.210 124.665 ;
        RECT 35.560 119.615 41.525 124.435 ;
        POLYGON 41.525 124.435 44.630 124.435 41.525 119.615 ;
        POLYGON 63.100 124.435 63.100 123.910 62.765 123.910 ;
        RECT 63.100 124.390 211.210 124.440 ;
        POLYGON 211.210 124.665 211.585 124.665 211.210 124.390 ;
        POLYGON 265.175 124.665 265.370 124.665 265.370 124.390 ;
        RECT 265.370 124.390 274.450 124.665 ;
        RECT 63.100 124.150 210.865 124.390 ;
        POLYGON 210.865 124.390 211.210 124.390 210.865 124.150 ;
        POLYGON 265.370 124.390 265.540 124.390 265.540 124.150 ;
        RECT 265.540 124.150 274.450 124.390 ;
        RECT 63.100 124.125 210.825 124.150 ;
        POLYGON 210.825 124.150 210.860 124.150 210.825 124.125 ;
        POLYGON 265.540 124.150 265.555 124.150 265.555 124.125 ;
        RECT 265.555 124.125 274.450 124.150 ;
        RECT 63.100 123.910 210.425 124.125 ;
        POLYGON 62.765 123.910 62.765 121.105 60.990 121.105 ;
        RECT 62.765 123.875 210.425 123.910 ;
        POLYGON 210.425 124.125 210.825 124.125 210.425 123.875 ;
        POLYGON 265.555 124.125 265.730 124.125 265.730 123.875 ;
        RECT 265.730 123.875 274.450 124.125 ;
        RECT 62.765 123.630 210.015 123.875 ;
        POLYGON 210.015 123.875 210.425 123.875 210.015 123.630 ;
        POLYGON 265.730 123.875 265.900 123.875 265.900 123.635 ;
        RECT 265.900 123.630 274.450 123.875 ;
        RECT 62.765 123.400 209.580 123.630 ;
        POLYGON 209.580 123.630 210.015 123.630 209.580 123.400 ;
        POLYGON 265.900 123.630 265.950 123.630 265.950 123.565 ;
        RECT 265.950 123.565 274.450 123.630 ;
        POLYGON 265.950 123.565 266.055 123.565 266.055 123.400 ;
        RECT 266.055 123.400 274.450 123.565 ;
        RECT 62.765 123.175 209.130 123.400 ;
        POLYGON 209.130 123.400 209.580 123.400 209.130 123.175 ;
        POLYGON 266.055 123.400 266.195 123.400 266.195 123.180 ;
        RECT 266.195 123.175 274.450 123.400 ;
        RECT 62.765 122.965 208.660 123.175 ;
        POLYGON 208.660 123.175 209.130 123.175 208.660 122.965 ;
        POLYGON 266.195 123.175 266.330 123.175 266.330 122.965 ;
        RECT 266.330 122.965 274.450 123.175 ;
        RECT 62.765 122.760 208.165 122.965 ;
        POLYGON 208.165 122.965 208.660 122.965 208.165 122.760 ;
        POLYGON 266.330 122.965 266.460 122.965 266.460 122.760 ;
        RECT 266.460 122.760 274.450 122.965 ;
        RECT 62.765 122.720 208.060 122.760 ;
        POLYGON 208.060 122.760 208.165 122.760 208.060 122.720 ;
        POLYGON 266.460 122.760 266.485 122.760 266.485 122.725 ;
        RECT 266.485 122.720 274.450 122.760 ;
        RECT 62.765 122.560 207.645 122.720 ;
        POLYGON 207.645 122.720 208.060 122.720 207.645 122.560 ;
        POLYGON 266.485 122.720 266.590 122.720 266.590 122.560 ;
        RECT 266.590 122.560 274.450 122.720 ;
        RECT 62.765 122.190 206.525 122.560 ;
        POLYGON 206.525 122.560 207.645 122.560 206.525 122.190 ;
        POLYGON 266.590 122.560 266.825 122.560 266.825 122.190 ;
        RECT 266.825 122.190 274.450 122.560 ;
        RECT 62.765 122.130 206.310 122.190 ;
        POLYGON 206.310 122.190 206.525 122.190 206.310 122.130 ;
        POLYGON 266.825 122.190 266.860 122.190 266.860 122.135 ;
        RECT 266.860 122.130 274.450 122.190 ;
        RECT 62.765 121.850 205.285 122.130 ;
        POLYGON 205.285 122.130 206.310 122.130 205.285 121.850 ;
        POLYGON 266.860 122.130 267.040 122.130 267.040 121.850 ;
        RECT 267.040 121.850 274.450 122.130 ;
        RECT 62.765 121.640 204.295 121.850 ;
        POLYGON 204.295 121.850 205.285 121.850 204.295 121.640 ;
        POLYGON 267.040 121.850 267.175 121.850 267.175 121.640 ;
        RECT 267.175 121.640 274.450 121.850 ;
        RECT 62.765 121.230 202.385 121.640 ;
        POLYGON 202.385 121.640 204.295 121.640 202.385 121.230 ;
        POLYGON 267.175 121.640 267.435 121.640 267.435 121.230 ;
        RECT 267.435 121.230 274.450 121.640 ;
        RECT 62.765 121.200 202.170 121.230 ;
        POLYGON 202.170 121.230 202.385 121.230 202.170 121.200 ;
        POLYGON 267.435 121.230 267.455 121.230 267.455 121.200 ;
        RECT 267.455 121.200 274.450 121.230 ;
        RECT 62.765 121.105 199.925 121.200 ;
        POLYGON 60.990 121.105 60.990 119.615 60.140 119.615 ;
        RECT 60.990 120.850 199.925 121.105 ;
        POLYGON 199.925 121.200 202.165 121.200 199.925 120.850 ;
        POLYGON 267.455 121.200 267.680 121.200 267.680 120.850 ;
        RECT 267.680 120.850 274.450 121.200 ;
        RECT 60.990 120.680 198.835 120.850 ;
        POLYGON 198.835 120.850 199.925 120.850 198.835 120.680 ;
        POLYGON 267.680 120.850 267.785 120.850 267.785 120.685 ;
        RECT 267.785 120.680 274.450 120.850 ;
        RECT 60.990 120.590 198.080 120.680 ;
        POLYGON 198.080 120.680 198.835 120.680 198.080 120.590 ;
        POLYGON 267.785 120.680 267.845 120.680 267.845 120.590 ;
        RECT 60.990 120.585 198.035 120.590 ;
        POLYGON 198.035 120.590 198.075 120.590 198.035 120.585 ;
        RECT 267.845 120.585 274.450 120.680 ;
        RECT 60.990 120.580 198.005 120.585 ;
        POLYGON 198.005 120.585 198.035 120.585 198.005 120.580 ;
        POLYGON 267.845 120.585 267.850 120.585 267.850 120.580 ;
        RECT 267.850 120.580 274.450 120.585 ;
        RECT 60.990 120.565 197.880 120.580 ;
        POLYGON 197.880 120.580 198.000 120.580 197.880 120.565 ;
        POLYGON 267.850 120.580 267.860 120.580 267.860 120.565 ;
        RECT 267.860 120.565 274.450 120.580 ;
        RECT 60.990 120.560 197.810 120.565 ;
        POLYGON 197.810 120.565 197.880 120.565 197.810 120.560 ;
        POLYGON 267.860 120.565 267.865 120.565 267.865 120.560 ;
        RECT 267.865 120.560 274.450 120.565 ;
        RECT 60.990 120.535 197.600 120.560 ;
        POLYGON 197.600 120.560 197.810 120.560 197.600 120.535 ;
        POLYGON 267.865 120.560 267.880 120.560 267.880 120.535 ;
        RECT 60.990 120.530 197.585 120.535 ;
        POLYGON 197.585 120.535 197.600 120.535 197.585 120.530 ;
        RECT 267.880 120.530 274.450 120.560 ;
        RECT 60.990 120.525 197.510 120.530 ;
        POLYGON 197.510 120.530 197.580 120.530 197.510 120.525 ;
        POLYGON 267.880 120.530 267.885 120.530 267.885 120.525 ;
        RECT 267.885 120.525 274.450 120.530 ;
        RECT 60.990 120.485 197.205 120.525 ;
        POLYGON 197.205 120.525 197.510 120.525 197.205 120.485 ;
        POLYGON 267.885 120.525 267.910 120.525 267.910 120.485 ;
        RECT 267.910 120.485 274.450 120.525 ;
        RECT 60.990 120.475 197.100 120.485 ;
        POLYGON 197.100 120.485 197.200 120.485 197.100 120.475 ;
        POLYGON 267.910 120.485 267.915 120.485 267.915 120.480 ;
        RECT 267.915 120.475 274.450 120.485 ;
        RECT 60.990 120.445 196.860 120.475 ;
        POLYGON 196.860 120.475 197.095 120.475 196.860 120.445 ;
        POLYGON 267.915 120.475 267.935 120.475 267.935 120.450 ;
        RECT 267.935 120.445 274.450 120.475 ;
        RECT 60.990 120.410 196.580 120.445 ;
        POLYGON 196.580 120.445 196.860 120.445 196.580 120.410 ;
        POLYGON 267.935 120.445 267.960 120.445 267.960 120.410 ;
        RECT 267.960 120.410 274.450 120.445 ;
        RECT 60.990 120.400 196.470 120.410 ;
        POLYGON 196.470 120.410 196.575 120.410 196.470 120.400 ;
        POLYGON 267.960 120.410 267.965 120.410 267.965 120.400 ;
        RECT 267.965 120.400 274.450 120.410 ;
        RECT 60.990 120.345 196.025 120.400 ;
        POLYGON 196.025 120.400 196.465 120.400 196.025 120.345 ;
        POLYGON 267.965 120.400 268.000 120.400 268.000 120.345 ;
        RECT 268.000 120.345 274.450 120.400 ;
        RECT 60.990 120.340 195.955 120.345 ;
        POLYGON 195.955 120.345 196.020 120.345 195.955 120.340 ;
        POLYGON 268.000 120.345 268.005 120.345 268.005 120.340 ;
        RECT 268.005 120.340 274.450 120.345 ;
        RECT 60.990 120.285 195.530 120.340 ;
        POLYGON 195.530 120.340 195.955 120.340 195.530 120.285 ;
        POLYGON 268.005 120.340 268.040 120.340 268.040 120.285 ;
        RECT 268.040 120.285 274.450 120.340 ;
        RECT 60.990 120.250 195.225 120.285 ;
        POLYGON 195.225 120.285 195.525 120.285 195.225 120.250 ;
        POLYGON 268.040 120.285 268.060 120.285 268.060 120.250 ;
        RECT 268.060 120.250 274.450 120.285 ;
        RECT 60.990 120.240 195.130 120.250 ;
        POLYGON 195.130 120.250 195.225 120.250 195.130 120.240 ;
        POLYGON 268.060 120.250 268.065 120.250 268.065 120.245 ;
        RECT 268.065 120.240 274.450 120.250 ;
        RECT 60.990 120.220 194.985 120.240 ;
        POLYGON 194.985 120.240 195.130 120.240 194.985 120.220 ;
        POLYGON 268.065 120.240 268.080 120.240 268.080 120.220 ;
        RECT 268.080 120.220 274.450 120.240 ;
        RECT 60.990 120.165 194.510 120.220 ;
        POLYGON 194.510 120.220 194.980 120.220 194.510 120.165 ;
        POLYGON 268.080 120.220 268.115 120.220 268.115 120.165 ;
        RECT 268.115 120.165 274.450 120.220 ;
        RECT 60.990 120.155 194.400 120.165 ;
        POLYGON 194.400 120.165 194.510 120.165 194.400 120.155 ;
        POLYGON 268.115 120.165 268.120 120.165 268.120 120.155 ;
        RECT 268.120 120.155 274.450 120.165 ;
        RECT 60.990 120.090 193.750 120.155 ;
        POLYGON 193.750 120.155 194.390 120.155 193.750 120.090 ;
        POLYGON 268.120 120.155 268.160 120.155 268.160 120.095 ;
        RECT 268.160 120.090 274.450 120.155 ;
        RECT 60.990 120.065 193.465 120.090 ;
        POLYGON 193.465 120.090 193.750 120.090 193.465 120.065 ;
        POLYGON 268.160 120.090 268.180 120.090 268.180 120.065 ;
        RECT 268.180 120.065 274.450 120.090 ;
        RECT 60.990 120.025 193.065 120.065 ;
        POLYGON 193.065 120.065 193.465 120.065 193.065 120.025 ;
        POLYGON 268.180 120.065 268.205 120.065 268.205 120.025 ;
        RECT 268.205 120.025 274.450 120.065 ;
        RECT 60.990 119.980 192.580 120.025 ;
        POLYGON 192.580 120.025 193.060 120.025 192.580 119.980 ;
        POLYGON 268.205 120.025 268.230 120.025 268.230 119.985 ;
        RECT 268.230 119.980 274.450 120.025 ;
        RECT 60.990 119.965 192.440 119.980 ;
        POLYGON 192.440 119.980 192.580 119.980 192.440 119.965 ;
        POLYGON 268.230 119.980 268.240 119.980 268.240 119.970 ;
        RECT 268.240 119.965 274.450 119.980 ;
        RECT 60.990 119.955 192.330 119.965 ;
        POLYGON 192.330 119.965 192.435 119.965 192.330 119.955 ;
        POLYGON 268.240 119.965 268.250 119.965 268.250 119.955 ;
        RECT 268.250 119.955 274.450 119.965 ;
        RECT 60.990 119.880 191.555 119.955 ;
        POLYGON 191.555 119.955 192.330 119.955 191.555 119.880 ;
        POLYGON 268.250 119.955 268.295 119.955 268.295 119.885 ;
        RECT 268.295 119.880 274.450 119.955 ;
        RECT 60.990 119.855 191.315 119.880 ;
        POLYGON 191.315 119.880 191.550 119.880 191.315 119.855 ;
        POLYGON 268.295 119.880 268.310 119.880 268.310 119.860 ;
        RECT 268.310 119.855 274.450 119.880 ;
        RECT 60.990 119.800 190.740 119.855 ;
        POLYGON 190.740 119.855 191.315 119.855 190.740 119.800 ;
        POLYGON 268.310 119.855 268.345 119.855 268.345 119.805 ;
        RECT 268.345 119.800 274.450 119.855 ;
        RECT 60.990 119.735 190.095 119.800 ;
        POLYGON 190.095 119.800 190.735 119.800 190.095 119.735 ;
        POLYGON 268.345 119.800 268.390 119.800 268.390 119.735 ;
        RECT 268.390 119.735 274.450 119.800 ;
        RECT 60.990 119.720 189.930 119.735 ;
        POLYGON 189.930 119.735 190.090 119.735 189.930 119.720 ;
        POLYGON 268.390 119.735 268.400 119.735 268.400 119.720 ;
        RECT 60.990 119.715 189.875 119.720 ;
        POLYGON 189.875 119.720 189.930 119.720 189.875 119.715 ;
        RECT 268.400 119.715 274.450 119.735 ;
        RECT 60.990 119.660 189.300 119.715 ;
        POLYGON 189.300 119.715 189.875 119.715 189.300 119.660 ;
        POLYGON 268.400 119.715 268.435 119.715 268.435 119.665 ;
        RECT 268.435 119.660 274.450 119.715 ;
        RECT 60.990 119.625 188.975 119.660 ;
        POLYGON 188.975 119.660 189.300 119.660 188.975 119.625 ;
        POLYGON 268.435 119.660 268.445 119.660 268.445 119.650 ;
        RECT 268.445 119.650 274.450 119.660 ;
        POLYGON 268.445 119.650 268.455 119.650 268.455 119.630 ;
        RECT 268.455 119.625 274.450 119.650 ;
        RECT 60.990 119.615 188.785 119.625 ;
        RECT 35.560 119.145 40.375 119.615 ;
        POLYGON 31.170 119.145 31.170 111.535 27.225 111.535 ;
        RECT 31.170 117.660 40.375 119.145 ;
        POLYGON 40.375 119.615 41.525 119.615 40.375 117.660 ;
        POLYGON 60.140 119.610 60.140 117.660 59.030 117.660 ;
        RECT 60.140 119.605 188.785 119.615 ;
        POLYGON 188.785 119.625 188.970 119.625 188.785 119.605 ;
        POLYGON 268.455 119.625 268.470 119.625 268.470 119.605 ;
        RECT 268.470 119.605 274.450 119.625 ;
        RECT 60.140 119.520 188.030 119.605 ;
        POLYGON 188.030 119.605 188.785 119.605 188.030 119.520 ;
        POLYGON 268.470 119.605 268.520 119.605 268.520 119.520 ;
        RECT 268.520 119.520 274.450 119.605 ;
        RECT 60.140 119.450 187.385 119.520 ;
        POLYGON 187.385 119.520 188.030 119.520 187.385 119.450 ;
        POLYGON 268.520 119.520 268.560 119.520 268.560 119.455 ;
        RECT 268.560 119.450 274.450 119.520 ;
        RECT 60.140 119.430 187.180 119.450 ;
        POLYGON 187.180 119.450 187.385 119.450 187.180 119.430 ;
        POLYGON 268.560 119.450 268.575 119.450 268.575 119.430 ;
        RECT 268.575 119.430 274.450 119.450 ;
        RECT 60.140 119.415 187.050 119.430 ;
        POLYGON 187.050 119.430 187.180 119.430 187.050 119.415 ;
        POLYGON 268.575 119.430 268.585 119.430 268.585 119.415 ;
        RECT 268.585 119.415 274.450 119.430 ;
        RECT 60.140 119.305 186.035 119.415 ;
        POLYGON 186.035 119.415 187.050 119.415 186.035 119.305 ;
        POLYGON 268.585 119.415 268.650 119.415 268.650 119.305 ;
        RECT 268.650 119.305 274.450 119.415 ;
        RECT 60.140 119.290 185.900 119.305 ;
        POLYGON 185.900 119.305 186.030 119.305 185.900 119.290 ;
        POLYGON 268.650 119.305 268.660 119.305 268.660 119.290 ;
        RECT 268.660 119.290 274.450 119.305 ;
        RECT 60.140 119.190 184.980 119.290 ;
        POLYGON 184.980 119.290 185.900 119.290 184.980 119.190 ;
        POLYGON 268.660 119.290 268.720 119.290 268.720 119.190 ;
        RECT 268.720 119.190 274.450 119.290 ;
        RECT 60.140 119.120 184.335 119.190 ;
        POLYGON 184.335 119.190 184.980 119.190 184.335 119.120 ;
        POLYGON 268.720 119.190 268.760 119.190 268.760 119.120 ;
        RECT 268.760 119.165 274.450 119.190 ;
        POLYGON 274.450 126.505 278.835 119.165 274.450 119.165 ;
        POLYGON 303.120 122.680 303.120 122.640 303.025 122.640 ;
        POLYGON 303.025 122.640 303.025 122.485 302.605 122.485 ;
        RECT 303.025 122.485 303.120 122.640 ;
        POLYGON 302.605 122.485 302.605 122.165 301.645 122.165 ;
        RECT 302.605 122.165 303.120 122.485 ;
        POLYGON 301.645 122.165 301.645 122.115 301.490 122.115 ;
        RECT 301.645 122.115 303.120 122.165 ;
        POLYGON 301.490 122.115 301.490 122.055 301.275 122.055 ;
        RECT 301.490 122.055 303.120 122.115 ;
        POLYGON 301.275 122.055 301.275 121.770 300.250 121.770 ;
        RECT 301.275 121.770 303.120 122.055 ;
        POLYGON 300.250 121.770 300.250 121.560 299.260 121.560 ;
        RECT 300.250 121.560 303.120 121.770 ;
        POLYGON 299.260 121.560 299.260 121.155 297.355 121.155 ;
        RECT 299.260 121.155 303.120 121.560 ;
        POLYGON 297.355 121.155 297.355 121.120 297.130 121.120 ;
        RECT 297.355 121.120 303.120 121.155 ;
        POLYGON 297.130 121.120 297.130 120.775 294.895 120.775 ;
        RECT 297.130 120.775 303.120 121.120 ;
        POLYGON 294.895 120.775 294.895 120.695 294.380 120.695 ;
        RECT 294.895 120.695 303.120 120.775 ;
        POLYGON 294.380 120.695 294.380 120.605 293.805 120.605 ;
        RECT 294.380 120.605 303.120 120.695 ;
        POLYGON 293.805 120.605 293.805 120.455 292.555 120.455 ;
        RECT 293.805 120.455 303.120 120.605 ;
        POLYGON 292.550 120.455 292.550 120.165 290.110 120.165 ;
        RECT 292.550 120.165 303.120 120.455 ;
        POLYGON 290.105 120.165 290.105 120.090 289.485 120.090 ;
        RECT 290.105 120.090 303.120 120.165 ;
        POLYGON 289.485 120.090 289.485 119.905 287.555 119.905 ;
        RECT 289.485 119.905 303.120 120.090 ;
        POLYGON 287.555 119.905 287.555 119.845 286.945 119.845 ;
        RECT 287.555 119.845 303.120 119.905 ;
        POLYGON 286.940 119.845 286.940 119.645 284.905 119.645 ;
        RECT 286.940 119.645 303.120 119.845 ;
        POLYGON 284.905 119.645 284.905 119.585 284.280 119.585 ;
        RECT 284.905 119.585 303.120 119.645 ;
        POLYGON 284.280 119.585 284.280 119.365 282.160 119.365 ;
        RECT 284.280 119.365 303.120 119.585 ;
        POLYGON 282.155 119.365 282.155 119.165 280.260 119.165 ;
        RECT 282.155 119.165 303.120 119.365 ;
        RECT 268.760 119.120 278.835 119.165 ;
        RECT 60.140 119.070 183.890 119.120 ;
        POLYGON 183.890 119.120 184.325 119.120 183.890 119.070 ;
        POLYGON 268.760 119.120 268.790 119.120 268.790 119.070 ;
        RECT 268.790 119.070 278.835 119.120 ;
        POLYGON 278.835 119.165 278.885 119.070 278.835 119.070 ;
        POLYGON 280.260 119.165 280.260 119.070 279.360 119.070 ;
        RECT 280.260 119.070 303.120 119.165 ;
        RECT 60.140 118.950 182.765 119.070 ;
        POLYGON 182.765 119.070 183.890 119.070 182.765 118.950 ;
        POLYGON 268.790 119.070 268.860 119.070 268.860 118.955 ;
        RECT 268.860 119.040 278.885 119.070 ;
        POLYGON 278.885 119.070 278.900 119.040 278.885 119.040 ;
        POLYGON 279.320 119.070 279.320 119.040 279.045 119.040 ;
        RECT 279.320 119.040 303.120 119.070 ;
        RECT 268.860 119.025 278.900 119.040 ;
        POLYGON 278.900 119.040 278.910 119.025 278.900 119.025 ;
        POLYGON 279.030 119.040 279.030 119.025 278.910 119.025 ;
        RECT 279.030 119.025 303.120 119.040 ;
        RECT 268.860 118.950 303.120 119.025 ;
        RECT 60.140 118.940 182.665 118.950 ;
        POLYGON 182.665 118.950 182.765 118.950 182.665 118.940 ;
        POLYGON 268.860 118.950 268.865 118.950 268.865 118.945 ;
        RECT 268.865 118.940 303.120 118.950 ;
        RECT 60.140 118.825 181.610 118.940 ;
        POLYGON 181.610 118.940 182.665 118.940 181.610 118.825 ;
        POLYGON 268.865 118.940 268.935 118.940 268.935 118.830 ;
        RECT 268.935 118.825 303.120 118.940 ;
        RECT 60.140 118.800 181.400 118.825 ;
        POLYGON 181.400 118.825 181.605 118.825 181.400 118.800 ;
        POLYGON 268.935 118.825 268.950 118.825 268.950 118.805 ;
        RECT 268.950 118.800 303.120 118.825 ;
        RECT 60.140 118.750 180.925 118.800 ;
        POLYGON 180.925 118.800 181.400 118.800 180.925 118.750 ;
        POLYGON 268.950 118.800 268.980 118.800 268.980 118.755 ;
        RECT 268.980 118.750 303.120 118.800 ;
        RECT 60.140 118.695 180.420 118.750 ;
        POLYGON 180.420 118.750 180.925 118.750 180.420 118.695 ;
        POLYGON 268.980 118.750 269.015 118.750 269.015 118.695 ;
        RECT 269.015 118.695 303.120 118.750 ;
        RECT 60.140 118.565 179.200 118.695 ;
        POLYGON 179.200 118.695 180.415 118.695 179.200 118.565 ;
        POLYGON 269.015 118.695 269.090 118.695 269.090 118.570 ;
        RECT 269.090 118.565 303.120 118.695 ;
        RECT 60.140 118.555 179.105 118.565 ;
        POLYGON 179.105 118.565 179.200 118.565 179.105 118.555 ;
        POLYGON 269.090 118.565 269.100 118.565 269.100 118.555 ;
        RECT 269.100 118.555 303.120 118.565 ;
        RECT 60.140 118.475 178.370 118.555 ;
        POLYGON 178.370 118.555 179.105 118.555 178.370 118.475 ;
        POLYGON 269.100 118.555 269.145 118.555 269.145 118.480 ;
        RECT 269.145 118.475 303.120 118.555 ;
        RECT 60.140 118.425 177.945 118.475 ;
        POLYGON 177.945 118.475 178.370 118.475 177.945 118.425 ;
        POLYGON 269.145 118.475 269.175 118.475 269.175 118.430 ;
        RECT 269.175 118.425 303.120 118.475 ;
        RECT 60.140 118.345 177.210 118.425 ;
        POLYGON 177.210 118.425 177.945 118.425 177.210 118.345 ;
        POLYGON 269.175 118.425 269.225 118.425 269.225 118.345 ;
        RECT 269.225 118.345 303.120 118.425 ;
        RECT 60.140 118.290 176.670 118.345 ;
        POLYGON 176.670 118.345 177.210 118.345 176.670 118.290 ;
        POLYGON 269.225 118.345 269.255 118.345 269.255 118.295 ;
        RECT 269.255 118.290 303.120 118.345 ;
        RECT 60.140 118.260 176.415 118.290 ;
        POLYGON 176.415 118.290 176.665 118.290 176.415 118.260 ;
        POLYGON 269.255 118.290 269.275 118.290 269.275 118.260 ;
        RECT 269.275 118.260 303.120 118.290 ;
        RECT 60.140 118.080 175.360 118.260 ;
        POLYGON 175.360 118.260 176.415 118.260 175.360 118.080 ;
        POLYGON 269.275 118.260 269.380 118.260 269.380 118.085 ;
        RECT 269.380 118.080 303.120 118.260 ;
        RECT 60.140 118.065 175.260 118.080 ;
        POLYGON 175.260 118.080 175.360 118.080 175.260 118.065 ;
        POLYGON 269.380 118.080 269.390 118.080 269.390 118.070 ;
        RECT 269.390 118.065 303.120 118.080 ;
        RECT 60.140 118.060 175.235 118.065 ;
        POLYGON 175.235 118.065 175.255 118.065 175.235 118.060 ;
        POLYGON 269.390 118.065 269.395 118.065 269.395 118.060 ;
        RECT 269.395 118.060 303.120 118.065 ;
        RECT 60.140 117.855 174.030 118.060 ;
        POLYGON 174.030 118.060 175.235 118.060 174.030 117.855 ;
        POLYGON 269.395 118.060 269.445 118.060 269.445 117.980 ;
        RECT 269.445 117.980 303.120 118.060 ;
        POLYGON 269.445 117.980 269.510 117.980 269.510 117.870 ;
        RECT 269.510 117.870 303.120 117.980 ;
        POLYGON 269.500 117.870 269.500 117.860 269.445 117.860 ;
        RECT 269.500 117.860 303.120 117.870 ;
        POLYGON 269.430 117.860 269.430 117.855 269.395 117.855 ;
        RECT 269.430 117.855 303.120 117.860 ;
        RECT 60.140 117.715 173.185 117.855 ;
        POLYGON 173.185 117.855 174.025 117.855 173.185 117.715 ;
        POLYGON 269.395 117.855 269.395 117.720 268.480 117.720 ;
        RECT 269.395 117.720 303.120 117.855 ;
        POLYGON 268.480 117.720 268.480 117.715 268.445 117.715 ;
        RECT 268.480 117.715 303.120 117.720 ;
        RECT 60.140 117.660 172.670 117.715 ;
        RECT 31.170 114.715 38.655 117.660 ;
        POLYGON 38.655 117.660 40.375 117.660 38.655 114.715 ;
        POLYGON 59.030 117.660 59.030 117.380 58.870 117.380 ;
        RECT 59.030 117.625 172.670 117.660 ;
        POLYGON 172.670 117.715 173.185 117.715 172.670 117.625 ;
        POLYGON 268.445 117.715 268.445 117.625 267.835 117.625 ;
        RECT 268.445 117.625 303.120 117.715 ;
        RECT 59.030 117.525 172.055 117.625 ;
        POLYGON 172.055 117.625 172.665 117.625 172.055 117.525 ;
        POLYGON 267.835 117.625 267.835 117.525 267.155 117.525 ;
        RECT 267.835 117.525 303.120 117.625 ;
        RECT 59.030 117.390 171.285 117.525 ;
        POLYGON 171.285 117.525 172.055 117.525 171.285 117.390 ;
        POLYGON 267.155 117.525 267.155 117.510 267.055 117.510 ;
        RECT 267.155 117.510 303.120 117.525 ;
        POLYGON 267.050 117.510 267.050 117.390 266.240 117.390 ;
        RECT 267.050 117.390 303.120 117.510 ;
        RECT 59.030 117.380 171.070 117.390 ;
        POLYGON 58.870 117.380 58.870 117.155 58.745 117.155 ;
        RECT 58.870 117.355 171.070 117.380 ;
        POLYGON 171.070 117.390 171.280 117.390 171.070 117.355 ;
        POLYGON 266.240 117.390 266.240 117.360 266.035 117.360 ;
        RECT 266.240 117.360 303.120 117.390 ;
        POLYGON 266.035 117.360 266.035 117.355 266.000 117.355 ;
        RECT 266.035 117.355 303.120 117.360 ;
        RECT 58.870 117.155 169.875 117.355 ;
        POLYGON 169.875 117.355 171.065 117.355 169.875 117.155 ;
        POLYGON 266.000 117.355 266.000 117.195 264.920 117.195 ;
        RECT 266.000 117.195 303.120 117.355 ;
        POLYGON 264.920 117.195 264.920 117.160 264.740 117.160 ;
        RECT 264.920 117.160 303.120 117.195 ;
        POLYGON 264.740 117.160 264.740 117.155 264.715 117.155 ;
        RECT 264.740 117.155 303.120 117.160 ;
        POLYGON 58.745 117.155 58.745 114.715 57.510 114.715 ;
        RECT 58.745 116.985 168.875 117.155 ;
        POLYGON 168.875 117.155 169.875 117.155 168.875 116.985 ;
        POLYGON 264.715 117.155 264.715 116.990 263.865 116.990 ;
        RECT 264.715 116.990 303.120 117.155 ;
        POLYGON 263.865 116.990 263.865 116.985 263.840 116.985 ;
        RECT 263.865 116.985 303.120 116.990 ;
        RECT 58.745 116.970 168.775 116.985 ;
        POLYGON 168.775 116.985 168.875 116.985 168.775 116.970 ;
        POLYGON 263.840 116.985 263.840 116.975 263.790 116.975 ;
        RECT 263.840 116.975 303.120 116.985 ;
        POLYGON 263.785 116.975 263.785 116.970 263.770 116.970 ;
        RECT 263.785 116.970 303.120 116.975 ;
        RECT 58.745 116.910 168.445 116.970 ;
        POLYGON 168.445 116.970 168.770 116.970 168.445 116.910 ;
        POLYGON 263.770 116.970 263.770 116.915 263.490 116.915 ;
        RECT 263.770 116.915 303.120 116.970 ;
        POLYGON 263.490 116.915 263.490 116.910 263.465 116.910 ;
        RECT 263.490 116.910 303.120 116.915 ;
        RECT 58.745 116.665 166.995 116.910 ;
        POLYGON 166.995 116.910 168.445 116.910 166.995 116.665 ;
        POLYGON 263.465 116.910 263.465 116.665 262.215 116.665 ;
        RECT 263.465 116.665 303.120 116.910 ;
        RECT 58.745 116.605 166.620 116.665 ;
        POLYGON 166.620 116.665 166.995 116.665 166.620 116.605 ;
        POLYGON 262.215 116.665 262.215 116.605 261.910 116.605 ;
        RECT 262.215 116.605 303.120 116.665 ;
        RECT 58.745 116.535 166.205 116.605 ;
        POLYGON 166.205 116.605 166.615 116.605 166.205 116.535 ;
        POLYGON 261.910 116.605 261.910 116.540 261.580 116.540 ;
        RECT 261.910 116.540 303.120 116.605 ;
        POLYGON 261.580 116.540 261.580 116.535 261.550 116.535 ;
        RECT 261.580 116.535 303.120 116.540 ;
        RECT 58.745 116.370 165.525 116.535 ;
        POLYGON 165.525 116.535 166.205 116.535 165.525 116.370 ;
        POLYGON 261.550 116.535 261.550 116.460 261.170 116.460 ;
        RECT 261.550 116.460 303.120 116.535 ;
        POLYGON 261.170 116.460 261.170 116.370 260.790 116.370 ;
        RECT 261.170 116.370 303.120 116.460 ;
        RECT 58.745 116.345 165.410 116.370 ;
        POLYGON 165.410 116.370 165.525 116.370 165.410 116.345 ;
        POLYGON 260.790 116.370 260.790 116.345 260.685 116.345 ;
        RECT 260.790 116.345 303.120 116.370 ;
        RECT 58.745 116.075 164.290 116.345 ;
        POLYGON 164.290 116.345 165.405 116.345 164.290 116.075 ;
        POLYGON 260.685 116.345 260.685 116.280 260.410 116.280 ;
        RECT 260.685 116.280 303.120 116.345 ;
        POLYGON 260.410 116.280 260.410 116.080 259.565 116.080 ;
        RECT 260.410 116.080 303.120 116.280 ;
        POLYGON 259.565 116.080 259.565 116.075 259.545 116.075 ;
        RECT 259.565 116.075 303.120 116.080 ;
        RECT 58.745 116.040 164.145 116.075 ;
        POLYGON 164.145 116.075 164.290 116.075 164.145 116.040 ;
        POLYGON 259.545 116.075 259.545 116.040 259.395 116.040 ;
        RECT 259.545 116.040 303.120 116.075 ;
        RECT 58.745 115.665 162.565 116.040 ;
        POLYGON 162.565 116.040 164.145 116.040 162.565 115.665 ;
        POLYGON 259.395 116.040 259.395 115.840 258.550 115.840 ;
        RECT 259.395 115.840 303.120 116.040 ;
        POLYGON 258.550 115.840 258.550 115.665 257.810 115.665 ;
        RECT 258.550 115.665 303.120 115.840 ;
        RECT 58.745 115.520 161.965 115.665 ;
        POLYGON 161.965 115.665 162.565 115.665 161.965 115.520 ;
        POLYGON 257.810 115.665 257.810 115.630 257.660 115.630 ;
        RECT 257.810 115.630 303.120 115.665 ;
        POLYGON 257.660 115.630 257.660 115.520 257.260 115.520 ;
        RECT 257.660 115.520 303.120 115.630 ;
        RECT 58.745 115.515 161.945 115.520 ;
        POLYGON 161.945 115.520 161.965 115.520 161.945 115.515 ;
        POLYGON 257.260 115.520 257.260 115.515 257.240 115.515 ;
        RECT 257.260 115.515 303.120 115.520 ;
        RECT 58.745 115.505 161.890 115.515 ;
        POLYGON 161.890 115.515 161.945 115.515 161.890 115.505 ;
        POLYGON 257.240 115.515 257.240 115.505 257.205 115.505 ;
        RECT 257.240 115.505 303.120 115.515 ;
        RECT 58.745 115.465 161.735 115.505 ;
        POLYGON 161.735 115.505 161.890 115.505 161.735 115.465 ;
        POLYGON 257.205 115.505 257.205 115.465 257.060 115.465 ;
        RECT 257.205 115.465 303.120 115.505 ;
        RECT 58.745 115.210 160.850 115.465 ;
        POLYGON 160.850 115.465 161.735 115.465 160.850 115.210 ;
        POLYGON 257.060 115.465 257.060 115.440 256.970 115.440 ;
        RECT 257.060 115.440 303.120 115.465 ;
        POLYGON 256.970 115.440 256.970 115.215 256.155 115.215 ;
        RECT 256.970 115.215 303.120 115.440 ;
        POLYGON 256.155 115.215 256.155 115.210 256.135 115.210 ;
        RECT 256.155 115.210 303.120 115.215 ;
        RECT 58.745 114.790 159.430 115.210 ;
        POLYGON 159.430 115.210 160.850 115.210 159.430 114.790 ;
        POLYGON 256.135 115.210 256.135 115.130 255.845 115.130 ;
        RECT 256.135 115.130 303.120 115.210 ;
        POLYGON 255.840 115.130 255.840 114.790 254.615 114.790 ;
        RECT 255.840 114.790 303.120 115.130 ;
        RECT 58.745 114.715 157.495 114.790 ;
        RECT 31.170 111.535 36.040 114.715 ;
        POLYGON 27.225 111.535 27.225 103.685 23.730 103.685 ;
        RECT 27.225 109.770 36.040 111.535 ;
        POLYGON 36.040 114.715 38.655 114.715 36.040 109.770 ;
        POLYGON 57.510 114.715 57.510 114.200 57.250 114.200 ;
        RECT 57.510 114.225 157.495 114.715 ;
        POLYGON 157.495 114.790 159.430 114.790 157.495 114.225 ;
        POLYGON 254.615 114.790 254.615 114.700 254.290 114.700 ;
        RECT 254.615 114.700 303.120 114.790 ;
        POLYGON 254.290 114.700 254.290 114.230 252.820 114.230 ;
        RECT 254.290 114.230 303.120 114.700 ;
        POLYGON 252.820 114.230 252.820 114.225 252.805 114.225 ;
        RECT 252.820 114.225 303.120 114.230 ;
        RECT 57.510 114.200 157.305 114.225 ;
        POLYGON 57.250 114.200 57.250 113.150 56.720 113.150 ;
        RECT 57.250 114.160 157.305 114.200 ;
        POLYGON 157.305 114.225 157.495 114.225 157.305 114.160 ;
        POLYGON 252.805 114.225 252.805 114.160 252.600 114.160 ;
        RECT 252.805 114.160 303.120 114.225 ;
        RECT 57.250 114.105 157.145 114.160 ;
        POLYGON 157.145 114.160 157.305 114.160 157.145 114.105 ;
        POLYGON 252.600 114.160 252.600 114.105 252.430 114.105 ;
        RECT 252.600 114.105 303.120 114.160 ;
        RECT 57.250 113.835 156.375 114.105 ;
        POLYGON 156.375 114.105 157.145 114.105 156.375 113.835 ;
        POLYGON 252.430 114.105 252.430 113.835 251.585 113.835 ;
        RECT 252.430 113.835 303.120 114.105 ;
        RECT 57.250 113.570 155.615 113.835 ;
        POLYGON 155.615 113.835 156.370 113.835 155.615 113.570 ;
        POLYGON 251.585 113.835 251.585 113.640 250.970 113.640 ;
        RECT 251.585 113.640 303.120 113.835 ;
        POLYGON 250.970 113.640 250.970 113.625 250.935 113.625 ;
        RECT 250.970 113.625 303.120 113.640 ;
        POLYGON 250.935 113.625 250.935 113.570 250.785 113.570 ;
        RECT 250.935 113.570 303.120 113.625 ;
        RECT 57.250 113.290 154.815 113.570 ;
        POLYGON 154.815 113.570 155.615 113.570 154.815 113.290 ;
        POLYGON 250.785 113.570 250.785 113.290 250.020 113.290 ;
        RECT 250.785 113.290 303.120 113.570 ;
        RECT 57.250 113.150 154.070 113.290 ;
        POLYGON 56.720 113.150 56.720 109.770 55.215 109.770 ;
        RECT 56.720 113.030 154.070 113.150 ;
        POLYGON 154.070 113.290 154.815 113.290 154.070 113.030 ;
        POLYGON 250.020 113.290 250.020 113.030 249.310 113.030 ;
        RECT 250.020 113.030 303.120 113.290 ;
        RECT 56.720 112.775 153.340 113.030 ;
        POLYGON 153.340 113.030 154.070 113.030 153.340 112.775 ;
        POLYGON 249.310 113.030 249.310 112.775 248.610 112.775 ;
        RECT 249.310 112.775 303.120 113.030 ;
        RECT 56.720 112.600 152.895 112.775 ;
        POLYGON 152.895 112.775 153.340 112.775 152.895 112.600 ;
        POLYGON 248.610 112.775 248.610 112.600 248.130 112.600 ;
        RECT 248.610 112.600 303.120 112.775 ;
        RECT 56.720 112.540 152.745 112.600 ;
        POLYGON 152.745 112.600 152.895 112.600 152.745 112.540 ;
        POLYGON 248.130 112.600 248.130 112.540 247.970 112.540 ;
        RECT 248.130 112.540 303.120 112.600 ;
        RECT 56.720 112.425 152.465 112.540 ;
        POLYGON 152.465 112.540 152.745 112.540 152.465 112.425 ;
        POLYGON 247.970 112.540 247.970 112.425 247.655 112.425 ;
        RECT 247.970 112.425 303.120 112.540 ;
        RECT 56.720 112.405 152.415 112.425 ;
        POLYGON 152.415 112.425 152.465 112.425 152.415 112.405 ;
        POLYGON 247.655 112.425 247.655 112.405 247.600 112.405 ;
        RECT 247.655 112.405 303.120 112.425 ;
        RECT 56.720 112.060 151.550 112.405 ;
        POLYGON 151.550 112.405 152.415 112.405 151.550 112.060 ;
        POLYGON 247.600 112.405 247.600 112.230 247.120 112.230 ;
        RECT 247.600 112.230 303.120 112.405 ;
        POLYGON 247.120 112.230 247.120 112.075 246.755 112.075 ;
        RECT 247.120 112.075 303.120 112.230 ;
        POLYGON 246.755 112.075 246.755 112.065 246.730 112.065 ;
        RECT 246.755 112.065 303.120 112.075 ;
        POLYGON 246.730 112.065 246.730 112.060 246.720 112.060 ;
        RECT 246.730 112.060 303.120 112.065 ;
        RECT 56.720 111.995 151.390 112.060 ;
        POLYGON 151.390 112.060 151.550 112.060 151.390 111.995 ;
        POLYGON 246.720 112.060 246.720 111.995 246.565 111.995 ;
        RECT 246.720 111.995 303.120 112.060 ;
        RECT 56.720 111.985 151.360 111.995 ;
        POLYGON 151.360 111.995 151.390 111.995 151.360 111.985 ;
        POLYGON 246.565 111.995 246.565 111.985 246.540 111.985 ;
        RECT 246.565 111.985 303.120 111.995 ;
        RECT 56.720 111.980 151.355 111.985 ;
        RECT 56.720 111.970 151.350 111.980 ;
        POLYGON 151.350 111.980 151.355 111.980 151.350 111.975 ;
        POLYGON 246.540 111.985 246.540 111.975 246.515 111.975 ;
        RECT 246.540 111.975 303.120 111.985 ;
        POLYGON 246.515 111.975 246.515 111.970 246.505 111.970 ;
        RECT 246.515 111.970 303.120 111.975 ;
        RECT 56.720 111.920 151.325 111.970 ;
        POLYGON 151.325 111.970 151.350 111.970 151.325 111.925 ;
        POLYGON 246.505 111.970 246.505 111.925 246.400 111.925 ;
        RECT 246.505 111.925 303.120 111.970 ;
        POLYGON 246.400 111.925 246.400 111.920 246.385 111.920 ;
        RECT 246.400 111.920 303.120 111.925 ;
        RECT 56.720 111.660 151.200 111.920 ;
        POLYGON 151.200 111.920 151.325 111.920 151.200 111.660 ;
        POLYGON 246.385 111.920 246.385 111.780 246.055 111.780 ;
        RECT 246.385 111.780 303.120 111.920 ;
        POLYGON 246.055 111.780 246.055 111.660 245.770 111.660 ;
        RECT 246.055 111.660 303.120 111.780 ;
        RECT 56.720 111.595 151.170 111.660 ;
        POLYGON 151.170 111.660 151.200 111.660 151.170 111.600 ;
        POLYGON 245.770 111.660 245.770 111.600 245.630 111.600 ;
        RECT 245.770 111.600 303.120 111.660 ;
        POLYGON 245.630 111.600 245.630 111.595 245.620 111.595 ;
        RECT 245.630 111.595 303.120 111.600 ;
        RECT 56.720 111.480 151.115 111.595 ;
        POLYGON 151.115 111.595 151.170 111.595 151.115 111.485 ;
        POLYGON 245.620 111.595 245.620 111.485 245.360 111.485 ;
        RECT 245.620 111.485 303.120 111.595 ;
        RECT 56.720 111.130 150.950 111.480 ;
        POLYGON 150.950 111.480 151.115 111.480 150.950 111.135 ;
        POLYGON 245.360 111.485 245.360 111.135 244.535 111.135 ;
        RECT 245.360 111.135 303.120 111.485 ;
        RECT 56.720 111.095 150.935 111.130 ;
        POLYGON 150.935 111.130 150.950 111.130 150.935 111.100 ;
        POLYGON 244.535 111.135 244.535 111.100 244.450 111.100 ;
        RECT 244.535 111.100 303.120 111.135 ;
        POLYGON 244.450 111.100 244.450 111.095 244.440 111.095 ;
        RECT 244.450 111.095 303.120 111.100 ;
        RECT 56.720 110.625 150.715 111.095 ;
        POLYGON 150.715 111.095 150.935 111.095 150.715 110.630 ;
        POLYGON 244.440 111.095 244.440 110.995 244.205 110.995 ;
        RECT 244.440 110.995 303.120 111.095 ;
        POLYGON 244.205 110.995 244.205 110.660 243.405 110.660 ;
        RECT 244.205 110.660 303.120 110.995 ;
        POLYGON 243.405 110.660 243.405 110.630 243.345 110.630 ;
        RECT 243.405 110.630 303.120 110.660 ;
        POLYGON 243.345 110.630 243.345 110.625 243.335 110.625 ;
        RECT 243.345 110.625 303.120 110.630 ;
        RECT 56.720 110.450 150.630 110.625 ;
        POLYGON 150.630 110.625 150.715 110.625 150.630 110.450 ;
        POLYGON 243.335 110.625 243.335 110.450 242.970 110.450 ;
        RECT 243.335 110.450 303.120 110.625 ;
        RECT 56.720 110.290 150.555 110.450 ;
        POLYGON 150.555 110.450 150.630 110.450 150.555 110.290 ;
        POLYGON 242.970 110.450 242.970 110.290 242.640 110.290 ;
        RECT 242.970 110.290 303.120 110.450 ;
        RECT 56.720 110.125 150.490 110.290 ;
        POLYGON 150.490 110.290 150.555 110.290 150.490 110.125 ;
        POLYGON 242.640 110.290 242.640 110.125 242.300 110.125 ;
        RECT 242.640 110.125 303.120 110.290 ;
        RECT 56.720 109.770 150.315 110.125 ;
        RECT 27.225 108.755 35.560 109.770 ;
        POLYGON 35.560 109.770 36.040 109.770 35.560 108.755 ;
        POLYGON 55.215 109.770 55.215 109.480 55.085 109.480 ;
        RECT 55.215 109.685 150.315 109.770 ;
        POLYGON 150.315 110.125 150.490 110.125 150.315 109.685 ;
        POLYGON 242.300 110.125 242.300 109.685 241.390 109.685 ;
        RECT 242.300 109.685 303.120 110.125 ;
        RECT 55.215 109.635 150.295 109.685 ;
        POLYGON 150.295 109.685 150.315 109.685 150.295 109.635 ;
        POLYGON 241.390 109.685 241.390 109.635 241.290 109.635 ;
        RECT 241.390 109.635 303.120 109.685 ;
        RECT 55.215 109.480 150.170 109.635 ;
        POLYGON 55.085 109.480 55.085 109.090 54.910 109.090 ;
        RECT 55.085 109.320 150.170 109.480 ;
        POLYGON 150.170 109.635 150.295 109.635 150.170 109.320 ;
        POLYGON 241.290 109.635 241.290 109.595 241.205 109.595 ;
        RECT 241.290 109.595 303.120 109.635 ;
        POLYGON 241.205 109.595 241.205 109.320 240.635 109.320 ;
        RECT 241.205 109.320 303.120 109.595 ;
        RECT 55.085 109.090 150.075 109.320 ;
        POLYGON 54.910 109.090 54.910 108.755 54.780 108.755 ;
        RECT 54.910 109.080 150.075 109.090 ;
        POLYGON 150.075 109.320 150.170 109.320 150.075 109.080 ;
        POLYGON 240.635 109.320 240.635 109.080 240.135 109.080 ;
        RECT 240.635 109.080 303.120 109.320 ;
        RECT 54.910 108.865 149.990 109.080 ;
        POLYGON 149.990 109.080 150.075 109.080 149.990 108.865 ;
        POLYGON 240.135 109.080 240.135 108.935 239.835 108.935 ;
        RECT 240.135 108.935 303.120 109.080 ;
        POLYGON 239.835 108.935 239.835 108.865 239.710 108.865 ;
        RECT 239.835 108.865 303.120 108.935 ;
        RECT 54.910 108.755 149.930 108.865 ;
        RECT 27.225 104.440 33.520 108.755 ;
        POLYGON 33.520 108.755 35.560 108.755 33.520 104.440 ;
        POLYGON 54.780 108.755 54.780 104.985 53.325 104.985 ;
        RECT 54.780 108.715 149.930 108.755 ;
        POLYGON 149.930 108.865 149.990 108.865 149.930 108.715 ;
        POLYGON 239.710 108.865 239.710 108.715 239.435 108.715 ;
        RECT 239.710 108.715 303.120 108.865 ;
        RECT 54.780 108.545 149.865 108.715 ;
        POLYGON 149.865 108.715 149.930 108.715 149.865 108.550 ;
        POLYGON 239.435 108.715 239.435 108.550 239.135 108.550 ;
        RECT 239.435 108.550 303.120 108.715 ;
        POLYGON 239.135 108.550 239.135 108.545 239.125 108.545 ;
        RECT 239.135 108.545 303.120 108.550 ;
        RECT 54.780 108.310 149.770 108.545 ;
        POLYGON 149.770 108.545 149.865 108.545 149.770 108.310 ;
        POLYGON 239.125 108.545 239.125 108.310 238.695 108.310 ;
        RECT 239.125 108.310 303.120 108.545 ;
        RECT 54.780 108.135 149.700 108.310 ;
        POLYGON 149.700 108.310 149.770 108.310 149.700 108.135 ;
        POLYGON 238.695 108.310 238.695 108.135 238.380 108.135 ;
        RECT 238.695 108.135 303.120 108.310 ;
        RECT 54.780 108.070 149.675 108.135 ;
        POLYGON 149.675 108.135 149.700 108.135 149.675 108.070 ;
        POLYGON 238.380 108.135 238.380 108.070 238.260 108.070 ;
        RECT 238.380 108.070 303.120 108.135 ;
        RECT 54.780 108.010 149.650 108.070 ;
        POLYGON 149.650 108.070 149.675 108.070 149.650 108.015 ;
        POLYGON 238.260 108.070 238.260 108.015 238.160 108.015 ;
        RECT 238.260 108.015 303.120 108.070 ;
        RECT 54.780 107.545 149.465 108.010 ;
        POLYGON 149.465 108.010 149.650 108.010 149.465 107.545 ;
        POLYGON 238.160 108.015 238.160 107.545 237.305 107.545 ;
        RECT 238.160 107.545 303.120 108.015 ;
        RECT 54.780 107.430 149.420 107.545 ;
        POLYGON 149.420 107.545 149.465 107.545 149.420 107.435 ;
        POLYGON 237.305 107.545 237.305 107.435 237.105 107.435 ;
        RECT 237.305 107.435 303.120 107.545 ;
        RECT 54.780 106.875 149.200 107.430 ;
        POLYGON 149.200 107.430 149.420 107.430 149.200 106.875 ;
        POLYGON 237.105 107.435 237.105 107.395 237.030 107.395 ;
        RECT 237.105 107.395 303.120 107.435 ;
        POLYGON 237.025 107.395 237.025 107.060 236.410 107.060 ;
        RECT 237.025 107.060 303.120 107.395 ;
        POLYGON 236.410 107.060 236.410 107.045 236.385 107.045 ;
        RECT 236.410 107.045 303.120 107.060 ;
        POLYGON 236.385 107.045 236.385 106.875 236.110 106.875 ;
        RECT 236.385 106.875 303.120 107.045 ;
        RECT 54.780 106.670 149.120 106.875 ;
        POLYGON 149.120 106.875 149.200 106.875 149.120 106.675 ;
        POLYGON 236.110 106.875 236.110 106.675 235.790 106.675 ;
        RECT 236.110 106.675 303.120 106.875 ;
        POLYGON 235.790 106.675 235.790 106.670 235.780 106.670 ;
        RECT 235.790 106.670 303.120 106.675 ;
        RECT 54.780 106.435 149.025 106.670 ;
        POLYGON 149.025 106.670 149.120 106.670 149.025 106.435 ;
        POLYGON 235.780 106.670 235.780 106.435 235.400 106.435 ;
        RECT 235.780 106.435 303.120 106.670 ;
        RECT 54.780 106.315 148.980 106.435 ;
        POLYGON 148.980 106.435 149.025 106.435 148.980 106.320 ;
        POLYGON 235.400 106.435 235.400 106.320 235.215 106.320 ;
        RECT 235.400 106.320 303.120 106.435 ;
        POLYGON 235.215 106.320 235.215 106.315 235.205 106.315 ;
        RECT 235.215 106.315 303.120 106.320 ;
        RECT 54.780 105.725 148.745 106.315 ;
        POLYGON 148.745 106.315 148.980 106.315 148.745 105.730 ;
        POLYGON 235.205 106.315 235.205 105.730 234.260 105.730 ;
        RECT 235.205 105.730 303.120 106.315 ;
        POLYGON 234.260 105.730 234.260 105.725 234.255 105.725 ;
        RECT 234.260 105.725 303.120 105.730 ;
        RECT 54.780 105.225 148.545 105.725 ;
        POLYGON 148.545 105.725 148.745 105.725 148.545 105.225 ;
        POLYGON 234.255 105.725 234.255 105.225 233.445 105.225 ;
        RECT 234.255 105.225 303.120 105.725 ;
        RECT 54.780 105.140 148.515 105.225 ;
        POLYGON 148.515 105.225 148.545 105.225 148.515 105.145 ;
        POLYGON 233.445 105.225 233.445 105.145 233.320 105.145 ;
        RECT 233.445 105.145 303.120 105.225 ;
        RECT 54.780 105.110 148.505 105.140 ;
        POLYGON 148.505 105.140 148.515 105.140 148.505 105.110 ;
        POLYGON 233.320 105.145 233.320 105.110 233.260 105.110 ;
        RECT 233.320 105.110 303.120 105.145 ;
        RECT 54.780 104.985 148.330 105.110 ;
        POLYGON 53.325 104.985 53.325 104.440 53.145 104.440 ;
        RECT 53.325 104.600 148.330 104.985 ;
        POLYGON 148.330 105.110 148.505 105.110 148.330 104.605 ;
        POLYGON 233.260 105.110 233.260 105.035 233.140 105.035 ;
        RECT 233.260 105.035 303.120 105.110 ;
        POLYGON 233.140 105.035 233.140 104.605 232.520 104.605 ;
        RECT 233.140 104.605 303.120 105.035 ;
        RECT 53.325 104.585 148.325 104.600 ;
        POLYGON 148.325 104.600 148.330 104.600 148.325 104.585 ;
        POLYGON 232.520 104.605 232.520 104.585 232.490 104.585 ;
        RECT 232.520 104.585 303.120 104.605 ;
        RECT 53.325 104.500 148.295 104.585 ;
        POLYGON 148.295 104.585 148.325 104.585 148.295 104.500 ;
        POLYGON 232.490 104.585 232.490 104.500 232.370 104.500 ;
        RECT 232.490 104.500 303.120 104.585 ;
        RECT 53.325 104.440 148.120 104.500 ;
        RECT 27.225 103.685 31.250 104.440 ;
        POLYGON 23.730 103.685 23.730 99.165 22.040 99.165 ;
        RECT 23.730 99.165 31.250 103.685 ;
        POLYGON 22.040 99.165 22.040 95.610 20.715 95.610 ;
        RECT 22.040 99.020 31.250 99.165 ;
        POLYGON 31.250 104.440 33.520 104.440 31.250 99.020 ;
        POLYGON 53.145 104.440 53.145 100.840 51.955 100.840 ;
        RECT 53.145 103.990 148.120 104.440 ;
        POLYGON 148.120 104.500 148.295 104.500 148.120 103.995 ;
        POLYGON 232.370 104.500 232.370 103.995 231.640 103.995 ;
        RECT 232.370 103.995 303.120 104.500 ;
        POLYGON 231.640 103.995 231.640 103.990 231.635 103.990 ;
        RECT 231.640 103.990 303.120 103.995 ;
        RECT 53.145 103.975 148.115 103.990 ;
        POLYGON 148.115 103.990 148.120 103.990 148.115 103.980 ;
        POLYGON 231.635 103.990 231.635 103.980 231.620 103.980 ;
        RECT 231.635 103.980 303.120 103.990 ;
        POLYGON 231.620 103.980 231.620 103.975 231.610 103.975 ;
        RECT 231.620 103.975 303.120 103.980 ;
        RECT 53.145 103.400 147.915 103.975 ;
        POLYGON 147.915 103.975 148.115 103.975 147.915 103.405 ;
        POLYGON 231.610 103.975 231.610 103.970 231.605 103.970 ;
        RECT 231.610 103.970 303.120 103.975 ;
        POLYGON 231.605 103.970 231.605 103.850 231.435 103.850 ;
        RECT 231.605 103.850 303.120 103.970 ;
        POLYGON 231.435 103.850 231.435 103.405 230.795 103.405 ;
        RECT 231.435 103.405 303.120 103.850 ;
        RECT 53.145 102.875 147.735 103.400 ;
        POLYGON 147.735 103.400 147.915 103.400 147.735 102.875 ;
        POLYGON 230.795 103.405 230.795 102.875 230.030 102.875 ;
        RECT 230.795 102.875 303.120 103.405 ;
        RECT 53.145 102.660 147.660 102.875 ;
        POLYGON 147.660 102.875 147.735 102.875 147.660 102.660 ;
        POLYGON 230.030 102.875 230.030 102.870 230.025 102.870 ;
        RECT 230.030 102.870 303.120 102.875 ;
        POLYGON 230.025 102.870 230.025 102.660 229.755 102.660 ;
        RECT 230.025 102.660 303.120 102.870 ;
        RECT 53.145 102.630 147.650 102.660 ;
        POLYGON 147.650 102.660 147.660 102.660 147.650 102.635 ;
        POLYGON 229.755 102.660 229.755 102.635 229.725 102.635 ;
        RECT 229.755 102.635 303.120 102.660 ;
        RECT 53.145 101.790 147.390 102.630 ;
        POLYGON 147.390 102.630 147.650 102.630 147.390 101.795 ;
        POLYGON 229.725 102.635 229.725 101.795 228.645 101.795 ;
        RECT 229.725 101.795 303.120 102.635 ;
        RECT 53.145 101.525 147.310 101.790 ;
        POLYGON 147.310 101.790 147.390 101.790 147.310 101.530 ;
        POLYGON 228.645 101.795 228.645 101.530 228.305 101.530 ;
        RECT 228.645 101.530 303.120 101.795 ;
        POLYGON 228.305 101.530 228.305 101.525 228.300 101.525 ;
        RECT 228.305 101.525 303.120 101.530 ;
        RECT 53.145 101.285 147.235 101.525 ;
        POLYGON 147.235 101.525 147.310 101.525 147.235 101.285 ;
        POLYGON 228.300 101.525 228.300 101.285 227.990 101.285 ;
        RECT 228.300 101.285 303.120 101.525 ;
        RECT 53.145 100.840 147.090 101.285 ;
        POLYGON 51.955 100.840 51.955 99.020 51.460 99.020 ;
        RECT 51.955 100.815 147.090 100.840 ;
        POLYGON 147.090 101.285 147.235 101.285 147.090 100.820 ;
        POLYGON 227.990 101.285 227.990 100.820 227.395 100.820 ;
        RECT 227.990 100.820 303.120 101.285 ;
        POLYGON 227.395 100.820 227.395 100.815 227.390 100.815 ;
        RECT 227.395 100.815 303.120 100.820 ;
        RECT 51.955 100.670 147.045 100.815 ;
        POLYGON 147.045 100.815 147.090 100.815 147.045 100.675 ;
        POLYGON 227.390 100.815 227.390 100.675 227.210 100.675 ;
        RECT 227.390 100.675 303.120 100.815 ;
        POLYGON 227.210 100.675 227.210 100.670 227.200 100.670 ;
        RECT 227.210 100.670 303.120 100.675 ;
        RECT 51.955 100.590 147.020 100.670 ;
        POLYGON 147.020 100.670 147.045 100.670 147.020 100.590 ;
        POLYGON 227.200 100.670 227.200 100.590 227.100 100.590 ;
        RECT 227.200 100.590 303.120 100.670 ;
        RECT 51.955 100.545 147.005 100.590 ;
        POLYGON 147.005 100.590 147.020 100.590 147.005 100.550 ;
        POLYGON 227.100 100.590 227.100 100.550 227.050 100.550 ;
        RECT 227.100 100.550 303.120 100.590 ;
        RECT 51.955 100.335 146.940 100.545 ;
        POLYGON 146.940 100.545 147.005 100.545 146.940 100.340 ;
        POLYGON 227.050 100.550 227.050 100.385 226.865 100.385 ;
        RECT 227.050 100.385 303.120 100.550 ;
        POLYGON 226.865 100.385 226.865 100.340 226.815 100.340 ;
        RECT 226.865 100.340 303.120 100.385 ;
        RECT 51.955 100.075 146.860 100.335 ;
        POLYGON 146.860 100.335 146.940 100.335 146.860 100.075 ;
        POLYGON 226.815 100.340 226.815 100.075 226.510 100.075 ;
        RECT 226.815 100.075 303.120 100.340 ;
        RECT 51.955 100.045 146.855 100.075 ;
        POLYGON 146.855 100.075 146.860 100.075 146.855 100.045 ;
        POLYGON 226.510 100.075 226.510 100.045 226.475 100.045 ;
        RECT 226.510 100.045 303.120 100.075 ;
        RECT 51.955 99.865 146.805 100.045 ;
        POLYGON 146.805 100.045 146.855 100.045 146.805 99.870 ;
        POLYGON 226.475 100.045 226.475 99.870 226.275 99.870 ;
        RECT 226.475 99.870 303.120 100.045 ;
        RECT 51.955 99.465 146.695 99.865 ;
        POLYGON 146.695 99.865 146.805 99.865 146.695 99.465 ;
        POLYGON 226.275 99.870 226.275 99.465 225.810 99.465 ;
        RECT 226.275 99.465 303.120 99.870 ;
        RECT 51.955 99.425 146.685 99.465 ;
        POLYGON 146.685 99.465 146.695 99.465 146.685 99.430 ;
        POLYGON 225.810 99.465 225.810 99.430 225.770 99.430 ;
        RECT 225.810 99.430 303.120 99.465 ;
        POLYGON 225.770 99.430 225.770 99.425 225.765 99.425 ;
        RECT 225.770 99.425 303.120 99.430 ;
        RECT 51.955 99.020 146.570 99.425 ;
        RECT 22.040 98.805 31.170 99.020 ;
        POLYGON 31.170 99.020 31.250 99.020 31.170 98.805 ;
        POLYGON 51.460 99.020 51.460 98.930 51.435 98.930 ;
        RECT 51.460 99.005 146.570 99.020 ;
        POLYGON 146.570 99.425 146.685 99.425 146.570 99.010 ;
        POLYGON 225.765 99.425 225.765 99.010 225.290 99.010 ;
        RECT 225.765 99.010 303.120 99.425 ;
        POLYGON 225.290 99.010 225.290 99.005 225.285 99.005 ;
        RECT 225.290 99.005 303.120 99.010 ;
        RECT 51.460 98.930 146.510 99.005 ;
        POLYGON 51.435 98.930 51.435 98.805 51.400 98.805 ;
        RECT 51.435 98.805 146.510 98.930 ;
        RECT 22.040 95.610 29.215 98.805 ;
        POLYGON 20.715 95.610 20.715 87.330 18.180 87.330 ;
        RECT 20.715 93.500 29.215 95.610 ;
        POLYGON 29.215 98.805 31.170 98.805 29.215 93.500 ;
        POLYGON 51.400 98.805 51.400 98.210 51.235 98.210 ;
        RECT 51.400 98.795 146.510 98.805 ;
        POLYGON 146.510 99.005 146.570 99.005 146.510 98.800 ;
        POLYGON 225.285 99.005 225.285 98.800 225.050 98.800 ;
        RECT 225.285 98.800 303.120 99.005 ;
        RECT 51.400 98.610 146.460 98.795 ;
        POLYGON 146.460 98.795 146.510 98.795 146.460 98.615 ;
        POLYGON 225.050 98.800 225.050 98.615 224.840 98.615 ;
        RECT 225.050 98.615 303.120 98.800 ;
        RECT 51.400 98.355 146.390 98.610 ;
        POLYGON 146.390 98.610 146.460 98.610 146.390 98.360 ;
        POLYGON 224.840 98.615 224.840 98.360 224.545 98.360 ;
        RECT 224.840 98.360 303.120 98.615 ;
        POLYGON 224.545 98.360 224.545 98.355 224.540 98.355 ;
        RECT 224.545 98.355 303.120 98.360 ;
        RECT 51.400 98.225 146.355 98.355 ;
        POLYGON 146.355 98.355 146.390 98.355 146.355 98.230 ;
        POLYGON 224.540 98.355 224.540 98.230 224.400 98.230 ;
        RECT 224.540 98.230 303.120 98.355 ;
        POLYGON 224.400 98.230 224.400 98.225 224.390 98.225 ;
        RECT 224.400 98.225 303.120 98.230 ;
        RECT 51.400 98.210 146.150 98.225 ;
        POLYGON 51.235 98.210 51.235 96.665 50.815 96.665 ;
        RECT 51.235 97.490 146.150 98.210 ;
        POLYGON 146.150 98.225 146.355 98.225 146.150 97.495 ;
        POLYGON 224.390 98.225 224.390 98.140 224.295 98.140 ;
        RECT 224.390 98.140 303.120 98.225 ;
        POLYGON 224.295 98.140 224.295 97.495 223.640 97.495 ;
        RECT 224.295 97.495 303.120 98.140 ;
        RECT 51.235 97.470 146.145 97.490 ;
        POLYGON 146.145 97.490 146.150 97.490 146.145 97.470 ;
        POLYGON 223.640 97.495 223.640 97.470 223.610 97.470 ;
        RECT 223.640 97.470 303.120 97.495 ;
        RECT 51.235 97.160 146.070 97.470 ;
        POLYGON 146.070 97.470 146.145 97.470 146.070 97.165 ;
        POLYGON 223.610 97.470 223.610 97.165 223.300 97.165 ;
        RECT 223.610 97.165 303.120 97.470 ;
        RECT 51.235 96.840 145.995 97.160 ;
        POLYGON 145.995 97.160 146.070 97.160 145.995 96.850 ;
        POLYGON 223.300 97.165 223.300 96.850 222.980 96.850 ;
        RECT 223.300 96.850 303.120 97.165 ;
        RECT 51.235 96.810 145.985 96.840 ;
        POLYGON 145.985 96.840 145.995 96.840 145.985 96.815 ;
        POLYGON 222.980 96.850 222.980 96.815 222.945 96.815 ;
        RECT 222.980 96.815 303.120 96.850 ;
        RECT 51.235 96.665 145.945 96.810 ;
        POLYGON 50.815 96.665 50.815 93.500 50.120 93.500 ;
        RECT 50.815 96.645 145.945 96.665 ;
        POLYGON 145.945 96.810 145.985 96.810 145.945 96.645 ;
        POLYGON 222.945 96.815 222.945 96.805 222.935 96.805 ;
        RECT 222.945 96.805 303.120 96.815 ;
        POLYGON 222.935 96.805 222.935 96.645 222.770 96.645 ;
        RECT 222.935 96.645 303.120 96.805 ;
        RECT 50.815 96.530 145.920 96.645 ;
        POLYGON 145.920 96.645 145.945 96.645 145.920 96.540 ;
        POLYGON 222.770 96.645 222.770 96.540 222.665 96.540 ;
        RECT 222.770 96.540 303.120 96.645 ;
        RECT 50.815 96.470 145.905 96.530 ;
        POLYGON 145.905 96.530 145.920 96.530 145.905 96.480 ;
        POLYGON 222.665 96.540 222.665 96.480 222.605 96.480 ;
        RECT 222.665 96.480 303.120 96.540 ;
        POLYGON 222.605 96.480 222.605 96.470 222.595 96.470 ;
        RECT 222.605 96.470 303.120 96.480 ;
        RECT 50.815 96.355 145.875 96.470 ;
        POLYGON 145.875 96.470 145.905 96.470 145.875 96.355 ;
        POLYGON 222.595 96.470 222.595 96.355 222.475 96.355 ;
        RECT 222.595 96.355 303.120 96.470 ;
        RECT 50.815 96.145 145.825 96.355 ;
        POLYGON 145.825 96.355 145.875 96.355 145.825 96.155 ;
        POLYGON 222.475 96.355 222.475 96.155 222.270 96.155 ;
        RECT 222.475 96.155 303.120 96.355 ;
        RECT 50.815 96.055 145.805 96.145 ;
        POLYGON 145.805 96.145 145.825 96.145 145.805 96.065 ;
        POLYGON 222.270 96.155 222.270 96.065 222.180 96.065 ;
        RECT 222.270 96.065 303.120 96.155 ;
        POLYGON 222.180 96.065 222.180 96.055 222.170 96.055 ;
        RECT 222.180 96.055 303.120 96.065 ;
        RECT 50.815 95.860 145.755 96.055 ;
        POLYGON 145.755 96.055 145.805 96.055 145.755 95.865 ;
        POLYGON 222.170 96.055 222.170 95.865 221.975 95.865 ;
        RECT 222.170 95.865 303.120 96.055 ;
        RECT 50.815 94.845 145.510 95.860 ;
        POLYGON 145.510 95.860 145.755 95.860 145.510 94.845 ;
        POLYGON 221.975 95.865 221.975 95.585 221.690 95.585 ;
        RECT 221.975 95.585 303.120 95.865 ;
        POLYGON 221.690 95.585 221.690 94.845 221.020 94.845 ;
        RECT 221.690 94.845 303.120 95.585 ;
        RECT 50.815 94.745 145.490 94.845 ;
        POLYGON 145.490 94.845 145.510 94.845 145.490 94.750 ;
        POLYGON 221.020 94.845 221.020 94.750 220.935 94.750 ;
        RECT 221.020 94.750 303.120 94.845 ;
        POLYGON 220.935 94.750 220.935 94.745 220.930 94.745 ;
        RECT 220.935 94.745 303.120 94.750 ;
        RECT 50.815 94.605 145.460 94.745 ;
        POLYGON 145.460 94.745 145.490 94.745 145.460 94.615 ;
        POLYGON 220.930 94.745 220.930 94.615 220.810 94.615 ;
        RECT 220.930 94.615 303.120 94.745 ;
        RECT 50.815 93.655 145.265 94.605 ;
        POLYGON 145.265 94.605 145.460 94.605 145.265 93.665 ;
        POLYGON 220.810 94.615 220.810 93.665 219.950 93.665 ;
        RECT 220.810 93.665 303.120 94.615 ;
        POLYGON 219.950 93.665 219.950 93.655 219.940 93.655 ;
        RECT 219.950 93.655 303.120 93.665 ;
        RECT 50.815 93.500 145.020 93.655 ;
        RECT 20.715 87.885 27.420 93.500 ;
        POLYGON 27.420 93.500 29.215 93.500 27.420 87.885 ;
        POLYGON 50.120 93.500 50.120 92.455 49.890 92.455 ;
        RECT 50.120 92.635 145.020 93.500 ;
        RECT 50.120 92.630 124.065 92.635 ;
        POLYGON 124.065 92.635 124.070 92.635 124.065 92.630 ;
        RECT 50.120 92.615 124.055 92.630 ;
        POLYGON 124.055 92.630 124.065 92.630 124.055 92.615 ;
        POLYGON 124.070 92.630 124.070 92.615 124.065 92.615 ;
        RECT 124.070 92.615 145.020 92.635 ;
        RECT 50.120 92.580 124.025 92.615 ;
        POLYGON 124.025 92.615 124.055 92.615 124.025 92.580 ;
        POLYGON 124.065 92.610 124.065 92.580 124.055 92.580 ;
        RECT 124.065 92.580 145.020 92.615 ;
        RECT 50.120 92.485 123.945 92.580 ;
        POLYGON 123.945 92.580 124.025 92.580 123.945 92.485 ;
        POLYGON 124.055 92.580 124.055 92.485 124.025 92.485 ;
        RECT 124.055 92.490 145.020 92.580 ;
        POLYGON 145.020 93.655 145.265 93.655 145.020 92.490 ;
        POLYGON 219.940 93.655 219.940 92.910 219.265 92.910 ;
        RECT 219.940 92.910 303.120 93.655 ;
        POLYGON 219.265 92.910 219.265 92.490 218.930 92.490 ;
        RECT 219.265 92.490 303.120 92.910 ;
        RECT 124.055 92.485 144.985 92.490 ;
        RECT 50.120 92.480 123.940 92.485 ;
        POLYGON 123.940 92.485 123.945 92.485 123.940 92.480 ;
        RECT 50.120 92.455 123.810 92.480 ;
        POLYGON 49.890 92.455 49.890 88.230 49.195 88.230 ;
        RECT 49.890 92.330 123.810 92.455 ;
        POLYGON 123.810 92.480 123.940 92.480 123.810 92.330 ;
        POLYGON 124.025 92.480 124.025 92.330 123.975 92.330 ;
        RECT 124.025 92.330 144.985 92.485 ;
        POLYGON 144.985 92.490 145.020 92.490 144.985 92.330 ;
        POLYGON 218.930 92.490 218.930 92.390 218.850 92.390 ;
        RECT 218.930 92.390 303.120 92.490 ;
        POLYGON 218.850 92.390 218.850 92.330 218.800 92.330 ;
        RECT 218.850 92.330 303.120 92.390 ;
        RECT 49.890 91.810 123.380 92.330 ;
        POLYGON 123.380 92.330 123.810 92.330 123.380 91.810 ;
        POLYGON 123.975 92.325 123.975 92.280 123.960 92.280 ;
        RECT 123.975 92.320 144.985 92.330 ;
        RECT 123.975 92.280 144.975 92.320 ;
        POLYGON 123.960 92.275 123.960 91.810 123.810 91.810 ;
        RECT 123.960 92.270 144.975 92.280 ;
        POLYGON 144.975 92.320 144.985 92.320 144.975 92.275 ;
        POLYGON 218.800 92.330 218.800 92.280 218.760 92.280 ;
        RECT 218.800 92.280 303.120 92.330 ;
        RECT 123.960 92.200 144.960 92.270 ;
        POLYGON 144.960 92.270 144.975 92.270 144.960 92.200 ;
        POLYGON 218.760 92.275 218.760 92.205 218.700 92.205 ;
        RECT 218.760 92.205 303.120 92.280 ;
        RECT 123.960 91.810 144.885 92.200 ;
        RECT 49.890 91.765 123.345 91.810 ;
        POLYGON 123.345 91.810 123.380 91.810 123.345 91.765 ;
        POLYGON 123.810 91.810 123.810 91.765 123.795 91.765 ;
        RECT 123.810 91.770 144.885 91.810 ;
        POLYGON 144.885 92.200 144.960 92.200 144.885 91.770 ;
        POLYGON 218.700 92.200 218.700 91.770 218.355 91.770 ;
        RECT 218.700 91.770 303.120 92.205 ;
        RECT 123.810 91.765 144.810 91.770 ;
        RECT 49.890 91.345 122.995 91.765 ;
        POLYGON 122.995 91.765 123.345 91.765 122.995 91.345 ;
        POLYGON 123.795 91.765 123.795 91.355 123.665 91.355 ;
        RECT 123.795 91.355 144.810 91.765 ;
        POLYGON 123.665 91.350 123.665 91.345 123.660 91.345 ;
        RECT 123.665 91.345 144.810 91.355 ;
        POLYGON 144.810 91.770 144.885 91.770 144.810 91.350 ;
        POLYGON 218.355 91.770 218.355 91.350 218.015 91.350 ;
        RECT 218.355 91.350 303.120 91.770 ;
        RECT 49.890 91.150 122.830 91.345 ;
        POLYGON 122.830 91.345 122.995 91.345 122.830 91.150 ;
        RECT 123.660 91.340 144.810 91.345 ;
        POLYGON 123.660 91.340 123.660 91.165 123.605 91.165 ;
        RECT 123.660 91.165 144.780 91.340 ;
        POLYGON 144.780 91.340 144.810 91.340 144.780 91.170 ;
        POLYGON 218.015 91.345 218.015 91.170 217.875 91.170 ;
        RECT 218.015 91.170 303.120 91.350 ;
        RECT 123.605 91.160 144.780 91.165 ;
        POLYGON 217.875 91.170 217.875 91.160 217.865 91.160 ;
        RECT 217.875 91.160 303.120 91.170 ;
        POLYGON 123.605 91.160 123.605 91.150 123.600 91.150 ;
        RECT 123.605 91.150 144.605 91.160 ;
        RECT 49.890 90.770 122.545 91.150 ;
        POLYGON 122.545 91.150 122.830 91.150 122.545 90.770 ;
        POLYGON 123.600 91.150 123.600 90.775 123.480 90.775 ;
        RECT 123.600 90.775 144.605 91.150 ;
        RECT 49.890 90.145 122.080 90.770 ;
        POLYGON 122.080 90.770 122.545 90.770 122.080 90.145 ;
        POLYGON 123.480 90.770 123.480 90.155 123.280 90.155 ;
        RECT 123.480 90.155 144.605 90.775 ;
        POLYGON 144.605 91.160 144.780 91.160 144.605 90.170 ;
        POLYGON 217.865 91.160 217.865 90.735 217.525 90.735 ;
        RECT 217.865 90.735 303.120 91.160 ;
        POLYGON 217.525 90.735 217.525 90.170 217.070 90.170 ;
        RECT 217.525 90.170 303.120 90.735 ;
        RECT 49.890 88.960 121.200 90.145 ;
        POLYGON 121.200 90.145 122.080 90.145 121.200 88.960 ;
        POLYGON 123.280 90.145 123.280 88.965 122.900 88.965 ;
        RECT 123.280 89.540 144.495 90.155 ;
        POLYGON 144.495 90.155 144.605 90.155 144.495 89.540 ;
        POLYGON 217.070 90.170 217.070 90.155 217.055 90.155 ;
        RECT 217.070 90.155 303.120 90.170 ;
        POLYGON 217.055 90.150 217.055 90.115 217.025 90.115 ;
        RECT 217.055 90.115 303.120 90.155 ;
        POLYGON 217.025 90.115 217.025 89.540 216.620 89.540 ;
        RECT 217.025 89.540 303.120 90.115 ;
        RECT 123.280 88.965 144.415 89.540 ;
        POLYGON 144.415 89.540 144.495 89.540 144.415 88.975 ;
        POLYGON 216.620 89.540 216.620 88.975 216.220 88.975 ;
        RECT 216.620 88.975 303.120 89.540 ;
        POLYGON 216.220 88.970 216.220 88.965 216.215 88.965 ;
        RECT 216.220 88.965 303.120 88.975 ;
        RECT 49.890 88.565 120.905 88.960 ;
        POLYGON 120.905 88.960 121.200 88.960 120.905 88.565 ;
        POLYGON 122.900 88.960 122.900 88.580 122.780 88.580 ;
        RECT 122.900 88.580 144.360 88.965 ;
        POLYGON 144.360 88.965 144.415 88.965 144.360 88.590 ;
        POLYGON 216.215 88.965 216.215 88.590 215.950 88.590 ;
        RECT 216.215 88.590 303.120 88.965 ;
        RECT 122.780 88.575 144.360 88.580 ;
        POLYGON 215.950 88.590 215.950 88.575 215.940 88.575 ;
        RECT 215.950 88.575 303.120 88.590 ;
        POLYGON 122.780 88.575 122.780 88.565 122.775 88.565 ;
        RECT 122.780 88.565 144.355 88.575 ;
        RECT 49.890 88.540 120.890 88.565 ;
        POLYGON 120.890 88.565 120.905 88.565 120.890 88.540 ;
        POLYGON 122.775 88.565 122.775 88.540 122.765 88.540 ;
        RECT 122.775 88.540 144.355 88.565 ;
        POLYGON 144.355 88.575 144.360 88.575 144.355 88.555 ;
        POLYGON 215.940 88.575 215.940 88.555 215.925 88.555 ;
        RECT 215.940 88.555 303.120 88.575 ;
        POLYGON 215.925 88.550 215.925 88.540 215.915 88.540 ;
        RECT 215.925 88.540 303.120 88.555 ;
        RECT 49.890 88.230 120.350 88.540 ;
        POLYGON 49.195 88.230 49.195 87.885 49.155 87.885 ;
        RECT 49.195 87.885 120.350 88.230 ;
        RECT 20.715 87.330 27.225 87.885 ;
        POLYGON 18.180 87.330 18.180 78.870 16.145 78.870 ;
        RECT 18.180 87.160 27.225 87.330 ;
        POLYGON 27.225 87.885 27.420 87.885 27.225 87.160 ;
        POLYGON 49.155 87.870 49.155 87.160 49.075 87.160 ;
        RECT 49.155 87.730 120.350 87.885 ;
        POLYGON 120.350 88.540 120.890 88.540 120.350 87.730 ;
        POLYGON 122.765 88.535 122.765 88.110 122.630 88.110 ;
        RECT 122.765 88.110 144.290 88.540 ;
        POLYGON 122.630 88.105 122.630 87.845 122.545 87.845 ;
        RECT 122.630 88.095 144.290 88.110 ;
        POLYGON 144.290 88.540 144.355 88.540 144.290 88.105 ;
        POLYGON 215.915 88.540 215.915 88.105 215.610 88.105 ;
        RECT 215.915 88.105 303.120 88.540 ;
        RECT 122.630 87.845 144.240 88.095 ;
        POLYGON 122.545 87.845 122.545 87.740 122.515 87.740 ;
        RECT 122.545 87.740 144.240 87.845 ;
        POLYGON 144.240 88.095 144.290 88.095 144.240 87.745 ;
        POLYGON 215.610 88.105 215.610 87.745 215.355 87.745 ;
        RECT 215.610 87.745 303.120 88.105 ;
        RECT 49.155 87.160 119.810 87.730 ;
        RECT 18.180 82.175 25.870 87.160 ;
        POLYGON 25.870 87.160 27.225 87.160 25.870 82.175 ;
        POLYGON 49.075 87.145 49.075 83.980 48.725 83.980 ;
        RECT 49.075 86.915 119.810 87.160 ;
        POLYGON 119.810 87.730 120.350 87.730 119.810 86.915 ;
        POLYGON 122.515 87.730 122.515 87.170 122.360 87.170 ;
        RECT 122.515 87.170 144.160 87.740 ;
        POLYGON 144.160 87.740 144.240 87.740 144.160 87.180 ;
        POLYGON 215.355 87.740 215.355 87.210 214.980 87.210 ;
        RECT 215.355 87.210 303.120 87.745 ;
        POLYGON 214.980 87.210 214.980 87.180 214.960 87.180 ;
        RECT 214.980 87.180 303.120 87.210 ;
        POLYGON 214.960 87.180 214.960 87.175 214.955 87.175 ;
        RECT 214.960 87.175 303.120 87.180 ;
        POLYGON 122.360 87.165 122.360 86.925 122.295 86.925 ;
        RECT 122.360 86.925 144.125 87.170 ;
        POLYGON 144.125 87.170 144.160 87.170 144.125 86.935 ;
        POLYGON 214.955 87.170 214.955 87.015 214.850 87.015 ;
        RECT 214.955 87.015 303.120 87.175 ;
        POLYGON 214.850 87.015 214.850 86.935 214.800 86.935 ;
        RECT 214.850 86.935 303.120 87.015 ;
        POLYGON 214.800 86.935 214.800 86.930 214.795 86.930 ;
        RECT 214.800 86.930 303.120 86.935 ;
        POLYGON 122.295 86.925 122.295 86.915 122.290 86.915 ;
        RECT 122.295 86.915 144.115 86.925 ;
        RECT 49.075 86.500 119.535 86.915 ;
        POLYGON 119.535 86.915 119.810 86.915 119.535 86.500 ;
        POLYGON 122.290 86.905 122.290 86.505 122.180 86.505 ;
        RECT 122.290 86.865 144.115 86.915 ;
        POLYGON 144.115 86.925 144.125 86.925 144.115 86.865 ;
        POLYGON 214.795 86.925 214.795 86.865 214.755 86.865 ;
        RECT 214.795 86.865 303.120 86.930 ;
        RECT 122.290 86.505 144.010 86.865 ;
        RECT 49.075 85.905 119.135 86.500 ;
        POLYGON 119.135 86.500 119.535 86.500 119.135 85.905 ;
        POLYGON 122.180 86.500 122.180 85.915 122.020 85.915 ;
        RECT 122.180 85.915 144.010 86.505 ;
        POLYGON 144.010 86.865 144.115 86.865 144.010 85.920 ;
        POLYGON 214.755 86.865 214.755 86.505 214.525 86.505 ;
        RECT 214.755 86.505 303.120 86.865 ;
        POLYGON 214.525 86.500 214.525 85.920 214.155 85.920 ;
        RECT 214.525 85.920 303.120 86.505 ;
        RECT 49.075 85.245 118.750 85.905 ;
        POLYGON 118.750 85.905 119.135 85.905 118.750 85.245 ;
        POLYGON 122.020 85.905 122.020 85.255 121.840 85.255 ;
        RECT 122.020 85.255 143.935 85.915 ;
        POLYGON 143.935 85.915 144.010 85.915 143.935 85.255 ;
        POLYGON 214.155 85.915 214.155 85.720 214.030 85.720 ;
        RECT 214.155 85.720 303.120 85.920 ;
        POLYGON 214.030 85.720 214.030 85.255 213.750 85.255 ;
        RECT 214.030 85.255 303.120 85.720 ;
        RECT 121.840 85.250 143.935 85.255 ;
        RECT 49.075 83.980 118.000 85.245 ;
        POLYGON 48.725 83.980 48.725 82.205 48.625 82.205 ;
        RECT 48.725 83.970 118.000 83.980 ;
        POLYGON 118.000 85.245 118.750 85.245 118.000 83.970 ;
        POLYGON 121.840 85.245 121.840 84.090 121.525 84.090 ;
        RECT 121.840 84.935 143.900 85.250 ;
        POLYGON 143.900 85.250 143.935 85.250 143.900 84.935 ;
        POLYGON 213.750 85.250 213.750 84.935 213.560 84.935 ;
        RECT 213.750 84.935 303.120 85.255 ;
        RECT 121.840 84.175 143.815 84.935 ;
        POLYGON 143.815 84.935 143.900 84.935 143.815 84.175 ;
        POLYGON 213.560 84.935 213.560 84.205 213.125 84.205 ;
        RECT 213.560 84.205 303.120 84.935 ;
        POLYGON 213.125 84.205 213.125 84.175 213.110 84.175 ;
        RECT 213.125 84.175 303.120 84.205 ;
        RECT 121.840 84.090 143.810 84.175 ;
        POLYGON 143.810 84.175 143.815 84.175 143.810 84.090 ;
        POLYGON 213.110 84.175 213.110 84.095 213.065 84.095 ;
        RECT 213.110 84.095 303.120 84.175 ;
        POLYGON 121.525 84.090 121.525 83.970 121.490 83.970 ;
        RECT 121.525 84.080 143.810 84.090 ;
        RECT 121.525 83.970 143.795 84.080 ;
        RECT 48.725 83.175 117.530 83.970 ;
        POLYGON 117.530 83.970 118.000 83.970 117.530 83.175 ;
        POLYGON 121.490 83.960 121.490 83.795 121.445 83.795 ;
        RECT 121.490 83.795 143.795 83.970 ;
        POLYGON 121.445 83.790 121.445 83.780 121.440 83.780 ;
        RECT 121.445 83.780 143.795 83.795 ;
        POLYGON 143.795 84.080 143.810 84.080 143.795 83.790 ;
        POLYGON 213.065 84.090 213.065 83.845 212.930 83.845 ;
        RECT 213.065 83.845 303.120 84.095 ;
        POLYGON 212.930 83.845 212.930 83.790 212.900 83.790 ;
        RECT 212.930 83.790 303.120 83.845 ;
        RECT 121.440 83.775 143.795 83.780 ;
        POLYGON 212.900 83.790 212.900 83.775 212.890 83.775 ;
        RECT 212.900 83.775 303.120 83.790 ;
        POLYGON 121.440 83.775 121.440 83.730 121.425 83.730 ;
        RECT 121.440 83.730 143.790 83.775 ;
        POLYGON 143.790 83.775 143.795 83.775 143.790 83.730 ;
        POLYGON 159.075 83.775 159.075 83.730 157.505 83.730 ;
        RECT 159.075 83.770 159.455 83.775 ;
        POLYGON 159.455 83.775 160.505 83.770 159.455 83.770 ;
        RECT 159.075 83.740 160.850 83.770 ;
        POLYGON 160.850 83.770 161.710 83.740 160.850 83.740 ;
        POLYGON 212.890 83.770 212.890 83.750 212.875 83.750 ;
        RECT 212.890 83.755 303.120 83.775 ;
        RECT 212.890 83.750 253.990 83.755 ;
        RECT 212.875 83.745 253.990 83.750 ;
        POLYGON 253.990 83.755 254.220 83.755 253.990 83.745 ;
        POLYGON 254.290 83.755 254.625 83.755 254.625 83.750 ;
        RECT 254.625 83.750 303.120 83.755 ;
        POLYGON 255.160 83.750 255.495 83.750 255.495 83.745 ;
        RECT 255.495 83.745 303.120 83.750 ;
        POLYGON 212.875 83.745 212.875 83.740 212.870 83.740 ;
        RECT 212.875 83.740 253.395 83.745 ;
        RECT 159.075 83.730 161.735 83.740 ;
        POLYGON 161.735 83.740 161.865 83.730 161.735 83.730 ;
        POLYGON 212.870 83.735 212.870 83.730 212.865 83.730 ;
        RECT 212.870 83.730 253.395 83.740 ;
        POLYGON 253.395 83.745 253.975 83.745 253.395 83.730 ;
        POLYGON 255.495 83.745 255.830 83.745 255.830 83.740 ;
        RECT 255.830 83.740 303.120 83.745 ;
        POLYGON 255.905 83.740 256.115 83.740 256.115 83.730 ;
        RECT 256.115 83.730 303.120 83.740 ;
        POLYGON 121.425 83.720 121.425 83.710 121.420 83.710 ;
        RECT 121.425 83.710 143.790 83.730 ;
        POLYGON 157.495 83.730 157.495 83.720 157.305 83.720 ;
        RECT 157.495 83.720 161.965 83.730 ;
        POLYGON 157.305 83.720 157.305 83.710 157.145 83.710 ;
        RECT 157.305 83.710 161.965 83.720 ;
        POLYGON 121.420 83.705 121.420 83.665 121.410 83.665 ;
        RECT 121.420 83.665 143.790 83.710 ;
        RECT 121.410 83.660 143.790 83.665 ;
        POLYGON 157.140 83.710 157.140 83.660 156.370 83.660 ;
        RECT 157.140 83.705 161.965 83.710 ;
        POLYGON 161.965 83.730 162.565 83.705 161.965 83.705 ;
        POLYGON 212.865 83.725 212.865 83.710 212.855 83.710 ;
        RECT 212.865 83.715 252.820 83.730 ;
        POLYGON 252.820 83.730 253.380 83.730 252.820 83.715 ;
        POLYGON 256.115 83.730 256.330 83.730 256.330 83.720 ;
        RECT 256.330 83.720 303.120 83.730 ;
        POLYGON 256.330 83.720 256.455 83.720 256.455 83.715 ;
        RECT 256.455 83.715 303.120 83.720 ;
        RECT 212.865 83.710 252.715 83.715 ;
        POLYGON 252.715 83.715 252.815 83.715 252.715 83.710 ;
        POLYGON 256.455 83.715 256.585 83.715 256.585 83.710 ;
        RECT 256.585 83.710 303.120 83.715 ;
        RECT 212.855 83.705 252.570 83.710 ;
        POLYGON 252.570 83.710 252.710 83.710 252.570 83.705 ;
        POLYGON 256.585 83.710 256.715 83.710 256.715 83.705 ;
        RECT 256.715 83.705 303.120 83.710 ;
        RECT 157.140 83.660 162.565 83.705 ;
        POLYGON 121.410 83.660 121.410 83.610 121.395 83.610 ;
        RECT 121.410 83.610 143.785 83.660 ;
        POLYGON 143.785 83.660 143.790 83.660 143.785 83.610 ;
        POLYGON 156.370 83.660 156.370 83.610 155.615 83.610 ;
        RECT 156.370 83.610 162.565 83.660 ;
        POLYGON 121.395 83.610 121.395 83.520 121.370 83.520 ;
        RECT 121.395 83.595 143.785 83.610 ;
        RECT 121.395 83.520 143.780 83.595 ;
        POLYGON 143.780 83.595 143.785 83.595 143.780 83.520 ;
        POLYGON 155.615 83.610 155.615 83.520 154.815 83.520 ;
        RECT 155.615 83.580 162.565 83.610 ;
        POLYGON 162.565 83.705 164.145 83.580 162.565 83.580 ;
        POLYGON 212.855 83.705 212.855 83.590 212.790 83.590 ;
        RECT 212.855 83.665 251.985 83.705 ;
        POLYGON 251.985 83.705 252.570 83.705 251.985 83.665 ;
        POLYGON 256.715 83.705 257.105 83.705 257.105 83.690 ;
        RECT 257.105 83.690 303.120 83.705 ;
        POLYGON 257.110 83.690 257.340 83.690 257.340 83.680 ;
        RECT 257.340 83.680 303.120 83.690 ;
        POLYGON 257.340 83.680 257.485 83.680 257.485 83.665 ;
        RECT 257.485 83.665 303.120 83.680 ;
        RECT 212.855 83.640 251.655 83.665 ;
        POLYGON 251.655 83.665 251.985 83.665 251.655 83.640 ;
        POLYGON 257.495 83.665 257.655 83.665 257.655 83.650 ;
        RECT 257.655 83.650 303.120 83.665 ;
        POLYGON 257.660 83.650 257.785 83.650 257.785 83.640 ;
        RECT 257.785 83.640 303.120 83.650 ;
        RECT 212.855 83.600 251.105 83.640 ;
        POLYGON 251.105 83.640 251.650 83.640 251.105 83.600 ;
        POLYGON 257.785 83.640 258.295 83.640 258.295 83.600 ;
        RECT 258.295 83.600 303.120 83.640 ;
        RECT 212.855 83.590 250.985 83.600 ;
        POLYGON 250.985 83.600 251.105 83.600 250.985 83.590 ;
        POLYGON 258.295 83.600 258.415 83.600 258.415 83.590 ;
        RECT 258.415 83.590 303.120 83.600 ;
        POLYGON 212.790 83.590 212.790 83.585 212.785 83.585 ;
        RECT 212.790 83.585 250.945 83.590 ;
        POLYGON 250.945 83.590 250.970 83.590 250.945 83.585 ;
        POLYGON 258.415 83.590 258.475 83.590 258.475 83.585 ;
        RECT 258.475 83.585 303.120 83.590 ;
        RECT 155.615 83.560 164.145 83.580 ;
        POLYGON 164.145 83.580 164.290 83.560 164.145 83.560 ;
        POLYGON 212.785 83.580 212.785 83.575 212.780 83.575 ;
        RECT 212.785 83.575 250.495 83.585 ;
        POLYGON 212.780 83.570 212.780 83.560 212.770 83.560 ;
        RECT 212.780 83.560 250.495 83.575 ;
        RECT 155.615 83.520 164.295 83.560 ;
        POLYGON 121.370 83.520 121.370 83.445 121.350 83.445 ;
        RECT 121.370 83.495 143.780 83.520 ;
        RECT 121.370 83.445 143.775 83.495 ;
        POLYGON 121.350 83.440 121.350 83.320 121.315 83.320 ;
        RECT 121.350 83.400 143.775 83.445 ;
        POLYGON 143.775 83.495 143.780 83.495 143.775 83.440 ;
        POLYGON 154.815 83.520 154.815 83.440 154.070 83.440 ;
        RECT 154.815 83.440 164.295 83.520 ;
        RECT 121.350 83.320 143.770 83.400 ;
        POLYGON 121.315 83.315 121.315 83.215 121.285 83.215 ;
        RECT 121.315 83.305 143.770 83.320 ;
        POLYGON 143.770 83.400 143.775 83.400 143.770 83.315 ;
        POLYGON 154.070 83.440 154.070 83.315 153.345 83.315 ;
        RECT 154.070 83.405 164.295 83.440 ;
        POLYGON 164.295 83.560 165.405 83.405 164.295 83.405 ;
        POLYGON 212.770 83.555 212.770 83.410 212.690 83.410 ;
        RECT 212.770 83.535 250.495 83.560 ;
        POLYGON 250.495 83.585 250.945 83.585 250.495 83.535 ;
        POLYGON 258.475 83.585 258.655 83.585 258.655 83.570 ;
        RECT 258.655 83.570 303.120 83.585 ;
        POLYGON 258.660 83.570 258.775 83.570 258.775 83.560 ;
        RECT 258.775 83.560 303.120 83.570 ;
        POLYGON 258.775 83.560 258.970 83.560 258.970 83.535 ;
        RECT 258.970 83.535 303.120 83.560 ;
        RECT 212.770 83.500 250.200 83.535 ;
        POLYGON 250.200 83.535 250.495 83.535 250.200 83.500 ;
        POLYGON 258.970 83.535 259.250 83.535 259.250 83.500 ;
        RECT 259.250 83.500 303.120 83.535 ;
        RECT 212.770 83.410 249.465 83.500 ;
        POLYGON 249.465 83.500 250.200 83.500 249.465 83.410 ;
        POLYGON 259.250 83.500 259.450 83.500 259.450 83.475 ;
        RECT 259.450 83.475 303.120 83.500 ;
        POLYGON 259.450 83.475 259.815 83.475 259.815 83.425 ;
        RECT 259.815 83.425 303.120 83.475 ;
        POLYGON 259.820 83.425 259.935 83.425 259.935 83.410 ;
        RECT 259.935 83.410 303.120 83.425 ;
        POLYGON 212.690 83.410 212.690 83.405 212.685 83.405 ;
        RECT 212.690 83.405 249.345 83.410 ;
        RECT 154.070 83.390 165.410 83.405 ;
        POLYGON 165.410 83.405 165.525 83.390 165.410 83.390 ;
        POLYGON 212.685 83.400 212.685 83.395 212.680 83.395 ;
        RECT 212.685 83.395 249.345 83.405 ;
        POLYGON 249.345 83.410 249.465 83.410 249.345 83.395 ;
        POLYGON 259.935 83.410 260.050 83.410 260.050 83.395 ;
        RECT 260.050 83.395 303.120 83.410 ;
        RECT 212.680 83.390 249.315 83.395 ;
        POLYGON 249.315 83.395 249.345 83.395 249.315 83.390 ;
        POLYGON 260.050 83.395 260.085 83.395 260.085 83.390 ;
        RECT 260.085 83.390 303.120 83.395 ;
        RECT 154.070 83.315 165.525 83.390 ;
        RECT 121.315 83.215 143.765 83.305 ;
        POLYGON 143.765 83.305 143.770 83.305 143.765 83.215 ;
        POLYGON 153.340 83.315 153.340 83.215 152.745 83.215 ;
        RECT 153.340 83.255 165.525 83.315 ;
        POLYGON 165.525 83.390 166.205 83.255 165.525 83.255 ;
        POLYGON 212.680 83.390 212.680 83.255 212.605 83.255 ;
        RECT 212.680 83.255 248.495 83.390 ;
        POLYGON 248.495 83.390 249.315 83.390 248.495 83.255 ;
        POLYGON 260.085 83.390 260.165 83.390 260.165 83.380 ;
        RECT 260.165 83.380 303.120 83.390 ;
        POLYGON 260.165 83.380 260.580 83.380 260.580 83.310 ;
        RECT 260.580 83.310 303.120 83.380 ;
        POLYGON 260.585 83.310 260.880 83.310 260.880 83.255 ;
        RECT 260.880 83.255 303.120 83.310 ;
        RECT 153.340 83.215 166.205 83.255 ;
        POLYGON 121.285 83.205 121.285 83.175 121.275 83.175 ;
        RECT 121.285 83.175 143.765 83.215 ;
        POLYGON 152.745 83.215 152.745 83.175 152.575 83.175 ;
        RECT 152.745 83.175 166.205 83.215 ;
        POLYGON 166.205 83.255 166.615 83.175 166.205 83.175 ;
        POLYGON 212.605 83.255 212.605 83.175 212.560 83.175 ;
        RECT 212.605 83.175 247.770 83.255 ;
        RECT 48.725 82.690 117.280 83.175 ;
        POLYGON 117.280 83.175 117.530 83.175 117.280 82.690 ;
        POLYGON 121.275 83.170 121.275 83.150 121.270 83.150 ;
        RECT 121.275 83.150 143.760 83.175 ;
        POLYGON 143.760 83.175 143.765 83.175 143.760 83.150 ;
        POLYGON 152.575 83.175 152.575 83.150 152.465 83.150 ;
        RECT 152.575 83.150 166.620 83.175 ;
        POLYGON 121.270 83.150 121.270 82.940 121.210 82.940 ;
        RECT 121.270 83.110 143.760 83.150 ;
        RECT 121.270 82.940 143.750 83.110 ;
        POLYGON 143.750 83.110 143.760 83.110 143.750 82.940 ;
        POLYGON 152.465 83.150 152.465 82.940 151.550 82.940 ;
        RECT 152.465 83.100 166.620 83.150 ;
        POLYGON 166.620 83.175 166.995 83.100 166.620 83.100 ;
        POLYGON 212.560 83.175 212.560 83.115 212.525 83.115 ;
        RECT 212.560 83.130 247.770 83.175 ;
        POLYGON 247.770 83.255 248.495 83.255 247.770 83.130 ;
        POLYGON 260.880 83.255 260.965 83.255 260.965 83.240 ;
        RECT 260.965 83.240 303.120 83.255 ;
        POLYGON 260.970 83.240 261.165 83.240 261.165 83.205 ;
        RECT 261.165 83.205 303.120 83.240 ;
        POLYGON 261.170 83.205 261.535 83.205 261.535 83.140 ;
        RECT 261.535 83.140 303.120 83.205 ;
        POLYGON 261.535 83.140 261.575 83.140 261.575 83.130 ;
        RECT 261.575 83.130 303.120 83.140 ;
        RECT 212.560 83.115 247.700 83.130 ;
        POLYGON 247.700 83.130 247.770 83.130 247.700 83.115 ;
        POLYGON 261.575 83.130 261.640 83.130 261.640 83.115 ;
        RECT 261.640 83.115 303.120 83.130 ;
        POLYGON 212.525 83.110 212.525 83.105 212.520 83.105 ;
        RECT 212.525 83.105 247.125 83.115 ;
        RECT 152.465 82.940 166.995 83.100 ;
        POLYGON 121.210 82.930 121.210 82.690 121.145 82.690 ;
        RECT 121.210 82.915 143.750 82.940 ;
        RECT 121.210 82.690 143.740 82.915 ;
        POLYGON 143.740 82.915 143.750 82.915 143.740 82.725 ;
        POLYGON 151.550 82.940 151.550 82.725 150.735 82.725 ;
        RECT 151.550 82.755 166.995 82.940 ;
        POLYGON 166.995 83.100 168.440 82.755 166.995 82.755 ;
        POLYGON 212.520 83.100 212.520 82.760 212.330 82.760 ;
        RECT 212.520 82.995 247.125 83.105 ;
        POLYGON 247.125 83.115 247.700 83.115 247.125 82.995 ;
        POLYGON 261.640 83.115 261.685 83.115 261.685 83.105 ;
        RECT 261.685 83.105 303.120 83.115 ;
        POLYGON 261.690 83.105 262.110 83.105 262.110 83.010 ;
        RECT 262.110 83.010 303.120 83.105 ;
        POLYGON 262.115 83.010 262.180 83.010 262.180 82.995 ;
        RECT 262.180 82.995 303.120 83.010 ;
        RECT 212.520 82.990 247.120 82.995 ;
        POLYGON 247.120 82.995 247.125 82.995 247.120 82.990 ;
        POLYGON 262.180 82.995 262.200 82.995 262.200 82.990 ;
        RECT 262.200 82.990 303.120 82.995 ;
        RECT 212.520 82.980 247.075 82.990 ;
        POLYGON 247.075 82.990 247.120 82.990 247.075 82.980 ;
        POLYGON 262.200 82.990 262.245 82.990 262.245 82.980 ;
        RECT 262.245 82.980 303.120 82.990 ;
        RECT 212.520 82.875 246.585 82.980 ;
        POLYGON 246.585 82.980 247.075 82.980 246.585 82.875 ;
        POLYGON 262.245 82.980 262.720 82.980 262.720 82.875 ;
        RECT 262.720 82.875 303.120 82.980 ;
        RECT 212.520 82.800 246.220 82.875 ;
        POLYGON 246.220 82.875 246.585 82.875 246.220 82.800 ;
        POLYGON 262.720 82.875 262.765 82.875 262.765 82.865 ;
        RECT 262.765 82.865 303.120 82.875 ;
        POLYGON 262.770 82.865 262.915 82.865 262.915 82.830 ;
        RECT 262.915 82.830 303.120 82.865 ;
        POLYGON 262.915 82.830 263.025 82.830 263.025 82.800 ;
        RECT 263.025 82.800 303.120 82.830 ;
        RECT 212.520 82.760 246.055 82.800 ;
        RECT 212.330 82.755 246.055 82.760 ;
        POLYGON 246.055 82.800 246.220 82.800 246.055 82.755 ;
        POLYGON 263.025 82.800 263.200 82.800 263.200 82.755 ;
        RECT 263.200 82.755 303.120 82.800 ;
        RECT 151.550 82.725 168.445 82.755 ;
        POLYGON 212.330 82.755 212.330 82.750 212.325 82.750 ;
        RECT 212.330 82.750 245.960 82.755 ;
        POLYGON 150.735 82.725 150.735 82.690 150.605 82.690 ;
        RECT 150.735 82.690 168.445 82.725 ;
        RECT 48.725 82.205 116.600 82.690 ;
        RECT 18.180 78.870 24.555 82.175 ;
        POLYGON 16.145 78.870 16.145 70.245 14.625 70.245 ;
        RECT 16.145 76.355 24.555 78.870 ;
        POLYGON 24.555 82.175 25.870 82.175 24.555 76.355 ;
        POLYGON 48.625 82.175 48.625 79.725 48.485 79.725 ;
        RECT 48.625 81.365 116.600 82.205 ;
        POLYGON 116.600 82.690 117.280 82.690 116.600 81.365 ;
        POLYGON 121.145 82.690 121.145 82.635 121.130 82.635 ;
        RECT 121.145 82.635 143.735 82.690 ;
        POLYGON 121.130 82.630 121.130 82.545 121.105 82.545 ;
        RECT 121.130 82.625 143.735 82.635 ;
        POLYGON 143.735 82.690 143.740 82.690 143.735 82.630 ;
        POLYGON 150.605 82.690 150.605 82.630 150.380 82.630 ;
        RECT 150.605 82.660 168.445 82.690 ;
        POLYGON 168.445 82.750 168.770 82.660 168.445 82.660 ;
        POLYGON 212.325 82.750 212.325 82.680 212.285 82.680 ;
        RECT 212.325 82.730 245.960 82.750 ;
        POLYGON 245.960 82.755 246.055 82.755 245.960 82.730 ;
        POLYGON 263.200 82.755 263.240 82.755 263.240 82.745 ;
        RECT 263.240 82.745 303.120 82.755 ;
        POLYGON 263.240 82.745 263.295 82.745 263.295 82.730 ;
        RECT 263.295 82.730 303.120 82.745 ;
        RECT 212.325 82.680 245.755 82.730 ;
        RECT 212.285 82.675 245.755 82.680 ;
        POLYGON 245.755 82.730 245.960 82.730 245.755 82.675 ;
        POLYGON 263.295 82.730 263.500 82.730 263.500 82.675 ;
        RECT 263.500 82.675 303.120 82.730 ;
        POLYGON 212.285 82.675 212.285 82.660 212.275 82.660 ;
        RECT 212.285 82.660 245.605 82.675 ;
        RECT 150.605 82.630 168.775 82.660 ;
        POLYGON 168.775 82.660 168.875 82.630 168.775 82.630 ;
        POLYGON 212.275 82.660 212.275 82.635 212.260 82.635 ;
        RECT 212.275 82.635 245.605 82.660 ;
        POLYGON 245.605 82.675 245.755 82.675 245.605 82.635 ;
        POLYGON 263.500 82.675 263.650 82.675 263.650 82.635 ;
        RECT 263.650 82.635 303.120 82.675 ;
        RECT 121.130 82.545 143.730 82.625 ;
        POLYGON 143.730 82.625 143.735 82.625 143.730 82.545 ;
        POLYGON 150.380 82.630 150.380 82.545 150.100 82.545 ;
        RECT 150.380 82.545 168.875 82.630 ;
        POLYGON 121.105 82.545 121.105 82.285 121.035 82.285 ;
        RECT 121.105 82.530 143.730 82.545 ;
        RECT 121.105 82.285 143.715 82.530 ;
        POLYGON 143.715 82.530 143.730 82.530 143.715 82.285 ;
        POLYGON 150.100 82.545 150.100 82.285 149.230 82.285 ;
        RECT 150.100 82.350 168.875 82.545 ;
        POLYGON 168.875 82.630 169.875 82.350 168.875 82.350 ;
        POLYGON 212.260 82.630 212.260 82.360 212.120 82.360 ;
        RECT 212.260 82.435 244.865 82.635 ;
        POLYGON 244.865 82.635 245.605 82.635 244.865 82.435 ;
        POLYGON 263.650 82.635 263.820 82.635 263.820 82.590 ;
        RECT 263.820 82.590 303.120 82.635 ;
        POLYGON 263.820 82.590 264.330 82.590 264.330 82.450 ;
        RECT 264.330 82.450 303.120 82.590 ;
        POLYGON 264.330 82.450 264.355 82.450 264.355 82.445 ;
        RECT 264.355 82.445 303.120 82.450 ;
        POLYGON 264.355 82.445 264.385 82.445 264.385 82.435 ;
        RECT 264.385 82.435 303.120 82.445 ;
        RECT 212.260 82.395 244.705 82.435 ;
        POLYGON 244.705 82.435 244.860 82.435 244.705 82.395 ;
        POLYGON 264.385 82.435 264.510 82.435 264.510 82.395 ;
        RECT 264.510 82.395 303.120 82.435 ;
        RECT 212.260 82.360 244.595 82.395 ;
        POLYGON 244.595 82.395 244.705 82.395 244.595 82.360 ;
        POLYGON 264.510 82.395 264.625 82.395 264.625 82.360 ;
        RECT 264.625 82.360 303.120 82.395 ;
        POLYGON 212.120 82.355 212.120 82.350 212.115 82.350 ;
        RECT 212.120 82.350 244.040 82.360 ;
        RECT 150.100 82.285 169.875 82.350 ;
        POLYGON 121.035 82.285 121.035 82.270 121.030 82.270 ;
        RECT 121.035 82.270 143.715 82.285 ;
        POLYGON 149.230 82.285 149.230 82.270 149.190 82.270 ;
        RECT 149.230 82.270 169.875 82.285 ;
        POLYGON 121.030 82.270 121.030 82.250 121.025 82.250 ;
        RECT 121.030 82.250 143.715 82.270 ;
        POLYGON 149.190 82.270 149.190 82.250 149.125 82.250 ;
        RECT 149.190 82.250 169.875 82.270 ;
        POLYGON 121.025 82.250 121.025 82.140 120.995 82.140 ;
        RECT 121.025 82.240 143.715 82.250 ;
        RECT 121.025 82.140 143.700 82.240 ;
        POLYGON 120.995 82.140 120.995 81.905 120.940 81.905 ;
        RECT 120.995 81.905 143.700 82.140 ;
        POLYGON 143.700 82.240 143.715 82.240 143.700 81.950 ;
        POLYGON 149.125 82.250 149.125 81.950 148.235 81.950 ;
        RECT 149.125 81.960 169.875 82.250 ;
        POLYGON 169.875 82.350 171.065 81.960 169.875 81.960 ;
        POLYGON 212.115 82.345 212.115 81.960 211.915 81.960 ;
        RECT 212.115 82.180 244.040 82.350 ;
        POLYGON 244.040 82.360 244.595 82.360 244.040 82.180 ;
        POLYGON 264.625 82.360 264.850 82.360 264.850 82.290 ;
        RECT 264.850 82.290 303.120 82.360 ;
        POLYGON 264.850 82.290 264.915 82.290 264.915 82.270 ;
        RECT 264.915 82.270 303.120 82.290 ;
        POLYGON 264.920 82.270 265.210 82.270 265.210 82.180 ;
        RECT 265.210 82.180 303.120 82.270 ;
        RECT 212.115 82.100 243.780 82.180 ;
        POLYGON 243.780 82.180 244.040 82.180 243.780 82.100 ;
        POLYGON 265.210 82.180 265.455 82.180 265.455 82.105 ;
        RECT 265.455 82.105 303.120 82.180 ;
        POLYGON 265.455 82.105 265.470 82.105 265.470 82.100 ;
        RECT 265.470 82.100 303.120 82.105 ;
        RECT 212.115 81.980 243.410 82.100 ;
        POLYGON 243.410 82.100 243.780 82.100 243.410 81.980 ;
        POLYGON 265.470 82.100 265.810 82.100 265.810 81.995 ;
        RECT 265.810 81.995 303.120 82.100 ;
        POLYGON 265.810 81.995 265.850 81.995 265.850 81.980 ;
        RECT 265.850 81.980 303.120 81.995 ;
        RECT 212.115 81.960 243.345 81.980 ;
        POLYGON 243.345 81.980 243.405 81.980 243.345 81.960 ;
        POLYGON 265.850 81.980 265.905 81.980 265.905 81.960 ;
        RECT 265.905 81.960 303.120 81.980 ;
        RECT 149.125 81.950 171.065 81.960 ;
        POLYGON 148.235 81.950 148.235 81.905 148.100 81.905 ;
        RECT 148.235 81.905 171.065 81.950 ;
        POLYGON 120.940 81.895 120.940 81.765 120.910 81.765 ;
        RECT 120.940 81.765 143.690 81.905 ;
        POLYGON 120.910 81.760 120.910 81.485 120.845 81.485 ;
        RECT 120.910 81.755 143.690 81.765 ;
        POLYGON 143.690 81.905 143.700 81.905 143.690 81.760 ;
        POLYGON 148.100 81.905 148.100 81.760 147.715 81.760 ;
        RECT 148.100 81.890 171.065 81.905 ;
        POLYGON 171.065 81.960 171.280 81.890 171.065 81.890 ;
        POLYGON 211.915 81.955 211.915 81.900 211.885 81.900 ;
        RECT 211.915 81.920 243.220 81.960 ;
        POLYGON 243.220 81.960 243.345 81.960 243.220 81.920 ;
        POLYGON 265.905 81.960 265.950 81.960 265.950 81.945 ;
        RECT 265.950 81.945 303.120 81.960 ;
        POLYGON 265.950 81.945 266.020 81.945 266.020 81.920 ;
        RECT 266.020 81.920 303.120 81.945 ;
        RECT 211.915 81.900 243.165 81.920 ;
        POLYGON 243.165 81.920 243.220 81.920 243.165 81.900 ;
        POLYGON 266.020 81.920 266.075 81.920 266.075 81.900 ;
        RECT 266.075 81.900 303.120 81.920 ;
        POLYGON 211.885 81.895 211.885 81.890 211.880 81.890 ;
        RECT 211.885 81.890 242.720 81.900 ;
        RECT 148.100 81.760 171.285 81.890 ;
        RECT 120.910 81.485 143.675 81.755 ;
        POLYGON 143.675 81.755 143.690 81.755 143.675 81.485 ;
        POLYGON 147.715 81.760 147.715 81.485 146.995 81.485 ;
        RECT 147.715 81.600 171.285 81.760 ;
        POLYGON 171.285 81.890 172.055 81.600 171.285 81.600 ;
        POLYGON 211.880 81.885 211.880 81.605 211.735 81.605 ;
        RECT 211.880 81.735 242.720 81.890 ;
        POLYGON 242.720 81.900 243.165 81.900 242.720 81.735 ;
        POLYGON 266.075 81.900 266.470 81.900 266.470 81.760 ;
        RECT 266.470 81.760 303.120 81.900 ;
        POLYGON 266.470 81.760 266.540 81.760 266.540 81.735 ;
        RECT 266.540 81.735 303.120 81.760 ;
        RECT 211.880 81.605 242.375 81.735 ;
        POLYGON 242.375 81.735 242.720 81.735 242.375 81.605 ;
        POLYGON 266.540 81.735 266.830 81.735 266.830 81.635 ;
        RECT 266.830 81.635 303.120 81.735 ;
        POLYGON 266.830 81.635 266.915 81.635 266.915 81.605 ;
        RECT 266.915 81.605 303.120 81.635 ;
        RECT 147.715 81.485 172.055 81.600 ;
        POLYGON 120.845 81.475 120.845 81.365 120.820 81.365 ;
        RECT 120.845 81.465 143.675 81.485 ;
        RECT 120.845 81.365 143.670 81.465 ;
        POLYGON 143.670 81.465 143.675 81.465 143.670 81.365 ;
        POLYGON 146.995 81.485 146.995 81.365 146.710 81.365 ;
        RECT 146.995 81.375 172.055 81.485 ;
        POLYGON 172.055 81.600 172.665 81.375 172.055 81.375 ;
        POLYGON 211.735 81.600 211.735 81.390 211.625 81.390 ;
        RECT 211.735 81.580 242.310 81.605 ;
        POLYGON 242.310 81.605 242.375 81.605 242.310 81.580 ;
        POLYGON 266.915 81.605 266.985 81.605 266.985 81.580 ;
        RECT 266.985 81.580 303.120 81.605 ;
        RECT 211.735 81.390 241.790 81.580 ;
        RECT 211.625 81.385 241.790 81.390 ;
        POLYGON 241.790 81.580 242.310 81.580 241.790 81.385 ;
        POLYGON 266.985 81.580 267.015 81.580 267.015 81.570 ;
        RECT 267.015 81.570 303.120 81.580 ;
        POLYGON 267.015 81.570 267.430 81.570 267.430 81.425 ;
        RECT 267.430 81.425 303.120 81.570 ;
        POLYGON 267.430 81.425 267.525 81.425 267.525 81.385 ;
        RECT 267.525 81.385 303.120 81.425 ;
        POLYGON 211.625 81.385 211.625 81.380 211.620 81.380 ;
        RECT 211.625 81.380 241.765 81.385 ;
        RECT 211.620 81.375 241.765 81.380 ;
        POLYGON 241.765 81.385 241.790 81.385 241.765 81.375 ;
        POLYGON 267.525 81.385 267.550 81.385 267.550 81.375 ;
        RECT 267.550 81.375 303.120 81.385 ;
        RECT 146.995 81.365 172.665 81.375 ;
        RECT 48.625 80.375 116.095 81.365 ;
        POLYGON 116.095 81.365 116.600 81.365 116.095 80.375 ;
        POLYGON 120.820 81.365 120.820 81.080 120.755 81.080 ;
        RECT 120.820 81.080 143.655 81.365 ;
        POLYGON 143.655 81.365 143.670 81.365 143.655 81.080 ;
        POLYGON 146.710 81.365 146.710 81.080 146.025 81.080 ;
        RECT 146.710 81.160 172.665 81.365 ;
        POLYGON 172.665 81.375 173.180 81.160 172.665 81.160 ;
        POLYGON 211.620 81.375 211.620 81.165 211.510 81.165 ;
        RECT 211.620 81.340 241.680 81.375 ;
        POLYGON 241.680 81.375 241.765 81.375 241.680 81.340 ;
        POLYGON 267.550 81.375 267.575 81.375 267.575 81.365 ;
        RECT 267.575 81.365 303.120 81.375 ;
        POLYGON 267.575 81.365 267.635 81.365 267.635 81.340 ;
        RECT 267.635 81.340 303.120 81.365 ;
        RECT 211.620 81.165 241.275 81.340 ;
        POLYGON 241.275 81.340 241.680 81.340 241.275 81.165 ;
        POLYGON 267.635 81.340 267.780 81.340 267.780 81.280 ;
        RECT 267.780 81.280 303.120 81.340 ;
        POLYGON 267.780 81.280 268.055 81.280 268.055 81.165 ;
        RECT 268.055 81.165 303.120 81.280 ;
        RECT 146.710 81.080 173.185 81.160 ;
        POLYGON 120.755 81.080 120.755 81.035 120.745 81.035 ;
        RECT 120.755 81.035 143.655 81.080 ;
        POLYGON 146.020 81.080 146.020 81.035 145.910 81.035 ;
        RECT 146.020 81.035 173.185 81.080 ;
        POLYGON 120.745 81.035 120.745 80.770 120.685 80.770 ;
        RECT 120.745 80.770 143.640 81.035 ;
        POLYGON 143.640 81.035 143.655 81.035 143.640 80.785 ;
        POLYGON 145.910 81.035 145.910 80.785 145.375 80.785 ;
        RECT 145.910 80.810 173.185 81.035 ;
        POLYGON 173.185 81.160 174.025 80.810 173.185 80.810 ;
        POLYGON 211.510 81.160 211.510 81.095 211.475 81.095 ;
        RECT 211.510 81.095 240.745 81.165 ;
        POLYGON 211.475 81.095 211.475 80.810 211.340 80.810 ;
        RECT 211.475 80.935 240.745 81.095 ;
        POLYGON 240.745 81.165 241.275 81.165 240.745 80.935 ;
        POLYGON 268.055 81.165 268.615 81.165 268.615 80.935 ;
        RECT 268.615 80.935 303.120 81.165 ;
        RECT 211.475 80.900 240.665 80.935 ;
        POLYGON 240.665 80.935 240.745 80.935 240.665 80.900 ;
        POLYGON 268.615 80.935 268.705 80.935 268.705 80.900 ;
        RECT 268.705 80.900 303.120 80.935 ;
        RECT 211.475 80.810 240.345 80.900 ;
        RECT 145.910 80.785 174.025 80.810 ;
        RECT 120.685 80.760 143.640 80.770 ;
        POLYGON 145.375 80.785 145.375 80.760 145.320 80.760 ;
        RECT 145.375 80.760 174.025 80.785 ;
        POLYGON 120.685 80.760 120.685 80.550 120.635 80.550 ;
        RECT 120.685 80.550 143.630 80.760 ;
        POLYGON 143.630 80.760 143.640 80.760 143.630 80.595 ;
        POLYGON 145.315 80.760 145.315 80.595 144.950 80.595 ;
        RECT 145.315 80.595 174.025 80.760 ;
        POLYGON 144.950 80.595 144.950 80.550 144.850 80.550 ;
        RECT 144.950 80.550 174.025 80.595 ;
        POLYGON 120.635 80.550 120.635 80.375 120.595 80.375 ;
        RECT 120.635 80.375 143.620 80.550 ;
        POLYGON 143.620 80.550 143.630 80.550 143.620 80.400 ;
        POLYGON 144.850 80.550 144.850 80.400 144.555 80.400 ;
        RECT 144.850 80.400 174.025 80.550 ;
        POLYGON 144.555 80.400 144.555 80.375 144.505 80.375 ;
        RECT 144.555 80.375 174.025 80.400 ;
        RECT 48.625 80.145 115.990 80.375 ;
        POLYGON 115.990 80.375 116.095 80.375 115.990 80.145 ;
        POLYGON 120.595 80.375 120.595 80.150 120.545 80.150 ;
        RECT 120.595 80.150 143.605 80.375 ;
        RECT 48.625 80.065 115.955 80.145 ;
        POLYGON 115.955 80.145 115.990 80.145 115.955 80.065 ;
        POLYGON 120.545 80.145 120.545 80.065 120.525 80.065 ;
        RECT 120.545 80.065 143.605 80.150 ;
        POLYGON 143.605 80.375 143.620 80.375 143.605 80.145 ;
        POLYGON 144.505 80.375 144.505 80.145 144.050 80.145 ;
        RECT 144.505 80.250 174.025 80.375 ;
        POLYGON 174.025 80.810 175.235 80.250 174.025 80.250 ;
        POLYGON 211.340 80.805 211.340 80.250 211.080 80.250 ;
        RECT 211.340 80.765 240.345 80.810 ;
        POLYGON 240.345 80.900 240.660 80.900 240.345 80.765 ;
        POLYGON 268.705 80.900 268.730 80.900 268.730 80.895 ;
        RECT 268.730 80.895 303.120 80.900 ;
        POLYGON 268.730 80.895 268.935 80.895 268.935 80.810 ;
        RECT 268.935 80.810 303.120 80.895 ;
        POLYGON 268.935 80.810 269.010 80.810 269.010 80.780 ;
        RECT 269.010 80.780 303.120 80.810 ;
        POLYGON 269.010 80.780 269.040 80.780 269.040 80.765 ;
        RECT 269.040 80.765 303.120 80.780 ;
        RECT 211.340 80.515 239.835 80.765 ;
        POLYGON 239.835 80.765 240.345 80.765 239.835 80.515 ;
        POLYGON 269.040 80.765 269.570 80.765 269.570 80.515 ;
        RECT 269.570 80.515 303.120 80.765 ;
        RECT 211.340 80.435 239.670 80.515 ;
        POLYGON 239.670 80.515 239.835 80.515 239.670 80.435 ;
        POLYGON 269.570 80.515 269.605 80.515 269.605 80.500 ;
        RECT 269.605 80.500 303.120 80.515 ;
        POLYGON 269.610 80.500 269.745 80.500 269.745 80.435 ;
        RECT 269.745 80.435 303.120 80.500 ;
        RECT 211.340 80.255 239.305 80.435 ;
        POLYGON 239.305 80.435 239.670 80.435 239.305 80.255 ;
        POLYGON 269.745 80.435 269.885 80.435 269.885 80.370 ;
        RECT 269.885 80.370 303.120 80.435 ;
        POLYGON 269.885 80.370 270.130 80.370 270.130 80.255 ;
        RECT 270.130 80.255 303.120 80.370 ;
        RECT 211.340 80.250 239.170 80.255 ;
        RECT 144.505 80.190 175.235 80.250 ;
        POLYGON 175.235 80.250 175.355 80.190 175.235 80.190 ;
        POLYGON 211.080 80.250 211.080 80.190 211.050 80.190 ;
        RECT 211.080 80.190 239.170 80.250 ;
        POLYGON 239.170 80.255 239.300 80.255 239.170 80.190 ;
        POLYGON 270.130 80.255 270.270 80.255 270.270 80.190 ;
        RECT 270.270 80.190 303.120 80.255 ;
        RECT 144.505 80.145 175.360 80.190 ;
        POLYGON 144.050 80.145 144.050 80.065 143.895 80.065 ;
        RECT 144.050 80.065 175.360 80.145 ;
        RECT 48.625 79.900 115.885 80.065 ;
        POLYGON 115.885 80.065 115.955 80.065 115.885 79.900 ;
        POLYGON 120.525 80.065 120.525 80.025 120.515 80.025 ;
        RECT 120.525 80.025 143.600 80.065 ;
        POLYGON 143.600 80.065 143.605 80.065 143.600 80.025 ;
        POLYGON 143.895 80.065 143.895 80.025 143.815 80.025 ;
        RECT 143.895 80.025 175.360 80.065 ;
        POLYGON 120.515 80.020 120.515 79.910 120.490 79.910 ;
        RECT 120.515 80.010 143.600 80.025 ;
        RECT 120.515 79.910 143.595 80.010 ;
        POLYGON 143.595 80.010 143.600 80.010 143.595 79.915 ;
        POLYGON 143.815 80.025 143.815 79.915 143.615 79.915 ;
        RECT 143.815 79.915 175.360 80.025 ;
        RECT 120.490 79.905 143.595 79.910 ;
        POLYGON 143.615 79.915 143.615 79.905 143.595 79.905 ;
        RECT 143.615 79.905 175.360 79.915 ;
        RECT 48.625 79.725 115.350 79.900 ;
        POLYGON 48.485 79.725 48.485 76.885 48.475 76.885 ;
        RECT 48.485 78.690 115.350 79.725 ;
        POLYGON 115.350 79.900 115.885 79.900 115.350 78.690 ;
        POLYGON 120.490 79.900 120.490 79.585 120.415 79.585 ;
        RECT 120.490 79.650 175.360 79.905 ;
        POLYGON 175.360 80.190 176.415 79.650 175.360 79.650 ;
        POLYGON 211.050 80.185 211.050 80.135 211.025 80.135 ;
        RECT 211.050 80.135 239.055 80.190 ;
        POLYGON 239.055 80.190 239.170 80.190 239.055 80.135 ;
        POLYGON 270.270 80.190 270.390 80.190 270.390 80.135 ;
        RECT 270.390 80.135 303.120 80.190 ;
        POLYGON 211.025 80.135 211.025 79.930 210.930 79.930 ;
        RECT 211.025 80.085 238.955 80.135 ;
        POLYGON 238.955 80.135 239.055 80.135 238.955 80.085 ;
        POLYGON 270.390 80.135 270.500 80.135 270.500 80.085 ;
        RECT 270.500 80.085 303.120 80.135 ;
        RECT 211.025 79.945 238.710 80.085 ;
        POLYGON 238.710 80.085 238.955 80.085 238.710 79.945 ;
        POLYGON 270.500 80.085 270.555 80.085 270.555 80.060 ;
        RECT 270.555 80.060 303.120 80.085 ;
        POLYGON 270.555 80.060 270.585 80.060 270.585 80.045 ;
        RECT 270.585 80.045 303.120 80.060 ;
        POLYGON 270.585 80.045 270.775 80.045 270.775 79.945 ;
        RECT 270.775 79.945 303.120 80.045 ;
        RECT 211.025 79.930 238.210 79.945 ;
        POLYGON 210.930 79.930 210.930 79.675 210.810 79.675 ;
        RECT 210.930 79.675 238.210 79.930 ;
        RECT 210.810 79.670 238.210 79.675 ;
        POLYGON 238.210 79.945 238.710 79.945 238.210 79.670 ;
        POLYGON 270.775 79.945 271.005 79.945 271.005 79.825 ;
        RECT 271.005 79.825 303.120 79.945 ;
        POLYGON 271.005 79.825 271.295 79.825 271.295 79.670 ;
        RECT 271.295 79.670 303.120 79.825 ;
        POLYGON 210.810 79.670 210.810 79.655 210.800 79.655 ;
        RECT 210.810 79.655 237.960 79.670 ;
        RECT 120.490 79.585 176.415 79.650 ;
        POLYGON 120.415 79.575 120.415 79.535 120.405 79.535 ;
        RECT 120.415 79.535 176.415 79.585 ;
        POLYGON 120.405 79.525 120.405 79.470 120.390 79.470 ;
        RECT 120.405 79.520 176.415 79.535 ;
        POLYGON 176.415 79.650 176.665 79.520 176.415 79.520 ;
        POLYGON 210.800 79.650 210.800 79.530 210.740 79.530 ;
        RECT 210.800 79.530 237.960 79.655 ;
        POLYGON 237.960 79.670 238.210 79.670 237.960 79.530 ;
        POLYGON 271.295 79.670 271.490 79.670 271.490 79.570 ;
        RECT 271.490 79.570 303.120 79.670 ;
        POLYGON 271.490 79.570 271.565 79.570 271.565 79.530 ;
        RECT 271.565 79.530 303.120 79.570 ;
        POLYGON 210.740 79.525 210.740 79.520 210.735 79.520 ;
        RECT 210.740 79.520 237.940 79.530 ;
        POLYGON 237.940 79.530 237.960 79.530 237.940 79.520 ;
        POLYGON 271.565 79.530 271.585 79.530 271.585 79.520 ;
        RECT 271.585 79.520 303.120 79.530 ;
        RECT 120.405 79.470 176.670 79.520 ;
        POLYGON 120.390 79.465 120.390 79.005 120.285 79.005 ;
        RECT 120.390 79.215 176.670 79.470 ;
        POLYGON 176.670 79.520 177.210 79.215 176.670 79.215 ;
        POLYGON 210.735 79.515 210.735 79.505 210.730 79.505 ;
        RECT 210.735 79.505 237.775 79.520 ;
        POLYGON 210.730 79.505 210.730 79.230 210.610 79.230 ;
        RECT 210.730 79.430 237.775 79.505 ;
        POLYGON 237.775 79.520 237.940 79.520 237.775 79.430 ;
        POLYGON 271.585 79.520 271.755 79.520 271.755 79.430 ;
        RECT 271.755 79.430 303.120 79.520 ;
        RECT 210.730 79.335 237.605 79.430 ;
        POLYGON 237.605 79.430 237.775 79.430 237.605 79.335 ;
        POLYGON 271.755 79.430 271.935 79.430 271.935 79.335 ;
        RECT 271.935 79.335 303.120 79.430 ;
        RECT 210.730 79.230 237.435 79.335 ;
        POLYGON 237.435 79.335 237.605 79.335 237.435 79.230 ;
        POLYGON 271.935 79.335 272.045 79.335 272.045 79.280 ;
        RECT 272.045 79.280 303.120 79.335 ;
        POLYGON 272.045 79.280 272.060 79.280 272.060 79.275 ;
        RECT 272.060 79.275 303.120 79.280 ;
        POLYGON 272.060 79.275 272.135 79.275 272.135 79.230 ;
        RECT 272.135 79.230 303.120 79.275 ;
        POLYGON 210.610 79.225 210.610 79.215 210.605 79.215 ;
        RECT 210.610 79.215 236.875 79.230 ;
        RECT 120.390 79.005 177.210 79.215 ;
        POLYGON 120.285 78.995 120.285 78.880 120.255 78.880 ;
        RECT 120.285 78.880 177.210 79.005 ;
        POLYGON 120.255 78.870 120.255 78.695 120.215 78.695 ;
        RECT 120.255 78.800 177.210 78.880 ;
        POLYGON 177.210 79.215 177.945 78.800 177.210 78.800 ;
        POLYGON 210.605 79.215 210.605 78.820 210.435 78.820 ;
        RECT 210.605 78.880 236.875 79.215 ;
        POLYGON 236.875 79.230 237.435 79.230 236.875 78.880 ;
        POLYGON 272.135 79.230 272.340 79.230 272.340 79.110 ;
        RECT 272.340 79.110 303.120 79.230 ;
        POLYGON 272.340 79.110 272.520 79.110 272.520 79.005 ;
        RECT 272.520 79.005 303.120 79.110 ;
        POLYGON 272.525 79.005 272.735 79.005 272.735 78.880 ;
        RECT 272.735 78.880 303.120 79.005 ;
        RECT 210.605 78.820 236.765 78.880 ;
        RECT 210.435 78.815 236.765 78.820 ;
        POLYGON 236.765 78.880 236.870 78.880 236.765 78.815 ;
        POLYGON 272.735 78.880 272.845 78.880 272.845 78.815 ;
        RECT 272.845 78.815 303.120 78.880 ;
        POLYGON 210.435 78.815 210.435 78.800 210.425 78.800 ;
        RECT 210.435 78.800 236.610 78.815 ;
        RECT 120.255 78.695 177.945 78.800 ;
        RECT 48.485 77.520 114.835 78.690 ;
        POLYGON 114.835 78.690 115.350 78.690 114.835 77.520 ;
        POLYGON 120.215 78.690 120.215 78.255 120.115 78.255 ;
        RECT 120.215 78.540 177.945 78.695 ;
        POLYGON 177.945 78.800 178.370 78.540 177.945 78.540 ;
        POLYGON 210.425 78.795 210.425 78.565 210.325 78.565 ;
        RECT 210.425 78.720 236.610 78.800 ;
        POLYGON 236.610 78.815 236.765 78.815 236.610 78.720 ;
        POLYGON 272.845 78.815 272.965 78.815 272.965 78.745 ;
        RECT 272.965 78.745 303.120 78.815 ;
        POLYGON 272.965 78.745 273.005 78.745 273.005 78.720 ;
        RECT 273.005 78.720 303.120 78.745 ;
        RECT 210.425 78.595 236.410 78.720 ;
        POLYGON 236.410 78.720 236.610 78.720 236.410 78.595 ;
        POLYGON 273.005 78.720 273.120 78.720 273.120 78.655 ;
        RECT 273.120 78.655 303.120 78.720 ;
        POLYGON 273.120 78.655 273.225 78.655 273.225 78.595 ;
        RECT 273.225 78.595 303.120 78.655 ;
        RECT 210.425 78.565 236.355 78.595 ;
        RECT 210.325 78.560 236.355 78.565 ;
        POLYGON 236.355 78.595 236.410 78.595 236.355 78.560 ;
        POLYGON 273.225 78.595 273.285 78.595 273.285 78.560 ;
        RECT 273.285 78.560 303.120 78.595 ;
        POLYGON 210.325 78.560 210.325 78.540 210.315 78.540 ;
        RECT 210.325 78.540 236.290 78.560 ;
        RECT 120.215 78.255 178.370 78.540 ;
        POLYGON 120.115 78.250 120.115 78.010 120.060 78.010 ;
        RECT 120.115 78.085 178.370 78.255 ;
        POLYGON 178.370 78.540 179.105 78.085 178.370 78.085 ;
        POLYGON 210.315 78.540 210.315 78.100 210.125 78.100 ;
        RECT 210.315 78.520 236.290 78.540 ;
        POLYGON 236.290 78.560 236.355 78.560 236.290 78.520 ;
        POLYGON 273.285 78.560 273.355 78.560 273.355 78.520 ;
        RECT 273.355 78.520 303.120 78.560 ;
        RECT 210.315 78.325 236.005 78.520 ;
        POLYGON 236.005 78.520 236.290 78.520 236.005 78.325 ;
        POLYGON 273.355 78.520 273.365 78.520 273.365 78.515 ;
        RECT 273.365 78.515 303.120 78.520 ;
        POLYGON 273.365 78.515 273.525 78.515 273.525 78.420 ;
        RECT 273.525 78.420 303.120 78.515 ;
        POLYGON 273.525 78.420 273.535 78.420 273.535 78.415 ;
        RECT 273.535 78.415 303.120 78.420 ;
        POLYGON 273.535 78.415 273.670 78.415 273.670 78.325 ;
        RECT 273.670 78.325 303.120 78.415 ;
        RECT 210.315 78.100 235.675 78.325 ;
        RECT 210.125 78.095 235.675 78.100 ;
        POLYGON 235.675 78.325 236.005 78.325 235.675 78.095 ;
        POLYGON 273.670 78.325 273.720 78.325 273.720 78.295 ;
        RECT 273.720 78.295 303.120 78.325 ;
        POLYGON 273.720 78.295 273.840 78.295 273.840 78.215 ;
        RECT 273.840 78.215 303.120 78.295 ;
        POLYGON 273.840 78.215 274.025 78.215 274.025 78.095 ;
        RECT 274.025 78.095 303.120 78.215 ;
        POLYGON 210.125 78.095 210.125 78.090 210.120 78.090 ;
        RECT 210.125 78.090 235.610 78.095 ;
        RECT 120.115 78.030 179.105 78.085 ;
        POLYGON 179.105 78.085 179.200 78.030 179.105 78.030 ;
        POLYGON 210.120 78.085 210.120 78.055 210.105 78.055 ;
        RECT 210.120 78.055 235.610 78.090 ;
        RECT 210.105 78.050 235.610 78.055 ;
        POLYGON 235.610 78.095 235.675 78.095 235.610 78.050 ;
        POLYGON 274.025 78.095 274.095 78.095 274.095 78.050 ;
        RECT 274.095 78.050 303.120 78.095 ;
        POLYGON 210.105 78.050 210.105 78.030 210.095 78.030 ;
        RECT 210.105 78.030 235.275 78.050 ;
        RECT 120.115 78.010 179.200 78.030 ;
        POLYGON 120.060 78.000 120.060 77.720 119.995 77.720 ;
        RECT 120.060 77.720 179.200 78.010 ;
        POLYGON 119.995 77.720 119.995 77.595 119.965 77.595 ;
        RECT 119.995 77.595 179.200 77.720 ;
        POLYGON 119.965 77.590 119.965 77.525 119.950 77.525 ;
        RECT 119.965 77.525 179.200 77.595 ;
        RECT 48.485 77.375 114.780 77.520 ;
        POLYGON 114.780 77.520 114.835 77.520 114.780 77.375 ;
        POLYGON 119.950 77.520 119.950 77.375 119.915 77.375 ;
        RECT 119.950 77.375 179.200 77.525 ;
        RECT 48.485 76.885 113.755 77.375 ;
        RECT 16.145 71.820 23.730 76.355 ;
        POLYGON 23.730 76.355 24.555 76.355 23.730 71.820 ;
        POLYGON 48.475 76.355 48.475 75.465 48.470 75.465 ;
        RECT 48.475 75.465 113.755 76.885 ;
        POLYGON 48.470 75.465 48.485 75.465 48.485 75.165 ;
        RECT 48.485 75.165 113.755 75.465 ;
        POLYGON 48.485 75.165 48.645 75.165 48.645 71.915 ;
        RECT 48.645 74.620 113.755 75.165 ;
        POLYGON 113.755 77.375 114.780 77.375 113.755 74.620 ;
        POLYGON 119.915 77.370 119.915 76.905 119.810 76.905 ;
        RECT 119.915 77.215 179.200 77.375 ;
        POLYGON 179.200 78.030 180.415 77.215 179.200 77.215 ;
        POLYGON 210.095 78.030 210.095 77.890 210.035 77.890 ;
        RECT 210.095 77.890 235.275 78.030 ;
        POLYGON 210.035 77.890 210.035 77.215 209.770 77.215 ;
        RECT 210.035 77.815 235.275 77.890 ;
        POLYGON 235.275 78.050 235.610 78.050 235.275 77.815 ;
        POLYGON 274.095 78.050 274.275 78.050 274.275 77.935 ;
        RECT 274.275 77.935 303.120 78.050 ;
        POLYGON 274.275 77.935 274.460 77.935 274.460 77.815 ;
        RECT 274.460 77.815 303.120 77.935 ;
        RECT 210.035 77.750 235.175 77.815 ;
        POLYGON 235.175 77.815 235.275 77.815 235.175 77.750 ;
        POLYGON 274.460 77.815 274.500 77.815 274.500 77.790 ;
        RECT 274.500 77.790 303.120 77.815 ;
        POLYGON 274.500 77.790 274.560 77.790 274.560 77.750 ;
        RECT 274.560 77.750 303.120 77.790 ;
        RECT 210.035 77.635 235.015 77.750 ;
        POLYGON 235.015 77.750 235.175 77.750 235.015 77.635 ;
        POLYGON 274.560 77.750 274.735 77.750 274.735 77.635 ;
        RECT 274.735 77.635 303.120 77.750 ;
        RECT 210.035 77.215 234.465 77.635 ;
        POLYGON 234.465 77.635 235.015 77.635 234.465 77.215 ;
        POLYGON 274.735 77.635 274.785 77.635 274.785 77.605 ;
        RECT 274.785 77.605 303.120 77.635 ;
        POLYGON 274.785 77.605 274.950 77.605 274.950 77.500 ;
        RECT 274.950 77.500 303.120 77.605 ;
        POLYGON 274.950 77.500 275.095 77.500 275.095 77.400 ;
        RECT 275.095 77.400 303.120 77.500 ;
        POLYGON 275.095 77.400 275.260 77.400 275.260 77.280 ;
        RECT 275.260 77.280 303.120 77.400 ;
        POLYGON 275.260 77.280 275.350 77.280 275.350 77.215 ;
        RECT 275.350 77.215 303.120 77.280 ;
        RECT 119.915 76.905 180.420 77.215 ;
        POLYGON 119.810 76.900 119.810 76.330 119.680 76.330 ;
        RECT 119.810 76.850 180.420 76.905 ;
        POLYGON 180.420 77.215 180.920 76.850 180.420 76.850 ;
        POLYGON 209.770 77.215 209.770 76.875 209.635 76.875 ;
        RECT 209.770 77.150 234.380 77.215 ;
        POLYGON 234.380 77.215 234.465 77.215 234.380 77.150 ;
        POLYGON 275.350 77.215 275.440 77.215 275.440 77.150 ;
        RECT 275.440 77.150 303.120 77.215 ;
        RECT 209.770 76.875 234.010 77.150 ;
        RECT 209.635 76.870 234.010 76.875 ;
        POLYGON 234.010 77.150 234.380 77.150 234.010 76.870 ;
        POLYGON 275.440 77.150 275.635 77.150 275.635 77.015 ;
        RECT 275.635 77.015 303.120 77.150 ;
        POLYGON 275.635 77.015 275.695 77.015 275.695 76.970 ;
        RECT 275.695 76.970 303.120 77.015 ;
        POLYGON 275.695 76.970 275.835 76.970 275.835 76.870 ;
        RECT 275.835 76.870 303.120 76.970 ;
        POLYGON 209.635 76.870 209.635 76.850 209.625 76.850 ;
        RECT 209.635 76.850 233.980 76.870 ;
        RECT 119.810 76.505 180.925 76.850 ;
        RECT 209.625 76.845 233.980 76.850 ;
        POLYGON 233.980 76.870 234.010 76.870 233.980 76.845 ;
        POLYGON 275.835 76.870 275.870 76.870 275.870 76.845 ;
        RECT 275.870 76.845 303.120 76.870 ;
        POLYGON 180.925 76.845 181.400 76.505 180.925 76.505 ;
        POLYGON 209.625 76.845 209.625 76.530 209.500 76.530 ;
        RECT 209.625 76.770 233.880 76.845 ;
        POLYGON 233.880 76.845 233.980 76.845 233.880 76.770 ;
        POLYGON 275.870 76.845 275.975 76.845 275.975 76.770 ;
        RECT 275.975 76.770 303.120 76.845 ;
        RECT 209.625 76.690 233.775 76.770 ;
        POLYGON 233.775 76.770 233.880 76.770 233.775 76.690 ;
        POLYGON 275.975 76.770 276.090 76.770 276.090 76.690 ;
        RECT 276.090 76.690 303.120 76.770 ;
        RECT 209.625 76.560 233.620 76.690 ;
        POLYGON 233.620 76.690 233.775 76.690 233.620 76.560 ;
        POLYGON 276.090 76.690 276.115 76.690 276.115 76.675 ;
        RECT 276.115 76.675 303.120 76.690 ;
        POLYGON 276.115 76.675 276.270 76.675 276.270 76.560 ;
        RECT 276.270 76.560 303.120 76.675 ;
        RECT 209.625 76.530 233.580 76.560 ;
        RECT 209.500 76.525 233.580 76.530 ;
        POLYGON 233.580 76.560 233.620 76.560 233.580 76.525 ;
        POLYGON 276.270 76.560 276.320 76.560 276.320 76.525 ;
        RECT 276.320 76.525 303.120 76.560 ;
        POLYGON 209.500 76.525 209.500 76.505 209.490 76.505 ;
        RECT 209.500 76.505 233.385 76.525 ;
        RECT 119.810 76.355 181.400 76.505 ;
        POLYGON 181.400 76.505 181.605 76.355 181.400 76.355 ;
        POLYGON 209.490 76.505 209.490 76.365 209.435 76.365 ;
        RECT 209.490 76.365 233.385 76.505 ;
        RECT 209.435 76.360 233.385 76.365 ;
        POLYGON 233.385 76.525 233.580 76.525 233.385 76.360 ;
        POLYGON 276.320 76.525 276.330 76.525 276.330 76.520 ;
        RECT 276.330 76.520 303.120 76.525 ;
        POLYGON 276.330 76.520 276.450 76.520 276.450 76.425 ;
        RECT 276.450 76.425 303.120 76.520 ;
        POLYGON 276.450 76.425 276.535 76.425 276.535 76.360 ;
        RECT 276.535 76.360 303.120 76.425 ;
        POLYGON 209.435 76.360 209.435 76.355 209.430 76.355 ;
        RECT 209.435 76.355 233.145 76.360 ;
        RECT 119.810 76.350 181.605 76.355 ;
        POLYGON 181.605 76.355 181.610 76.350 181.605 76.350 ;
        RECT 119.810 76.330 181.610 76.350 ;
        POLYGON 119.680 76.330 119.680 76.175 119.650 76.175 ;
        RECT 119.680 76.175 181.610 76.330 ;
        POLYGON 119.650 76.165 119.650 76.135 119.645 76.135 ;
        RECT 119.650 76.135 181.610 76.175 ;
        POLYGON 119.645 76.125 119.645 75.445 119.520 75.445 ;
        RECT 119.645 75.520 181.610 76.135 ;
        POLYGON 181.610 76.350 182.665 75.520 181.610 75.520 ;
        POLYGON 209.430 76.350 209.430 76.250 209.390 76.250 ;
        RECT 209.430 76.250 233.145 76.355 ;
        POLYGON 209.390 76.250 209.390 76.155 209.355 76.155 ;
        RECT 209.390 76.155 233.145 76.250 ;
        POLYGON 233.145 76.360 233.385 76.360 233.145 76.155 ;
        POLYGON 276.535 76.360 276.770 76.360 276.770 76.180 ;
        RECT 276.770 76.180 303.120 76.360 ;
        POLYGON 276.770 76.180 276.800 76.180 276.800 76.155 ;
        RECT 276.800 76.155 303.120 76.180 ;
        RECT 209.355 76.150 233.140 76.155 ;
        POLYGON 233.140 76.155 233.145 76.155 233.140 76.150 ;
        POLYGON 276.800 76.155 276.805 76.155 276.805 76.150 ;
        RECT 276.805 76.150 303.120 76.155 ;
        POLYGON 209.355 76.150 209.355 75.545 209.140 75.545 ;
        RECT 209.355 75.950 232.910 76.150 ;
        POLYGON 232.910 76.150 233.140 76.150 232.910 75.950 ;
        POLYGON 276.805 76.150 276.895 76.150 276.895 76.080 ;
        RECT 276.895 76.080 303.120 76.150 ;
        POLYGON 276.895 76.080 277.050 76.080 277.050 75.960 ;
        RECT 277.050 75.960 303.120 76.080 ;
        POLYGON 277.050 75.960 277.060 75.960 277.060 75.950 ;
        RECT 277.060 75.950 303.120 75.960 ;
        RECT 209.355 75.675 232.580 75.950 ;
        POLYGON 232.580 75.950 232.910 75.950 232.580 75.675 ;
        POLYGON 277.060 75.950 277.205 75.950 277.205 75.840 ;
        RECT 277.205 75.840 303.120 75.950 ;
        POLYGON 277.205 75.840 277.285 75.840 277.285 75.775 ;
        RECT 277.285 75.775 303.120 75.840 ;
        POLYGON 277.290 75.775 277.410 75.775 277.410 75.675 ;
        RECT 277.410 75.675 303.120 75.775 ;
        RECT 209.355 75.545 232.435 75.675 ;
        RECT 209.140 75.540 232.435 75.545 ;
        POLYGON 232.435 75.675 232.580 75.675 232.435 75.540 ;
        POLYGON 277.410 75.675 277.455 75.675 277.455 75.640 ;
        RECT 277.455 75.640 303.120 75.675 ;
        POLYGON 277.455 75.640 277.490 75.640 277.490 75.615 ;
        RECT 277.490 75.615 303.120 75.640 ;
        POLYGON 277.490 75.615 277.585 75.615 277.585 75.540 ;
        RECT 277.585 75.540 303.120 75.615 ;
        POLYGON 209.140 75.540 209.140 75.520 209.130 75.520 ;
        RECT 209.140 75.520 232.390 75.540 ;
        RECT 119.645 75.445 182.665 75.520 ;
        POLYGON 182.665 75.520 182.765 75.445 182.665 75.445 ;
        POLYGON 209.130 75.515 209.130 75.450 209.105 75.450 ;
        RECT 209.130 75.500 232.390 75.520 ;
        POLYGON 232.390 75.540 232.435 75.540 232.390 75.500 ;
        POLYGON 277.585 75.540 277.635 75.540 277.635 75.500 ;
        RECT 277.635 75.500 303.120 75.540 ;
        RECT 209.130 75.450 232.340 75.500 ;
        POLYGON 232.340 75.500 232.390 75.500 232.340 75.450 ;
        POLYGON 277.635 75.500 277.650 75.500 277.650 75.490 ;
        RECT 277.650 75.490 303.120 75.500 ;
        POLYGON 277.655 75.490 277.695 75.490 277.695 75.450 ;
        RECT 277.695 75.450 303.120 75.490 ;
        POLYGON 119.520 75.440 119.520 75.420 119.515 75.420 ;
        RECT 119.520 75.420 182.765 75.445 ;
        POLYGON 119.515 75.415 119.515 74.630 119.370 74.630 ;
        RECT 119.515 74.630 182.765 75.420 ;
        RECT 48.645 74.605 113.750 74.620 ;
        POLYGON 113.750 74.620 113.755 74.620 113.750 74.605 ;
        RECT 48.645 71.865 112.930 74.605 ;
        POLYGON 112.930 74.605 113.750 74.605 112.930 71.865 ;
        POLYGON 119.370 74.605 119.370 73.815 119.225 73.815 ;
        RECT 119.370 74.490 182.765 74.630 ;
        POLYGON 182.765 75.445 183.890 74.490 182.765 74.490 ;
        POLYGON 209.105 75.445 209.105 74.595 208.805 74.595 ;
        RECT 209.105 75.355 232.240 75.450 ;
        POLYGON 232.240 75.450 232.340 75.450 232.240 75.355 ;
        POLYGON 277.695 75.450 277.775 75.450 277.775 75.385 ;
        RECT 277.775 75.385 303.120 75.450 ;
        POLYGON 277.775 75.385 277.795 75.385 277.795 75.370 ;
        RECT 277.795 75.370 303.120 75.385 ;
        POLYGON 277.795 75.370 277.810 75.370 277.810 75.355 ;
        RECT 277.810 75.355 303.120 75.370 ;
        RECT 209.105 75.040 231.900 75.355 ;
        POLYGON 231.900 75.355 232.240 75.355 231.900 75.040 ;
        POLYGON 277.810 75.355 277.860 75.355 277.860 75.310 ;
        RECT 277.860 75.310 303.120 75.355 ;
        POLYGON 277.860 75.310 277.885 75.310 277.885 75.295 ;
        RECT 277.885 75.295 303.120 75.310 ;
        POLYGON 277.885 75.295 277.905 75.295 277.905 75.270 ;
        RECT 277.905 75.270 303.120 75.295 ;
        POLYGON 277.910 75.270 277.915 75.270 277.915 75.265 ;
        RECT 277.915 75.265 303.120 75.270 ;
        POLYGON 277.915 75.265 278.175 75.265 278.175 75.040 ;
        RECT 278.175 75.040 303.120 75.265 ;
        RECT 209.105 74.740 231.580 75.040 ;
        POLYGON 231.580 75.040 231.900 75.040 231.580 74.740 ;
        POLYGON 278.175 75.040 278.530 75.040 278.530 74.740 ;
        RECT 278.530 74.740 303.120 75.040 ;
        RECT 209.105 74.595 231.425 74.740 ;
        POLYGON 231.425 74.740 231.580 74.740 231.425 74.595 ;
        POLYGON 278.530 74.740 278.700 74.740 278.700 74.595 ;
        RECT 278.700 74.595 303.120 74.740 ;
        POLYGON 208.805 74.595 208.805 74.500 208.775 74.500 ;
        RECT 208.805 74.500 231.335 74.595 ;
        POLYGON 231.335 74.595 231.425 74.595 231.335 74.500 ;
        POLYGON 278.700 74.595 278.810 74.595 278.810 74.500 ;
        RECT 278.810 74.500 303.120 74.595 ;
        RECT 119.370 74.095 183.890 74.490 ;
        POLYGON 183.890 74.490 184.325 74.095 183.890 74.095 ;
        POLYGON 208.775 74.490 208.775 74.100 208.655 74.100 ;
        RECT 208.775 74.445 231.280 74.500 ;
        POLYGON 231.280 74.500 231.335 74.500 231.280 74.445 ;
        POLYGON 278.810 74.500 278.875 74.500 278.875 74.445 ;
        RECT 278.875 74.445 303.120 74.500 ;
        RECT 208.775 74.300 231.140 74.445 ;
        POLYGON 231.140 74.445 231.280 74.445 231.140 74.300 ;
        POLYGON 278.875 74.445 278.960 74.445 278.960 74.375 ;
        RECT 278.960 74.375 303.120 74.445 ;
        POLYGON 278.960 74.375 279.040 74.375 279.040 74.300 ;
        RECT 279.040 74.300 303.120 74.375 ;
        RECT 208.775 74.155 231.005 74.300 ;
        POLYGON 231.005 74.300 231.140 74.300 231.005 74.155 ;
        POLYGON 279.040 74.300 279.195 74.300 279.195 74.155 ;
        RECT 279.195 74.155 303.120 74.300 ;
        RECT 208.775 74.100 230.950 74.155 ;
        POLYGON 230.950 74.155 231.005 74.155 230.950 74.100 ;
        POLYGON 279.195 74.155 279.255 74.155 279.255 74.100 ;
        RECT 279.255 74.100 303.120 74.155 ;
        RECT 119.370 74.085 184.325 74.095 ;
        POLYGON 184.325 74.095 184.335 74.085 184.325 74.085 ;
        RECT 119.370 73.945 184.335 74.085 ;
        POLYGON 208.655 74.095 208.655 74.080 208.650 74.080 ;
        RECT 208.655 74.080 230.745 74.100 ;
        RECT 119.370 73.940 156.975 73.945 ;
        POLYGON 156.975 73.945 157.285 73.945 156.975 73.940 ;
        POLYGON 157.710 73.945 157.885 73.945 157.885 73.940 ;
        RECT 157.885 73.940 184.335 73.945 ;
        RECT 119.370 73.935 156.650 73.940 ;
        POLYGON 156.650 73.940 156.970 73.940 156.650 73.935 ;
        POLYGON 157.885 73.940 158.065 73.940 158.065 73.935 ;
        RECT 158.065 73.935 184.335 73.940 ;
        RECT 119.370 73.925 156.410 73.935 ;
        POLYGON 156.410 73.935 156.650 73.935 156.410 73.925 ;
        POLYGON 158.065 73.935 158.245 73.935 158.245 73.930 ;
        RECT 158.245 73.930 184.335 73.935 ;
        POLYGON 158.245 73.930 158.415 73.930 158.415 73.925 ;
        RECT 158.415 73.925 184.335 73.930 ;
        RECT 119.370 73.900 155.855 73.925 ;
        POLYGON 155.855 73.925 156.400 73.925 155.855 73.900 ;
        POLYGON 158.435 73.925 158.720 73.925 158.720 73.905 ;
        RECT 158.720 73.905 184.335 73.925 ;
        POLYGON 158.740 73.905 158.840 73.905 158.840 73.900 ;
        RECT 158.840 73.900 184.335 73.905 ;
        RECT 119.370 73.880 155.615 73.900 ;
        POLYGON 155.615 73.900 155.855 73.900 155.615 73.880 ;
        POLYGON 158.840 73.900 159.045 73.900 159.045 73.890 ;
        RECT 159.045 73.890 184.335 73.900 ;
        POLYGON 159.075 73.890 159.135 73.890 159.135 73.880 ;
        RECT 159.135 73.880 184.335 73.890 ;
        RECT 119.370 73.875 155.505 73.880 ;
        POLYGON 155.505 73.880 155.610 73.880 155.505 73.875 ;
        POLYGON 159.145 73.880 159.200 73.880 159.200 73.875 ;
        RECT 159.200 73.875 184.335 73.880 ;
        RECT 119.370 73.855 155.285 73.875 ;
        POLYGON 155.285 73.875 155.500 73.875 155.285 73.855 ;
        POLYGON 159.200 73.875 159.430 73.875 159.430 73.855 ;
        RECT 159.430 73.855 184.335 73.875 ;
        RECT 119.370 73.840 155.065 73.855 ;
        POLYGON 155.065 73.855 155.285 73.855 155.065 73.840 ;
        POLYGON 159.430 73.855 159.605 73.855 159.605 73.840 ;
        RECT 159.605 73.840 184.335 73.855 ;
        RECT 119.370 73.815 154.775 73.840 ;
        RECT 119.225 73.810 154.775 73.815 ;
        POLYGON 154.775 73.840 155.065 73.840 154.775 73.810 ;
        POLYGON 159.605 73.840 159.840 73.840 159.840 73.820 ;
        RECT 159.840 73.820 184.335 73.840 ;
        POLYGON 159.865 73.820 159.945 73.820 159.945 73.810 ;
        RECT 159.945 73.810 184.335 73.820 ;
        POLYGON 119.225 73.805 119.225 73.040 119.085 73.040 ;
        RECT 119.225 73.755 154.275 73.810 ;
        POLYGON 154.275 73.810 154.770 73.810 154.275 73.755 ;
        POLYGON 159.945 73.810 160.395 73.810 160.395 73.755 ;
        RECT 160.395 73.755 184.335 73.810 ;
        RECT 119.225 73.730 154.120 73.755 ;
        POLYGON 154.120 73.755 154.275 73.755 154.120 73.730 ;
        POLYGON 160.395 73.755 160.520 73.755 160.520 73.740 ;
        RECT 160.520 73.740 184.335 73.755 ;
        POLYGON 160.520 73.740 160.595 73.740 160.595 73.730 ;
        RECT 160.595 73.730 184.335 73.740 ;
        RECT 119.225 73.725 154.070 73.730 ;
        POLYGON 154.070 73.730 154.120 73.730 154.070 73.725 ;
        POLYGON 160.595 73.730 160.635 73.730 160.635 73.725 ;
        RECT 160.635 73.725 184.335 73.730 ;
        RECT 119.225 73.720 154.050 73.725 ;
        POLYGON 154.050 73.725 154.070 73.725 154.050 73.720 ;
        POLYGON 160.635 73.725 160.670 73.725 160.670 73.720 ;
        RECT 160.670 73.720 184.335 73.725 ;
        RECT 119.225 73.640 153.490 73.720 ;
        POLYGON 153.490 73.720 154.045 73.720 153.490 73.640 ;
        POLYGON 160.670 73.720 160.845 73.720 160.845 73.695 ;
        RECT 160.845 73.695 184.335 73.720 ;
        POLYGON 160.850 73.695 160.970 73.695 160.970 73.675 ;
        RECT 160.970 73.675 184.335 73.695 ;
        POLYGON 160.970 73.675 161.175 73.675 161.175 73.645 ;
        RECT 161.175 73.645 184.335 73.675 ;
        POLYGON 161.175 73.645 161.205 73.645 161.205 73.640 ;
        RECT 161.205 73.640 184.335 73.645 ;
        RECT 119.225 73.615 153.335 73.640 ;
        POLYGON 153.335 73.640 153.490 73.640 153.335 73.615 ;
        POLYGON 161.205 73.640 161.365 73.640 161.365 73.615 ;
        RECT 161.365 73.615 184.335 73.640 ;
        RECT 119.225 73.550 152.955 73.615 ;
        POLYGON 152.955 73.615 153.335 73.615 152.955 73.550 ;
        POLYGON 161.365 73.615 161.430 73.615 161.430 73.605 ;
        RECT 161.430 73.605 184.335 73.615 ;
        POLYGON 161.430 73.605 161.720 73.605 161.720 73.550 ;
        RECT 161.720 73.550 184.335 73.605 ;
        RECT 119.225 73.510 152.745 73.550 ;
        POLYGON 152.745 73.550 152.950 73.550 152.745 73.510 ;
        POLYGON 161.720 73.550 161.800 73.550 161.800 73.535 ;
        RECT 161.800 73.535 184.335 73.550 ;
        POLYGON 161.805 73.535 161.940 73.535 161.940 73.510 ;
        RECT 161.940 73.510 184.335 73.535 ;
        RECT 119.225 73.505 152.710 73.510 ;
        POLYGON 152.710 73.510 152.745 73.510 152.710 73.505 ;
        POLYGON 161.940 73.510 161.965 73.510 161.965 73.505 ;
        RECT 161.965 73.505 184.335 73.510 ;
        RECT 119.225 73.490 152.645 73.505 ;
        POLYGON 152.645 73.505 152.710 73.505 152.645 73.490 ;
        POLYGON 161.965 73.505 162.050 73.505 162.050 73.490 ;
        RECT 162.050 73.495 184.335 73.505 ;
        POLYGON 184.335 74.080 184.980 73.495 184.335 73.495 ;
        POLYGON 208.650 74.075 208.650 73.525 208.485 73.525 ;
        RECT 208.650 73.890 230.745 74.080 ;
        POLYGON 230.745 74.100 230.950 74.100 230.745 73.890 ;
        POLYGON 279.255 74.100 279.440 74.100 279.440 73.925 ;
        RECT 279.440 73.925 303.120 74.100 ;
        POLYGON 251.650 73.925 251.650 73.900 251.105 73.900 ;
        RECT 251.650 73.900 252.820 73.925 ;
        POLYGON 252.820 73.925 253.370 73.900 252.820 73.900 ;
        POLYGON 279.440 73.925 279.465 73.925 279.465 73.900 ;
        RECT 279.465 73.900 303.120 73.925 ;
        POLYGON 251.105 73.900 251.105 73.890 250.980 73.890 ;
        RECT 251.105 73.895 253.380 73.900 ;
        POLYGON 253.380 73.900 253.395 73.895 253.380 73.895 ;
        POLYGON 279.465 73.900 279.475 73.900 279.475 73.895 ;
        RECT 279.475 73.895 303.120 73.900 ;
        RECT 251.105 73.890 253.405 73.895 ;
        RECT 208.650 73.640 230.505 73.890 ;
        POLYGON 230.505 73.890 230.745 73.890 230.505 73.640 ;
        POLYGON 250.945 73.890 250.945 73.870 250.495 73.870 ;
        RECT 250.945 73.870 253.405 73.890 ;
        POLYGON 253.405 73.895 253.970 73.870 253.405 73.870 ;
        POLYGON 279.475 73.895 279.500 73.895 279.500 73.870 ;
        RECT 279.500 73.870 303.120 73.895 ;
        POLYGON 250.495 73.870 250.495 73.840 250.200 73.840 ;
        RECT 250.495 73.845 253.990 73.870 ;
        POLYGON 253.990 73.870 254.220 73.845 253.990 73.845 ;
        POLYGON 279.500 73.870 279.525 73.870 279.525 73.845 ;
        RECT 279.525 73.845 303.120 73.870 ;
        RECT 250.495 73.840 254.220 73.845 ;
        POLYGON 254.220 73.845 254.285 73.840 254.220 73.840 ;
        POLYGON 279.525 73.845 279.530 73.845 279.530 73.840 ;
        RECT 279.530 73.840 303.120 73.845 ;
        POLYGON 250.195 73.840 250.195 73.760 249.345 73.760 ;
        RECT 250.195 73.805 254.290 73.840 ;
        POLYGON 254.290 73.840 254.665 73.805 254.290 73.805 ;
        POLYGON 279.530 73.840 279.570 73.840 279.570 73.805 ;
        RECT 279.570 73.805 303.120 73.840 ;
        RECT 250.195 73.760 254.670 73.805 ;
        POLYGON 254.670 73.805 255.160 73.760 254.670 73.760 ;
        POLYGON 279.570 73.805 279.620 73.805 279.620 73.760 ;
        RECT 279.620 73.760 303.120 73.805 ;
        POLYGON 249.345 73.760 249.345 73.640 248.530 73.640 ;
        RECT 249.345 73.660 255.160 73.760 ;
        POLYGON 255.160 73.760 255.830 73.660 255.160 73.660 ;
        POLYGON 279.620 73.760 279.725 73.760 279.725 73.660 ;
        RECT 279.725 73.660 303.120 73.760 ;
        RECT 249.345 73.650 255.830 73.660 ;
        POLYGON 255.830 73.660 255.905 73.650 255.830 73.650 ;
        POLYGON 279.725 73.660 279.735 73.660 279.735 73.650 ;
        RECT 279.735 73.650 303.120 73.660 ;
        RECT 249.345 73.640 255.905 73.650 ;
        RECT 208.650 73.525 230.390 73.640 ;
        RECT 208.485 73.520 230.390 73.525 ;
        POLYGON 230.390 73.640 230.505 73.640 230.390 73.520 ;
        POLYGON 248.530 73.640 248.530 73.635 248.495 73.635 ;
        RECT 248.530 73.635 255.905 73.640 ;
        POLYGON 248.490 73.635 248.490 73.595 248.205 73.595 ;
        RECT 248.490 73.595 255.905 73.635 ;
        POLYGON 248.205 73.595 248.205 73.520 247.820 73.520 ;
        RECT 248.205 73.590 255.905 73.595 ;
        POLYGON 255.905 73.650 256.330 73.590 255.905 73.590 ;
        POLYGON 279.735 73.650 279.800 73.650 279.800 73.590 ;
        RECT 279.800 73.590 303.120 73.650 ;
        RECT 248.205 73.520 256.330 73.590 ;
        POLYGON 256.330 73.590 256.690 73.520 256.330 73.520 ;
        POLYGON 279.800 73.590 279.875 73.590 279.875 73.520 ;
        RECT 279.875 73.520 303.120 73.590 ;
        POLYGON 208.485 73.520 208.485 73.495 208.475 73.495 ;
        RECT 208.485 73.495 230.285 73.520 ;
        RECT 162.050 73.490 184.980 73.495 ;
        RECT 119.225 73.350 151.970 73.490 ;
        POLYGON 151.970 73.490 152.640 73.490 151.970 73.350 ;
        POLYGON 162.050 73.490 162.220 73.490 162.220 73.455 ;
        RECT 162.220 73.455 184.980 73.490 ;
        POLYGON 162.220 73.455 162.565 73.455 162.565 73.380 ;
        RECT 162.565 73.380 184.980 73.455 ;
        POLYGON 162.565 73.380 162.695 73.380 162.695 73.350 ;
        RECT 162.695 73.350 184.980 73.380 ;
        RECT 119.225 73.345 151.940 73.350 ;
        POLYGON 151.940 73.350 151.965 73.350 151.940 73.345 ;
        POLYGON 162.695 73.350 162.715 73.350 162.715 73.345 ;
        RECT 162.715 73.345 184.980 73.350 ;
        RECT 119.225 73.310 151.790 73.345 ;
        POLYGON 151.790 73.345 151.940 73.345 151.790 73.310 ;
        POLYGON 162.715 73.345 162.870 73.345 162.870 73.310 ;
        RECT 162.870 73.310 184.980 73.345 ;
        RECT 119.225 73.255 151.550 73.310 ;
        POLYGON 151.550 73.310 151.790 73.310 151.550 73.255 ;
        POLYGON 162.870 73.310 162.915 73.310 162.915 73.300 ;
        RECT 162.915 73.300 184.980 73.310 ;
        POLYGON 162.920 73.300 163.105 73.300 163.105 73.260 ;
        RECT 163.105 73.260 184.980 73.300 ;
        POLYGON 163.105 73.260 163.125 73.260 163.125 73.255 ;
        RECT 163.125 73.255 184.980 73.260 ;
        RECT 119.225 73.195 151.320 73.255 ;
        POLYGON 151.320 73.255 151.550 73.255 151.320 73.195 ;
        POLYGON 163.125 73.255 163.145 73.255 163.145 73.250 ;
        RECT 163.145 73.250 184.980 73.255 ;
        POLYGON 163.145 73.250 163.355 73.250 163.355 73.195 ;
        RECT 163.355 73.195 184.980 73.250 ;
        RECT 119.225 73.160 151.170 73.195 ;
        POLYGON 151.170 73.195 151.320 73.195 151.170 73.160 ;
        POLYGON 163.355 73.195 163.490 73.195 163.490 73.160 ;
        RECT 163.490 73.160 184.980 73.195 ;
        RECT 119.225 73.040 150.700 73.160 ;
        POLYGON 119.085 73.035 119.085 72.665 119.015 72.665 ;
        RECT 119.085 73.030 150.700 73.040 ;
        POLYGON 150.700 73.160 151.170 73.160 150.700 73.030 ;
        POLYGON 163.490 73.160 163.995 73.160 163.995 73.030 ;
        RECT 163.995 73.030 184.980 73.160 ;
        RECT 119.085 73.015 150.635 73.030 ;
        POLYGON 150.635 73.030 150.695 73.030 150.635 73.015 ;
        POLYGON 164.000 73.030 164.050 73.030 164.050 73.015 ;
        RECT 164.050 73.015 184.980 73.030 ;
        RECT 119.085 72.955 150.415 73.015 ;
        POLYGON 150.415 73.015 150.630 73.015 150.415 72.955 ;
        POLYGON 164.050 73.015 164.125 73.015 164.125 72.990 ;
        RECT 164.125 72.990 184.980 73.015 ;
        POLYGON 164.125 72.990 164.145 72.990 164.145 72.985 ;
        RECT 164.145 72.985 184.980 72.990 ;
        POLYGON 164.145 72.985 164.245 72.985 164.245 72.955 ;
        RECT 164.245 72.955 184.980 72.985 ;
        RECT 119.085 72.945 150.380 72.955 ;
        POLYGON 150.380 72.955 150.415 72.955 150.380 72.945 ;
        POLYGON 164.245 72.955 164.275 72.955 164.275 72.945 ;
        RECT 164.275 72.945 184.980 72.955 ;
        RECT 119.085 72.750 149.750 72.945 ;
        POLYGON 149.750 72.945 150.380 72.945 149.750 72.750 ;
        POLYGON 164.275 72.945 164.930 72.945 164.930 72.750 ;
        RECT 164.930 72.750 184.980 72.945 ;
        RECT 119.085 72.725 149.665 72.750 ;
        POLYGON 149.665 72.750 149.745 72.750 149.665 72.725 ;
        POLYGON 164.930 72.750 165.005 72.750 165.005 72.725 ;
        RECT 165.005 72.725 184.980 72.750 ;
        RECT 119.085 72.665 149.485 72.725 ;
        RECT 119.015 72.660 149.485 72.665 ;
        POLYGON 149.485 72.725 149.665 72.725 149.485 72.660 ;
        POLYGON 165.005 72.725 165.040 72.725 165.040 72.715 ;
        RECT 165.040 72.715 184.980 72.725 ;
        POLYGON 165.045 72.715 165.115 72.715 165.115 72.690 ;
        RECT 165.115 72.690 184.980 72.715 ;
        POLYGON 165.115 72.690 165.205 72.690 165.205 72.660 ;
        RECT 165.205 72.660 184.980 72.690 ;
        POLYGON 119.015 72.655 119.015 71.865 118.870 71.865 ;
        RECT 119.015 72.575 149.230 72.660 ;
        POLYGON 149.230 72.660 149.485 72.660 149.230 72.575 ;
        POLYGON 165.205 72.660 165.460 72.660 165.460 72.575 ;
        RECT 165.460 72.590 184.980 72.660 ;
        POLYGON 184.980 73.495 185.900 72.590 184.980 72.590 ;
        POLYGON 208.475 73.490 208.475 73.225 208.395 73.225 ;
        RECT 208.475 73.410 230.285 73.495 ;
        POLYGON 230.285 73.520 230.390 73.520 230.285 73.410 ;
        POLYGON 247.820 73.520 247.820 73.510 247.770 73.510 ;
        RECT 247.820 73.510 256.690 73.520 ;
        POLYGON 247.770 73.510 247.770 73.410 247.235 73.410 ;
        RECT 247.770 73.440 256.690 73.510 ;
        POLYGON 256.690 73.520 257.110 73.440 256.690 73.440 ;
        POLYGON 279.875 73.520 279.960 73.520 279.960 73.440 ;
        RECT 279.960 73.440 303.120 73.520 ;
        RECT 247.770 73.410 257.115 73.440 ;
        RECT 208.475 73.225 230.085 73.410 ;
        POLYGON 208.395 73.225 208.395 72.600 208.205 72.600 ;
        RECT 208.395 73.205 230.085 73.225 ;
        POLYGON 230.085 73.410 230.285 73.410 230.085 73.205 ;
        POLYGON 247.235 73.410 247.235 73.390 247.125 73.390 ;
        RECT 247.235 73.395 257.115 73.410 ;
        POLYGON 257.115 73.440 257.335 73.395 257.115 73.395 ;
        POLYGON 279.960 73.440 280.010 73.440 280.010 73.395 ;
        RECT 280.010 73.395 303.120 73.440 ;
        RECT 247.235 73.390 257.340 73.395 ;
        POLYGON 247.120 73.390 247.120 73.380 247.075 73.380 ;
        RECT 247.120 73.380 257.340 73.390 ;
        POLYGON 247.075 73.380 247.075 73.260 246.585 73.260 ;
        RECT 247.075 73.365 257.340 73.380 ;
        POLYGON 257.340 73.395 257.495 73.365 257.340 73.365 ;
        POLYGON 280.010 73.395 280.040 73.395 280.040 73.365 ;
        RECT 280.040 73.365 303.120 73.395 ;
        RECT 247.075 73.330 257.495 73.365 ;
        POLYGON 257.495 73.365 257.655 73.330 257.495 73.330 ;
        POLYGON 280.040 73.365 280.080 73.365 280.080 73.330 ;
        RECT 280.080 73.330 303.120 73.365 ;
        RECT 247.075 73.260 257.660 73.330 ;
        POLYGON 246.585 73.260 246.585 73.205 246.360 73.205 ;
        RECT 246.585 73.205 257.660 73.260 ;
        RECT 208.395 73.145 230.025 73.205 ;
        POLYGON 230.025 73.205 230.085 73.205 230.025 73.145 ;
        POLYGON 246.360 73.205 246.360 73.170 246.220 73.170 ;
        RECT 246.360 73.175 257.660 73.205 ;
        POLYGON 257.660 73.330 258.295 73.175 257.660 73.175 ;
        POLYGON 280.080 73.330 280.205 73.330 280.205 73.215 ;
        RECT 280.205 73.215 303.120 73.330 ;
        POLYGON 280.205 73.215 280.240 73.215 280.240 73.175 ;
        RECT 280.240 73.175 303.120 73.215 ;
        RECT 246.360 73.170 258.295 73.175 ;
        POLYGON 246.220 73.170 246.220 73.145 246.110 73.145 ;
        RECT 246.220 73.145 258.295 73.170 ;
        RECT 208.395 73.025 229.910 73.145 ;
        POLYGON 229.910 73.145 230.025 73.145 229.910 73.025 ;
        POLYGON 246.110 73.145 246.110 73.110 245.960 73.110 ;
        RECT 246.110 73.110 258.295 73.145 ;
        POLYGON 245.960 73.110 245.960 73.025 245.670 73.025 ;
        RECT 245.960 73.085 258.295 73.110 ;
        POLYGON 258.295 73.175 258.660 73.085 258.295 73.085 ;
        POLYGON 280.240 73.175 280.330 73.175 280.330 73.085 ;
        RECT 280.330 73.085 303.120 73.175 ;
        RECT 245.960 73.050 258.660 73.085 ;
        POLYGON 258.660 73.085 258.775 73.050 258.660 73.050 ;
        POLYGON 280.330 73.085 280.365 73.085 280.365 73.050 ;
        RECT 280.365 73.050 303.120 73.085 ;
        RECT 245.960 73.025 258.775 73.050 ;
        RECT 208.395 73.010 229.895 73.025 ;
        POLYGON 229.895 73.025 229.910 73.025 229.895 73.010 ;
        POLYGON 245.670 73.025 245.670 73.010 245.620 73.010 ;
        RECT 245.670 73.010 258.775 73.025 ;
        RECT 208.395 72.835 229.745 73.010 ;
        POLYGON 229.745 73.010 229.895 73.010 229.745 72.835 ;
        POLYGON 245.620 73.010 245.620 72.835 245.030 72.835 ;
        RECT 245.620 72.855 258.775 73.010 ;
        POLYGON 258.775 73.050 259.450 72.855 258.775 72.855 ;
        POLYGON 280.365 73.050 280.560 73.050 280.560 72.855 ;
        RECT 280.560 72.855 303.120 73.050 ;
        RECT 245.620 72.835 259.455 72.855 ;
        RECT 208.395 72.600 229.545 72.835 ;
        POLYGON 229.545 72.835 229.745 72.835 229.545 72.600 ;
        POLYGON 245.030 72.835 245.030 72.785 244.860 72.785 ;
        RECT 245.030 72.785 259.455 72.835 ;
        POLYGON 244.860 72.785 244.860 72.730 244.705 72.730 ;
        RECT 244.860 72.745 259.455 72.785 ;
        POLYGON 259.455 72.855 259.820 72.745 259.455 72.745 ;
        POLYGON 280.560 72.855 280.670 72.855 280.670 72.745 ;
        RECT 280.670 72.745 303.120 72.855 ;
        RECT 244.860 72.730 259.820 72.745 ;
        POLYGON 244.705 72.730 244.705 72.600 244.330 72.600 ;
        RECT 244.705 72.630 259.820 72.730 ;
        POLYGON 259.820 72.745 260.165 72.630 259.820 72.630 ;
        POLYGON 280.670 72.745 280.785 72.745 280.785 72.630 ;
        RECT 280.785 72.630 303.120 72.745 ;
        RECT 244.705 72.600 260.165 72.630 ;
        POLYGON 260.165 72.630 260.250 72.600 260.165 72.600 ;
        POLYGON 280.785 72.630 280.810 72.630 280.810 72.600 ;
        RECT 280.810 72.600 303.120 72.630 ;
        RECT 165.460 72.575 185.900 72.590 ;
        RECT 119.015 72.470 148.920 72.575 ;
        POLYGON 148.920 72.575 149.230 72.575 148.920 72.470 ;
        POLYGON 165.460 72.575 165.520 72.575 165.520 72.555 ;
        RECT 165.520 72.555 185.900 72.575 ;
        POLYGON 165.525 72.555 165.575 72.555 165.575 72.535 ;
        RECT 165.575 72.535 185.900 72.555 ;
        POLYGON 165.575 72.535 165.760 72.535 165.760 72.470 ;
        RECT 165.760 72.470 185.900 72.535 ;
        RECT 119.015 72.435 148.830 72.470 ;
        POLYGON 148.830 72.470 148.920 72.470 148.830 72.435 ;
        POLYGON 165.760 72.470 165.790 72.470 165.790 72.460 ;
        RECT 165.790 72.460 185.900 72.470 ;
        POLYGON 165.790 72.460 165.855 72.460 165.855 72.435 ;
        RECT 165.855 72.455 185.900 72.460 ;
        POLYGON 185.900 72.590 186.035 72.455 185.900 72.455 ;
        POLYGON 208.205 72.590 208.205 72.475 208.170 72.475 ;
        RECT 208.205 72.530 229.485 72.600 ;
        POLYGON 229.485 72.600 229.545 72.600 229.485 72.530 ;
        POLYGON 244.330 72.600 244.330 72.530 244.125 72.530 ;
        RECT 244.330 72.530 260.250 72.600 ;
        RECT 208.205 72.475 229.440 72.530 ;
        POLYGON 229.440 72.530 229.485 72.530 229.440 72.480 ;
        POLYGON 244.125 72.530 244.125 72.500 244.040 72.500 ;
        RECT 244.125 72.500 260.250 72.530 ;
        POLYGON 244.040 72.500 244.040 72.480 243.980 72.480 ;
        RECT 244.040 72.485 260.250 72.500 ;
        POLYGON 260.250 72.600 260.585 72.485 260.250 72.485 ;
        POLYGON 280.810 72.600 280.925 72.600 280.925 72.485 ;
        RECT 280.925 72.485 303.120 72.600 ;
        RECT 244.040 72.480 260.585 72.485 ;
        POLYGON 243.980 72.480 243.980 72.475 243.970 72.475 ;
        RECT 243.980 72.475 260.585 72.480 ;
        POLYGON 260.585 72.485 260.610 72.475 260.585 72.475 ;
        POLYGON 280.925 72.485 280.935 72.485 280.935 72.475 ;
        RECT 280.935 72.475 303.120 72.485 ;
        POLYGON 208.170 72.475 208.170 72.460 208.165 72.460 ;
        RECT 208.170 72.460 229.305 72.475 ;
        RECT 165.855 72.435 186.035 72.455 ;
        RECT 119.015 72.255 148.355 72.435 ;
        POLYGON 148.355 72.435 148.830 72.435 148.355 72.255 ;
        POLYGON 165.855 72.435 166.050 72.435 166.050 72.365 ;
        RECT 166.050 72.365 186.035 72.435 ;
        POLYGON 166.050 72.365 166.070 72.365 166.070 72.355 ;
        RECT 166.070 72.355 186.035 72.365 ;
        POLYGON 166.070 72.355 166.335 72.355 166.335 72.255 ;
        RECT 166.335 72.255 186.035 72.355 ;
        RECT 119.015 72.190 148.190 72.255 ;
        POLYGON 148.190 72.255 148.355 72.255 148.190 72.190 ;
        POLYGON 166.335 72.255 166.510 72.255 166.510 72.190 ;
        RECT 166.510 72.190 186.035 72.255 ;
        RECT 119.015 72.155 148.100 72.190 ;
        POLYGON 148.100 72.190 148.190 72.190 148.100 72.155 ;
        POLYGON 166.510 72.190 166.595 72.190 166.595 72.160 ;
        RECT 166.595 72.160 186.035 72.190 ;
        POLYGON 166.595 72.160 166.605 72.160 166.605 72.155 ;
        RECT 166.605 72.155 186.035 72.160 ;
        RECT 119.015 72.090 147.945 72.155 ;
        POLYGON 147.945 72.155 148.100 72.155 147.945 72.090 ;
        POLYGON 166.605 72.155 166.630 72.155 166.630 72.145 ;
        RECT 166.630 72.145 186.035 72.155 ;
        POLYGON 166.630 72.145 166.755 72.145 166.755 72.090 ;
        RECT 166.755 72.090 186.035 72.145 ;
        RECT 119.015 71.890 147.470 72.090 ;
        POLYGON 147.470 72.090 147.945 72.090 147.470 71.890 ;
        POLYGON 166.755 72.090 166.995 72.090 166.995 71.990 ;
        RECT 166.995 71.990 186.035 72.090 ;
        POLYGON 166.995 71.990 167.020 71.990 167.020 71.980 ;
        RECT 167.020 71.980 186.035 71.990 ;
        POLYGON 167.020 71.980 167.135 71.980 167.135 71.930 ;
        RECT 167.135 71.930 186.035 71.980 ;
        POLYGON 167.135 71.930 167.225 71.930 167.225 71.890 ;
        RECT 167.225 71.890 186.035 71.930 ;
        RECT 119.015 71.865 147.245 71.890 ;
        RECT 48.645 71.820 112.885 71.865 ;
        RECT 16.145 70.440 23.480 71.820 ;
        POLYGON 23.480 71.820 23.730 71.820 23.480 70.440 ;
        POLYGON 48.645 71.820 48.680 71.820 48.680 71.205 ;
        RECT 48.680 71.660 112.885 71.820 ;
        POLYGON 112.885 71.865 112.930 71.865 112.885 71.660 ;
        POLYGON 118.870 71.850 118.870 71.660 118.835 71.660 ;
        RECT 118.870 71.790 147.245 71.865 ;
        POLYGON 147.245 71.890 147.470 71.890 147.245 71.790 ;
        POLYGON 167.225 71.890 167.455 71.890 167.455 71.795 ;
        RECT 167.455 71.795 186.035 71.890 ;
        POLYGON 167.455 71.795 167.465 71.795 167.465 71.790 ;
        RECT 167.465 71.790 186.035 71.795 ;
        RECT 118.870 71.720 147.090 71.790 ;
        POLYGON 147.090 71.790 147.245 71.790 147.090 71.720 ;
        POLYGON 167.465 71.790 167.610 71.790 167.610 71.720 ;
        RECT 167.610 71.720 186.035 71.790 ;
        RECT 118.870 71.675 146.995 71.720 ;
        POLYGON 146.995 71.720 147.090 71.720 146.995 71.675 ;
        POLYGON 167.610 71.720 167.705 71.720 167.705 71.675 ;
        RECT 167.705 71.675 186.035 71.720 ;
        RECT 118.870 71.660 146.765 71.675 ;
        RECT 48.680 71.205 112.260 71.660 ;
        POLYGON 48.680 71.205 48.725 71.205 48.725 70.785 ;
        RECT 48.725 70.785 112.260 71.205 ;
        POLYGON 48.725 70.785 48.760 70.785 48.760 70.445 ;
        RECT 48.760 70.440 112.260 70.785 ;
        RECT 16.145 70.245 22.645 70.440 ;
        POLYGON 14.625 70.245 14.625 65.420 14.030 65.420 ;
        RECT 14.625 65.420 22.645 70.245 ;
        POLYGON 14.030 65.420 14.030 60.390 13.610 60.390 ;
        RECT 14.030 64.415 22.645 65.420 ;
        POLYGON 22.645 70.440 23.480 70.440 22.645 64.415 ;
        POLYGON 48.760 70.440 48.805 70.440 48.805 70.005 ;
        RECT 48.805 70.000 112.260 70.440 ;
        RECT 14.030 60.390 22.335 64.415 ;
        POLYGON 13.610 60.390 13.610 60.000 13.590 60.000 ;
        RECT 13.610 60.000 22.335 60.390 ;
        POLYGON 22.335 64.415 22.645 64.415 22.335 60.000 ;
        RECT 25.000 62.000 45.000 70.000 ;
        POLYGON 48.805 70.000 49.125 70.000 49.125 66.950 ;
        RECT 49.125 68.985 112.260 70.000 ;
        POLYGON 112.260 71.660 112.885 71.660 112.260 68.985 ;
        POLYGON 118.835 71.660 118.835 71.440 118.795 71.440 ;
        RECT 118.835 71.570 146.765 71.660 ;
        POLYGON 146.765 71.675 146.995 71.675 146.765 71.570 ;
        POLYGON 167.705 71.675 167.925 71.675 167.925 71.570 ;
        RECT 167.925 71.570 186.035 71.675 ;
        RECT 118.835 71.440 146.380 71.570 ;
        POLYGON 118.795 71.435 118.795 71.005 118.715 71.005 ;
        RECT 118.795 71.380 146.380 71.440 ;
        POLYGON 146.380 71.570 146.765 71.570 146.380 71.380 ;
        POLYGON 167.925 71.570 167.950 71.570 167.950 71.560 ;
        RECT 167.950 71.560 186.035 71.570 ;
        POLYGON 167.950 71.560 168.255 71.560 168.255 71.420 ;
        RECT 168.255 71.415 186.035 71.560 ;
        POLYGON 168.255 71.415 168.325 71.415 168.325 71.380 ;
        RECT 168.325 71.380 186.035 71.415 ;
        POLYGON 186.035 72.455 187.050 71.380 186.035 71.380 ;
        POLYGON 208.165 72.455 208.165 71.845 207.980 71.845 ;
        RECT 208.165 72.320 229.305 72.460 ;
        POLYGON 229.305 72.475 229.440 72.475 229.305 72.320 ;
        POLYGON 243.970 72.475 243.970 72.410 243.780 72.410 ;
        RECT 243.970 72.410 260.610 72.475 ;
        POLYGON 243.780 72.410 243.780 72.320 243.560 72.320 ;
        RECT 243.780 72.350 260.610 72.410 ;
        POLYGON 260.610 72.475 260.970 72.350 260.610 72.350 ;
        POLYGON 280.935 72.475 281.060 72.475 281.060 72.350 ;
        RECT 281.060 72.350 303.120 72.475 ;
        RECT 243.780 72.320 260.970 72.350 ;
        RECT 208.165 72.205 229.205 72.320 ;
        POLYGON 229.205 72.320 229.305 72.320 229.205 72.205 ;
        POLYGON 243.560 72.320 243.560 72.260 243.410 72.260 ;
        RECT 243.560 72.270 260.970 72.320 ;
        POLYGON 260.970 72.350 261.170 72.270 260.970 72.270 ;
        POLYGON 281.060 72.350 281.140 72.350 281.140 72.270 ;
        RECT 281.140 72.270 303.120 72.350 ;
        RECT 243.560 72.260 261.170 72.270 ;
        POLYGON 243.405 72.260 243.405 72.205 243.270 72.205 ;
        RECT 243.405 72.205 261.170 72.260 ;
        RECT 208.165 72.185 229.190 72.205 ;
        POLYGON 229.190 72.205 229.205 72.205 229.190 72.185 ;
        POLYGON 243.270 72.205 243.270 72.185 243.220 72.185 ;
        RECT 243.270 72.185 261.170 72.205 ;
        RECT 208.165 71.915 228.955 72.185 ;
        POLYGON 228.955 72.185 229.190 72.185 228.955 71.915 ;
        POLYGON 243.220 72.185 243.220 71.980 242.720 71.980 ;
        RECT 243.220 72.125 261.170 72.185 ;
        POLYGON 261.170 72.270 261.535 72.125 261.170 72.125 ;
        POLYGON 281.140 72.270 281.285 72.270 281.285 72.125 ;
        RECT 281.285 72.125 303.120 72.270 ;
        RECT 243.220 72.065 261.535 72.125 ;
        POLYGON 261.535 72.125 261.690 72.065 261.535 72.065 ;
        POLYGON 281.285 72.125 281.345 72.125 281.345 72.065 ;
        RECT 281.345 72.065 303.120 72.125 ;
        RECT 243.220 71.980 261.690 72.065 ;
        POLYGON 242.720 71.980 242.720 71.915 242.575 71.915 ;
        RECT 242.720 71.915 261.690 71.980 ;
        RECT 208.165 71.845 228.705 71.915 ;
        POLYGON 207.980 71.845 207.980 71.565 207.915 71.565 ;
        RECT 207.980 71.620 228.705 71.845 ;
        POLYGON 228.705 71.915 228.955 71.915 228.705 71.620 ;
        POLYGON 242.575 71.915 242.575 71.795 242.310 71.795 ;
        RECT 242.575 71.895 261.690 71.915 ;
        POLYGON 261.690 72.065 262.115 71.895 261.690 71.895 ;
        POLYGON 281.345 72.065 281.405 72.065 281.405 72.005 ;
        RECT 281.405 72.005 303.120 72.065 ;
        POLYGON 281.405 72.005 281.500 72.005 281.500 71.900 ;
        RECT 281.500 71.895 303.120 72.005 ;
        RECT 242.575 71.795 262.115 71.895 ;
        POLYGON 242.310 71.795 242.310 71.620 241.930 71.620 ;
        RECT 242.310 71.620 262.115 71.795 ;
        RECT 207.980 71.565 228.655 71.620 ;
        RECT 207.915 71.560 228.655 71.565 ;
        POLYGON 228.655 71.620 228.705 71.620 228.655 71.560 ;
        POLYGON 241.930 71.620 241.930 71.560 241.800 71.560 ;
        RECT 241.930 71.595 262.115 71.620 ;
        POLYGON 262.115 71.895 262.770 71.595 262.115 71.595 ;
        POLYGON 281.500 71.895 281.775 71.895 281.775 71.595 ;
        RECT 281.775 71.595 303.120 71.895 ;
        RECT 241.930 71.560 262.770 71.595 ;
        POLYGON 262.770 71.595 262.845 71.560 262.770 71.560 ;
        POLYGON 281.775 71.595 281.805 71.595 281.805 71.560 ;
        RECT 281.805 71.560 303.120 71.595 ;
        POLYGON 207.915 71.560 207.915 71.415 207.880 71.415 ;
        RECT 207.915 71.415 228.525 71.560 ;
        RECT 207.880 71.410 228.525 71.415 ;
        POLYGON 228.525 71.560 228.655 71.560 228.525 71.410 ;
        POLYGON 241.800 71.560 241.800 71.545 241.765 71.545 ;
        RECT 241.800 71.545 262.845 71.560 ;
        POLYGON 241.765 71.545 241.765 71.505 241.680 71.505 ;
        RECT 241.765 71.530 262.845 71.545 ;
        POLYGON 262.845 71.560 262.915 71.530 262.845 71.530 ;
        POLYGON 281.805 71.560 281.830 71.560 281.830 71.535 ;
        RECT 281.830 71.530 303.120 71.560 ;
        RECT 241.765 71.505 262.915 71.530 ;
        POLYGON 241.680 71.505 241.680 71.410 241.500 71.410 ;
        RECT 241.680 71.410 262.915 71.505 ;
        RECT 207.880 71.405 228.520 71.410 ;
        POLYGON 228.520 71.410 228.525 71.410 228.520 71.405 ;
        POLYGON 241.500 71.410 241.500 71.405 241.490 71.405 ;
        RECT 241.500 71.405 262.915 71.410 ;
        POLYGON 262.915 71.530 263.185 71.405 262.915 71.405 ;
        POLYGON 281.830 71.530 281.945 71.530 281.945 71.405 ;
        RECT 281.945 71.405 303.120 71.530 ;
        POLYGON 207.880 71.405 207.880 71.380 207.870 71.380 ;
        RECT 207.880 71.380 228.400 71.405 ;
        RECT 118.795 71.225 146.070 71.380 ;
        POLYGON 146.070 71.380 146.380 71.380 146.070 71.225 ;
        POLYGON 168.325 71.380 168.445 71.380 168.445 71.320 ;
        RECT 168.445 71.320 187.050 71.380 ;
        POLYGON 168.445 71.320 168.625 71.320 168.625 71.225 ;
        RECT 168.625 71.230 187.050 71.320 ;
        POLYGON 187.050 71.380 187.180 71.230 187.050 71.230 ;
        POLYGON 207.870 71.370 207.870 71.250 207.840 71.250 ;
        RECT 207.870 71.250 228.400 71.380 ;
        POLYGON 228.400 71.405 228.520 71.405 228.400 71.250 ;
        POLYGON 241.490 71.405 241.490 71.250 241.195 71.250 ;
        RECT 241.490 71.380 263.185 71.405 ;
        POLYGON 263.185 71.405 263.240 71.380 263.185 71.380 ;
        POLYGON 281.945 71.405 281.970 71.405 281.970 71.380 ;
        RECT 281.970 71.380 303.120 71.405 ;
        RECT 241.490 71.250 263.240 71.380 ;
        POLYGON 263.240 71.380 263.490 71.250 263.240 71.250 ;
        POLYGON 281.970 71.380 282.085 71.380 282.085 71.250 ;
        RECT 282.085 71.250 303.120 71.380 ;
        POLYGON 207.840 71.245 207.840 71.230 207.835 71.230 ;
        RECT 207.840 71.230 228.385 71.250 ;
        POLYGON 228.385 71.250 228.400 71.250 228.385 71.230 ;
        POLYGON 241.195 71.250 241.195 71.230 241.155 71.230 ;
        RECT 241.195 71.230 263.490 71.250 ;
        RECT 168.625 71.225 187.180 71.230 ;
        RECT 118.795 71.140 145.910 71.225 ;
        POLYGON 145.910 71.225 146.070 71.225 145.910 71.140 ;
        POLYGON 168.625 71.225 168.790 71.225 168.790 71.140 ;
        RECT 168.790 71.140 187.180 71.225 ;
        RECT 118.795 71.005 145.530 71.140 ;
        POLYGON 118.715 70.995 118.715 70.620 118.645 70.620 ;
        RECT 118.715 70.935 145.530 71.005 ;
        POLYGON 145.530 71.140 145.910 71.140 145.530 70.935 ;
        POLYGON 168.790 71.140 168.840 71.140 168.840 71.115 ;
        RECT 168.840 71.115 187.180 71.140 ;
        POLYGON 168.840 71.115 169.045 71.115 169.045 71.010 ;
        RECT 169.045 71.010 187.180 71.115 ;
        POLYGON 169.045 71.010 169.175 71.010 169.175 70.935 ;
        RECT 169.175 71.000 187.180 71.010 ;
        POLYGON 187.180 71.230 187.385 71.000 187.180 71.000 ;
        POLYGON 207.835 71.220 207.835 71.005 207.785 71.005 ;
        RECT 207.835 71.005 228.210 71.230 ;
        POLYGON 228.210 71.230 228.385 71.230 228.210 71.005 ;
        POLYGON 241.155 71.230 241.155 71.015 240.745 71.015 ;
        RECT 241.155 71.080 263.490 71.230 ;
        POLYGON 263.490 71.250 263.820 71.080 263.490 71.080 ;
        POLYGON 282.085 71.250 282.240 71.250 282.240 71.080 ;
        RECT 282.240 71.080 303.120 71.250 ;
        RECT 241.155 71.015 263.820 71.080 ;
        POLYGON 240.745 71.015 240.745 71.005 240.725 71.005 ;
        RECT 240.745 71.005 263.820 71.015 ;
        POLYGON 263.820 71.080 263.965 71.005 263.820 71.005 ;
        POLYGON 282.240 71.080 282.310 71.080 282.310 71.005 ;
        RECT 282.310 71.005 303.120 71.080 ;
        RECT 169.175 70.935 187.385 71.000 ;
        POLYGON 207.785 71.005 207.785 70.995 207.780 70.995 ;
        RECT 207.785 70.995 227.890 71.005 ;
        RECT 118.715 70.910 145.485 70.935 ;
        POLYGON 145.485 70.935 145.530 70.935 145.485 70.910 ;
        POLYGON 169.175 70.935 169.215 70.935 169.215 70.910 ;
        RECT 169.215 70.910 187.385 70.935 ;
        RECT 118.715 70.860 145.385 70.910 ;
        POLYGON 145.385 70.910 145.485 70.910 145.385 70.860 ;
        POLYGON 169.215 70.910 169.305 70.910 169.305 70.860 ;
        RECT 169.305 70.860 187.385 70.910 ;
        RECT 118.715 70.620 144.850 70.860 ;
        POLYGON 118.645 70.610 118.645 70.415 118.610 70.415 ;
        RECT 118.645 70.545 144.850 70.620 ;
        POLYGON 144.850 70.860 145.385 70.860 144.850 70.545 ;
        POLYGON 169.305 70.860 169.690 70.860 169.690 70.640 ;
        RECT 169.690 70.640 187.385 70.860 ;
        POLYGON 169.690 70.640 169.820 70.640 169.820 70.565 ;
        RECT 169.820 70.565 187.385 70.640 ;
        POLYGON 169.820 70.565 169.850 70.565 169.850 70.545 ;
        RECT 169.850 70.545 187.385 70.565 ;
        RECT 118.645 70.480 144.740 70.545 ;
        POLYGON 144.740 70.545 144.850 70.545 144.740 70.480 ;
        POLYGON 169.850 70.545 169.875 70.545 169.875 70.530 ;
        RECT 169.875 70.530 187.385 70.545 ;
        POLYGON 169.875 70.530 169.955 70.530 169.955 70.480 ;
        RECT 169.955 70.480 187.385 70.530 ;
        RECT 118.645 70.470 144.720 70.480 ;
        POLYGON 144.720 70.480 144.740 70.480 144.720 70.470 ;
        POLYGON 169.955 70.480 169.970 70.480 169.970 70.470 ;
        RECT 169.970 70.470 187.385 70.480 ;
        RECT 118.645 70.450 144.690 70.470 ;
        POLYGON 144.690 70.470 144.720 70.470 144.690 70.450 ;
        POLYGON 169.970 70.470 170.000 70.470 170.000 70.450 ;
        RECT 170.000 70.450 187.385 70.470 ;
        RECT 118.645 70.415 144.065 70.450 ;
        POLYGON 118.610 70.415 118.610 69.805 118.525 69.805 ;
        RECT 118.610 70.060 144.065 70.415 ;
        POLYGON 144.065 70.450 144.690 70.450 144.065 70.060 ;
        POLYGON 170.000 70.450 170.455 70.450 170.455 70.170 ;
        RECT 170.455 70.265 187.385 70.450 ;
        POLYGON 187.385 70.995 188.030 70.265 187.385 70.265 ;
        POLYGON 207.780 70.985 207.780 70.275 207.615 70.275 ;
        RECT 207.780 70.600 227.890 70.995 ;
        POLYGON 227.890 71.005 228.210 71.005 227.890 70.600 ;
        POLYGON 240.725 71.005 240.725 70.975 240.660 70.975 ;
        RECT 240.725 70.975 263.965 71.005 ;
        POLYGON 240.660 70.975 240.660 70.785 240.345 70.785 ;
        RECT 240.660 70.820 263.965 70.975 ;
        POLYGON 263.965 71.005 264.330 70.820 263.965 70.820 ;
        POLYGON 282.310 71.005 282.475 71.005 282.475 70.820 ;
        RECT 282.475 70.820 303.120 71.005 ;
        RECT 240.660 70.805 264.330 70.820 ;
        POLYGON 264.330 70.820 264.355 70.805 264.330 70.805 ;
        POLYGON 282.475 70.820 282.490 70.820 282.490 70.805 ;
        RECT 282.490 70.805 303.120 70.820 ;
        RECT 240.660 70.785 264.355 70.805 ;
        POLYGON 240.345 70.785 240.345 70.600 240.025 70.600 ;
        RECT 240.345 70.600 264.355 70.785 ;
        RECT 207.780 70.515 227.830 70.600 ;
        POLYGON 227.830 70.600 227.890 70.600 227.830 70.515 ;
        POLYGON 240.025 70.600 240.025 70.515 239.880 70.515 ;
        RECT 240.025 70.525 264.355 70.600 ;
        POLYGON 264.355 70.805 264.850 70.525 264.355 70.525 ;
        POLYGON 282.490 70.805 282.550 70.805 282.550 70.740 ;
        RECT 282.550 70.740 303.120 70.805 ;
        POLYGON 282.550 70.740 282.725 70.740 282.725 70.530 ;
        RECT 282.725 70.525 303.120 70.740 ;
        RECT 240.025 70.515 264.850 70.525 ;
        RECT 207.780 70.275 227.650 70.515 ;
        RECT 207.615 70.270 227.650 70.275 ;
        POLYGON 227.650 70.515 227.830 70.515 227.650 70.270 ;
        POLYGON 239.880 70.515 239.880 70.490 239.835 70.490 ;
        RECT 239.880 70.490 264.850 70.515 ;
        POLYGON 239.835 70.490 239.835 70.390 239.670 70.390 ;
        RECT 239.835 70.485 264.850 70.490 ;
        POLYGON 264.850 70.525 264.920 70.485 264.850 70.485 ;
        POLYGON 282.725 70.525 282.760 70.525 282.760 70.485 ;
        RECT 282.760 70.485 303.120 70.525 ;
        RECT 239.835 70.390 264.920 70.485 ;
        POLYGON 239.670 70.390 239.670 70.270 239.485 70.270 ;
        RECT 239.670 70.270 264.920 70.390 ;
        POLYGON 264.920 70.485 265.290 70.270 264.920 70.270 ;
        POLYGON 282.760 70.485 282.940 70.485 282.940 70.270 ;
        RECT 282.940 70.270 303.120 70.485 ;
        RECT 170.455 70.170 188.030 70.265 ;
        POLYGON 207.615 70.270 207.615 70.260 207.610 70.260 ;
        RECT 207.615 70.260 227.520 70.270 ;
        POLYGON 170.455 70.170 170.575 70.170 170.575 70.095 ;
        RECT 170.575 70.095 188.030 70.170 ;
        POLYGON 170.575 70.095 170.625 70.095 170.625 70.060 ;
        RECT 170.625 70.060 188.030 70.095 ;
        RECT 118.610 70.035 144.025 70.060 ;
        POLYGON 144.025 70.060 144.065 70.060 144.025 70.035 ;
        POLYGON 170.625 70.060 170.660 70.060 170.660 70.035 ;
        RECT 170.660 70.035 188.030 70.060 ;
        RECT 118.610 69.945 143.900 70.035 ;
        POLYGON 143.900 70.035 144.025 70.035 143.900 69.945 ;
        POLYGON 170.660 70.035 170.790 70.035 170.790 69.945 ;
        RECT 170.790 69.945 188.030 70.035 ;
        RECT 118.610 69.920 143.885 69.945 ;
        POLYGON 143.885 69.945 143.900 69.945 143.885 69.935 ;
        POLYGON 170.790 69.945 170.805 69.945 170.805 69.935 ;
        RECT 170.805 69.935 188.030 69.945 ;
        POLYGON 170.805 69.935 170.820 69.935 170.820 69.925 ;
        RECT 170.820 69.925 188.030 69.935 ;
        POLYGON 143.885 69.925 143.890 69.920 143.885 69.920 ;
        POLYGON 170.820 69.925 170.830 69.925 170.830 69.920 ;
        RECT 170.830 69.920 188.030 69.925 ;
        RECT 118.610 69.830 143.890 69.920 ;
        POLYGON 170.830 69.920 170.875 69.920 170.875 69.890 ;
        RECT 170.875 69.890 188.030 69.920 ;
        POLYGON 143.890 69.890 143.900 69.830 143.890 69.830 ;
        POLYGON 170.875 69.890 170.960 69.890 170.960 69.830 ;
        RECT 170.960 69.830 188.030 69.890 ;
        RECT 118.610 69.805 143.900 69.830 ;
        POLYGON 118.525 69.795 118.525 69.550 118.490 69.550 ;
        RECT 118.525 69.645 143.900 69.805 ;
        POLYGON 143.900 69.830 143.920 69.645 143.900 69.645 ;
        RECT 118.525 69.600 143.920 69.645 ;
        POLYGON 170.960 69.830 171.260 69.830 171.260 69.630 ;
        RECT 171.260 69.630 188.030 69.830 ;
        POLYGON 171.260 69.630 171.285 69.630 171.285 69.615 ;
        RECT 171.285 69.615 188.030 69.630 ;
        POLYGON 143.920 69.615 143.925 69.600 143.920 69.600 ;
        RECT 118.525 69.550 143.925 69.600 ;
        POLYGON 171.285 69.615 171.345 69.615 171.345 69.570 ;
        RECT 171.345 69.570 188.030 69.615 ;
        POLYGON 118.490 69.540 118.490 69.335 118.460 69.335 ;
        RECT 118.490 69.505 143.925 69.550 ;
        POLYGON 143.925 69.570 143.935 69.505 143.925 69.505 ;
        POLYGON 171.345 69.570 171.435 69.570 171.435 69.505 ;
        RECT 171.435 69.505 188.030 69.570 ;
        RECT 118.490 69.370 143.935 69.505 ;
        POLYGON 143.935 69.505 143.950 69.370 143.935 69.370 ;
        RECT 118.490 69.335 143.950 69.370 ;
        POLYGON 171.435 69.505 171.640 69.505 171.640 69.355 ;
        RECT 171.640 69.355 188.030 69.505 ;
        POLYGON 118.460 69.330 118.460 68.985 118.410 68.985 ;
        RECT 118.460 69.185 143.950 69.335 ;
        POLYGON 143.950 69.355 143.970 69.185 143.950 69.185 ;
        POLYGON 171.640 69.355 171.875 69.355 171.875 69.185 ;
        RECT 171.875 69.335 188.030 69.355 ;
        POLYGON 188.030 70.260 188.785 69.335 188.030 69.335 ;
        POLYGON 207.610 70.255 207.610 69.355 207.400 69.355 ;
        RECT 207.610 70.090 227.520 70.260 ;
        POLYGON 227.520 70.270 227.650 70.270 227.520 70.090 ;
        POLYGON 239.485 70.270 239.485 70.150 239.300 70.150 ;
        RECT 239.485 70.175 265.290 70.270 ;
        POLYGON 265.290 70.270 265.455 70.175 265.290 70.175 ;
        POLYGON 282.940 70.270 283.020 70.270 283.020 70.175 ;
        RECT 283.020 70.175 303.120 70.270 ;
        RECT 239.485 70.150 265.455 70.175 ;
        POLYGON 239.300 70.150 239.300 70.090 239.210 70.090 ;
        RECT 239.300 70.090 265.455 70.150 ;
        RECT 207.610 69.780 227.300 70.090 ;
        POLYGON 227.300 70.090 227.520 70.090 227.300 69.780 ;
        POLYGON 239.210 70.090 239.210 69.925 238.955 69.925 ;
        RECT 239.210 69.945 265.455 70.090 ;
        POLYGON 265.455 70.175 265.810 69.945 265.455 69.945 ;
        POLYGON 283.020 70.175 283.210 70.175 283.210 69.950 ;
        RECT 283.210 69.945 303.120 70.175 ;
        RECT 239.210 69.925 265.810 69.945 ;
        POLYGON 238.955 69.925 238.955 69.780 238.740 69.780 ;
        RECT 238.955 69.920 265.810 69.925 ;
        POLYGON 265.810 69.945 265.850 69.920 265.810 69.920 ;
        POLYGON 283.210 69.945 283.235 69.945 283.235 69.920 ;
        RECT 283.235 69.920 303.120 69.945 ;
        RECT 238.955 69.855 265.850 69.920 ;
        POLYGON 265.850 69.920 265.950 69.855 265.850 69.855 ;
        POLYGON 283.235 69.920 283.285 69.920 283.285 69.860 ;
        RECT 283.285 69.855 303.120 69.920 ;
        RECT 238.955 69.780 265.950 69.855 ;
        RECT 207.610 69.775 227.295 69.780 ;
        POLYGON 227.295 69.780 227.300 69.780 227.295 69.775 ;
        POLYGON 238.740 69.780 238.740 69.775 238.730 69.775 ;
        RECT 238.740 69.775 265.950 69.780 ;
        RECT 207.610 69.450 227.075 69.775 ;
        POLYGON 227.075 69.775 227.295 69.775 227.075 69.450 ;
        POLYGON 238.730 69.775 238.730 69.760 238.710 69.760 ;
        RECT 238.730 69.760 265.950 69.775 ;
        POLYGON 238.710 69.760 238.710 69.450 238.285 69.450 ;
        RECT 238.710 69.490 265.950 69.760 ;
        POLYGON 265.950 69.855 266.470 69.490 265.950 69.490 ;
        POLYGON 283.285 69.855 283.590 69.855 283.590 69.495 ;
        RECT 283.590 69.490 303.120 69.855 ;
        RECT 238.710 69.450 266.470 69.490 ;
        RECT 207.610 69.355 227.010 69.450 ;
        POLYGON 227.010 69.450 227.075 69.450 227.010 69.355 ;
        POLYGON 238.285 69.450 238.285 69.355 238.155 69.355 ;
        RECT 238.285 69.355 266.470 69.450 ;
        RECT 171.875 69.185 188.785 69.335 ;
        POLYGON 207.400 69.350 207.400 69.330 207.395 69.330 ;
        RECT 207.400 69.330 226.845 69.355 ;
        RECT 118.460 69.140 143.970 69.185 ;
        POLYGON 171.875 69.185 171.885 69.185 171.885 69.175 ;
        RECT 171.885 69.175 188.785 69.185 ;
        POLYGON 143.970 69.175 143.975 69.140 143.970 69.140 ;
        RECT 118.460 69.050 143.975 69.140 ;
        POLYGON 171.885 69.175 171.980 69.175 171.980 69.105 ;
        RECT 171.980 69.105 188.785 69.175 ;
        POLYGON 188.785 69.330 188.970 69.105 188.785 69.105 ;
        POLYGON 207.395 69.330 207.395 69.115 207.345 69.115 ;
        RECT 207.395 69.115 226.845 69.330 ;
        RECT 207.345 69.110 226.845 69.115 ;
        POLYGON 226.845 69.355 227.010 69.355 226.845 69.110 ;
        POLYGON 238.155 69.355 238.155 69.200 237.940 69.200 ;
        RECT 238.155 69.220 266.470 69.355 ;
        POLYGON 266.470 69.490 266.830 69.220 266.470 69.220 ;
        POLYGON 283.590 69.490 283.645 69.490 283.645 69.430 ;
        RECT 283.645 69.430 303.120 69.490 ;
        POLYGON 283.645 69.430 283.700 69.430 283.700 69.355 ;
        RECT 283.700 69.355 303.120 69.430 ;
        POLYGON 283.700 69.355 283.805 69.355 283.805 69.220 ;
        RECT 283.805 69.220 303.120 69.355 ;
        RECT 238.155 69.200 266.830 69.220 ;
        POLYGON 237.940 69.200 237.940 69.110 237.815 69.110 ;
        RECT 237.940 69.110 266.830 69.200 ;
        POLYGON 266.830 69.220 266.970 69.110 266.830 69.110 ;
        POLYGON 283.805 69.220 283.885 69.220 283.885 69.115 ;
        RECT 283.885 69.110 303.120 69.220 ;
        POLYGON 171.980 69.105 171.985 69.105 171.985 69.100 ;
        RECT 171.985 69.100 188.970 69.105 ;
        POLYGON 188.970 69.105 188.975 69.100 188.970 69.100 ;
        POLYGON 207.345 69.105 207.345 69.100 207.340 69.100 ;
        RECT 207.345 69.100 226.785 69.110 ;
        POLYGON 143.975 69.100 143.985 69.050 143.975 69.050 ;
        RECT 118.460 68.985 143.985 69.050 ;
        POLYGON 171.985 69.100 172.060 69.100 172.060 69.045 ;
        RECT 172.060 69.045 188.975 69.100 ;
        RECT 49.125 68.520 112.180 68.985 ;
        POLYGON 112.180 68.985 112.260 68.985 112.180 68.520 ;
        POLYGON 118.410 68.960 118.410 68.520 118.345 68.520 ;
        RECT 118.410 68.910 143.985 68.985 ;
        POLYGON 143.985 69.045 144.000 68.910 143.985 68.910 ;
        RECT 118.410 68.775 144.000 68.910 ;
        POLYGON 172.060 69.045 172.270 69.045 172.270 68.880 ;
        RECT 172.270 68.880 188.975 69.045 ;
        POLYGON 144.000 68.880 144.015 68.775 144.000 68.775 ;
        RECT 118.410 68.730 144.015 68.775 ;
        POLYGON 172.270 68.880 172.445 68.880 172.445 68.740 ;
        RECT 172.445 68.740 188.975 68.880 ;
        POLYGON 144.015 68.740 144.020 68.730 144.015 68.730 ;
        RECT 118.410 68.680 144.020 68.730 ;
        POLYGON 172.445 68.740 172.480 68.740 172.480 68.710 ;
        RECT 172.480 68.710 188.975 68.740 ;
        POLYGON 144.020 68.710 144.025 68.680 144.020 68.680 ;
        RECT 118.410 68.635 144.025 68.680 ;
        POLYGON 172.480 68.710 172.545 68.710 172.545 68.660 ;
        RECT 172.545 68.670 188.975 68.710 ;
        POLYGON 188.975 69.100 189.300 68.670 188.975 68.670 ;
        POLYGON 207.340 69.095 207.340 68.965 207.310 68.965 ;
        RECT 207.340 69.020 226.785 69.100 ;
        POLYGON 226.785 69.110 226.845 69.110 226.785 69.020 ;
        POLYGON 237.815 69.110 237.815 69.080 237.775 69.080 ;
        RECT 237.815 69.080 266.970 69.110 ;
        POLYGON 237.775 69.080 237.775 69.020 237.700 69.020 ;
        RECT 237.775 69.075 266.970 69.080 ;
        POLYGON 266.970 69.110 267.015 69.075 266.970 69.075 ;
        POLYGON 283.885 69.110 283.915 69.110 283.915 69.075 ;
        RECT 283.915 69.075 303.120 69.110 ;
        RECT 237.775 69.020 267.015 69.075 ;
        RECT 207.340 68.965 226.730 69.020 ;
        POLYGON 207.310 68.965 207.310 68.680 207.260 68.680 ;
        RECT 207.310 68.940 226.730 68.965 ;
        POLYGON 226.730 69.020 226.785 69.020 226.730 68.940 ;
        POLYGON 237.700 69.020 237.700 68.940 237.605 68.940 ;
        RECT 237.700 68.940 267.015 69.020 ;
        RECT 207.310 68.680 226.570 68.940 ;
        POLYGON 226.570 68.940 226.730 68.940 226.570 68.685 ;
        POLYGON 237.605 68.940 237.605 68.685 237.290 68.685 ;
        RECT 237.605 68.745 267.015 68.940 ;
        POLYGON 267.015 69.075 267.430 68.745 267.015 68.745 ;
        POLYGON 283.915 69.075 284.165 69.075 284.165 68.750 ;
        RECT 284.165 68.745 303.120 69.075 ;
        RECT 237.605 68.685 267.430 68.745 ;
        POLYGON 237.290 68.685 237.290 68.680 237.285 68.680 ;
        RECT 237.290 68.680 267.430 68.685 ;
        POLYGON 267.430 68.745 267.505 68.680 267.430 68.680 ;
        POLYGON 284.165 68.745 284.215 68.745 284.215 68.680 ;
        RECT 284.215 68.680 303.120 68.745 ;
        RECT 172.545 68.660 189.300 68.670 ;
        POLYGON 156.240 68.660 156.240 68.650 155.855 68.650 ;
        POLYGON 156.240 68.660 156.400 68.655 156.240 68.655 ;
        POLYGON 172.545 68.660 172.550 68.660 172.550 68.655 ;
        RECT 172.550 68.655 189.300 68.660 ;
        RECT 156.240 68.650 156.650 68.655 ;
        POLYGON 156.650 68.655 156.900 68.650 156.650 68.650 ;
        POLYGON 172.550 68.655 172.555 68.655 172.555 68.650 ;
        RECT 172.555 68.650 189.300 68.655 ;
        POLYGON 155.835 68.650 155.835 68.645 155.615 68.645 ;
        RECT 155.835 68.645 156.975 68.650 ;
        POLYGON 155.595 68.645 155.595 68.640 155.500 68.640 ;
        RECT 155.595 68.640 156.975 68.645 ;
        POLYGON 144.025 68.640 144.030 68.635 144.025 68.635 ;
        RECT 118.410 68.590 144.030 68.635 ;
        POLYGON 155.500 68.640 155.500 68.630 155.285 68.630 ;
        RECT 155.500 68.635 156.975 68.640 ;
        POLYGON 156.975 68.650 157.285 68.635 156.975 68.635 ;
        POLYGON 172.555 68.650 172.575 68.650 172.575 68.635 ;
        RECT 172.575 68.635 189.300 68.650 ;
        RECT 155.500 68.630 157.305 68.635 ;
        POLYGON 155.285 68.630 155.285 68.620 155.065 68.620 ;
        RECT 155.285 68.620 157.305 68.630 ;
        POLYGON 157.305 68.635 157.595 68.620 157.305 68.620 ;
        POLYGON 172.575 68.635 172.595 68.635 172.595 68.620 ;
        RECT 172.595 68.620 189.300 68.635 ;
        POLYGON 155.065 68.620 155.065 68.600 154.770 68.600 ;
        RECT 155.065 68.615 157.600 68.620 ;
        POLYGON 157.600 68.620 157.710 68.615 157.600 68.615 ;
        POLYGON 172.595 68.620 172.600 68.620 172.600 68.615 ;
        RECT 172.600 68.615 189.300 68.620 ;
        RECT 155.065 68.600 157.710 68.615 ;
        POLYGON 144.030 68.600 144.035 68.590 144.030 68.590 ;
        RECT 118.410 68.545 144.035 68.590 ;
        POLYGON 154.770 68.600 154.770 68.555 154.275 68.555 ;
        RECT 154.770 68.575 157.710 68.600 ;
        POLYGON 157.710 68.615 158.245 68.575 157.710 68.575 ;
        POLYGON 172.600 68.615 172.615 68.615 172.615 68.605 ;
        RECT 172.615 68.605 189.300 68.615 ;
        POLYGON 172.615 68.605 172.650 68.605 172.650 68.580 ;
        RECT 172.650 68.580 189.300 68.605 ;
        POLYGON 172.650 68.580 172.655 68.580 172.655 68.575 ;
        RECT 172.655 68.575 189.300 68.580 ;
        RECT 154.770 68.560 158.245 68.575 ;
        POLYGON 158.245 68.575 158.435 68.560 158.245 68.560 ;
        POLYGON 172.655 68.575 172.670 68.575 172.670 68.560 ;
        RECT 172.670 68.560 189.300 68.575 ;
        RECT 154.770 68.555 158.435 68.560 ;
        POLYGON 144.035 68.555 144.040 68.545 144.035 68.545 ;
        POLYGON 154.275 68.555 154.275 68.545 154.120 68.545 ;
        RECT 154.275 68.545 158.435 68.555 ;
        RECT 118.410 68.520 144.040 68.545 ;
        POLYGON 154.115 68.545 154.115 68.540 154.070 68.540 ;
        RECT 154.115 68.540 158.435 68.545 ;
        POLYGON 154.070 68.540 154.070 68.535 154.045 68.535 ;
        RECT 154.070 68.535 158.435 68.540 ;
        RECT 49.125 67.565 112.015 68.520 ;
        POLYGON 112.015 68.520 112.180 68.520 112.015 67.565 ;
        POLYGON 118.345 68.505 118.345 68.110 118.290 68.110 ;
        RECT 118.345 68.500 144.040 68.520 ;
        POLYGON 144.040 68.535 144.045 68.500 144.040 68.500 ;
        RECT 118.345 68.455 144.045 68.500 ;
        POLYGON 154.045 68.535 154.045 68.465 153.490 68.465 ;
        RECT 154.045 68.490 158.435 68.535 ;
        POLYGON 158.435 68.560 159.045 68.490 158.435 68.490 ;
        POLYGON 172.670 68.560 172.760 68.560 172.760 68.490 ;
        RECT 172.760 68.490 189.300 68.560 ;
        RECT 154.045 68.485 159.045 68.490 ;
        POLYGON 159.045 68.490 159.070 68.485 159.045 68.485 ;
        POLYGON 172.760 68.490 172.770 68.490 172.770 68.485 ;
        RECT 172.770 68.485 189.300 68.490 ;
        RECT 154.045 68.475 159.075 68.485 ;
        POLYGON 159.075 68.485 159.145 68.475 159.075 68.475 ;
        POLYGON 172.770 68.485 172.780 68.485 172.780 68.475 ;
        RECT 172.780 68.475 189.300 68.485 ;
        RECT 154.045 68.465 159.145 68.475 ;
        POLYGON 144.045 68.465 144.050 68.455 144.045 68.455 ;
        RECT 118.345 68.405 144.050 68.455 ;
        POLYGON 153.490 68.465 153.490 68.450 153.335 68.450 ;
        RECT 153.490 68.450 159.145 68.465 ;
        POLYGON 144.050 68.450 144.055 68.405 144.050 68.405 ;
        RECT 118.345 68.360 144.055 68.405 ;
        POLYGON 153.335 68.450 153.335 68.385 152.950 68.385 ;
        RECT 153.335 68.385 159.145 68.450 ;
        POLYGON 152.950 68.385 152.950 68.375 152.890 68.375 ;
        RECT 152.950 68.375 159.145 68.385 ;
        POLYGON 144.055 68.375 144.060 68.360 144.055 68.360 ;
        RECT 118.345 68.225 144.060 68.360 ;
        POLYGON 152.890 68.375 152.890 68.350 152.745 68.350 ;
        RECT 152.890 68.370 159.145 68.375 ;
        POLYGON 159.145 68.475 159.845 68.370 159.145 68.370 ;
        POLYGON 172.780 68.475 172.790 68.475 172.790 68.470 ;
        RECT 172.790 68.470 189.300 68.475 ;
        POLYGON 172.790 68.470 172.905 68.470 172.905 68.370 ;
        RECT 172.905 68.370 189.300 68.470 ;
        RECT 152.890 68.365 159.845 68.370 ;
        POLYGON 159.845 68.370 159.865 68.365 159.845 68.365 ;
        POLYGON 172.905 68.370 172.910 68.370 172.910 68.365 ;
        RECT 172.910 68.365 189.300 68.370 ;
        RECT 152.890 68.350 159.865 68.365 ;
        POLYGON 152.745 68.350 152.745 68.345 152.715 68.345 ;
        RECT 152.745 68.345 159.865 68.350 ;
        POLYGON 152.710 68.345 152.710 68.335 152.640 68.335 ;
        RECT 152.710 68.335 159.865 68.345 ;
        POLYGON 144.060 68.335 144.075 68.225 144.060 68.225 ;
        RECT 118.345 68.180 144.075 68.225 ;
        POLYGON 152.640 68.335 152.640 68.220 152.090 68.220 ;
        RECT 152.640 68.240 159.865 68.335 ;
        POLYGON 159.865 68.365 160.520 68.240 159.865 68.240 ;
        POLYGON 172.910 68.365 173.060 68.365 173.060 68.240 ;
        RECT 173.060 68.240 189.300 68.365 ;
        RECT 152.640 68.220 160.520 68.240 ;
        POLYGON 152.090 68.220 152.090 68.195 151.970 68.195 ;
        RECT 152.090 68.210 160.520 68.220 ;
        POLYGON 160.520 68.240 160.635 68.210 160.520 68.210 ;
        POLYGON 173.060 68.240 173.095 68.240 173.095 68.210 ;
        RECT 173.095 68.210 189.300 68.240 ;
        RECT 152.090 68.195 160.635 68.210 ;
        POLYGON 151.965 68.195 151.965 68.190 151.940 68.190 ;
        RECT 151.965 68.190 160.635 68.195 ;
        POLYGON 144.075 68.190 144.080 68.180 144.075 68.180 ;
        RECT 118.345 68.130 144.080 68.180 ;
        POLYGON 151.935 68.190 151.935 68.150 151.790 68.150 ;
        RECT 151.935 68.160 160.635 68.190 ;
        POLYGON 160.635 68.210 160.850 68.160 160.635 68.160 ;
        POLYGON 173.095 68.210 173.155 68.210 173.155 68.160 ;
        RECT 173.155 68.160 189.300 68.210 ;
        RECT 151.935 68.150 160.850 68.160 ;
        POLYGON 144.080 68.150 144.085 68.130 144.080 68.130 ;
        RECT 118.345 68.110 144.085 68.130 ;
        POLYGON 118.290 68.105 118.290 67.570 118.215 67.570 ;
        RECT 118.290 68.085 144.085 68.110 ;
        POLYGON 151.790 68.150 151.790 68.095 151.550 68.095 ;
        RECT 151.790 68.130 160.850 68.150 ;
        POLYGON 160.850 68.160 160.970 68.130 160.850 68.130 ;
        POLYGON 173.155 68.160 173.190 68.160 173.190 68.130 ;
        RECT 173.190 68.130 189.300 68.160 ;
        RECT 151.790 68.095 160.970 68.130 ;
        POLYGON 144.085 68.095 144.090 68.085 144.085 68.085 ;
        RECT 118.290 68.040 144.090 68.085 ;
        POLYGON 151.550 68.095 151.550 68.070 151.455 68.070 ;
        RECT 151.550 68.085 160.970 68.095 ;
        POLYGON 160.970 68.130 161.175 68.085 160.970 68.085 ;
        POLYGON 173.190 68.130 173.245 68.130 173.245 68.085 ;
        RECT 173.245 68.085 189.300 68.130 ;
        RECT 151.550 68.070 161.175 68.085 ;
        POLYGON 144.090 68.070 144.095 68.040 144.090 68.040 ;
        RECT 118.290 67.995 144.095 68.040 ;
        POLYGON 151.455 68.070 151.455 68.035 151.320 68.035 ;
        RECT 151.455 68.035 161.175 68.070 ;
        POLYGON 144.095 68.035 144.100 67.995 144.095 67.995 ;
        RECT 118.290 67.860 144.100 67.995 ;
        POLYGON 151.320 68.035 151.320 67.990 151.175 67.990 ;
        RECT 151.320 68.010 161.175 68.035 ;
        POLYGON 161.175 68.085 161.430 68.010 161.175 68.010 ;
        POLYGON 173.245 68.085 173.275 68.085 173.275 68.060 ;
        RECT 173.275 68.060 189.300 68.085 ;
        POLYGON 173.275 68.060 173.330 68.060 173.330 68.010 ;
        RECT 173.330 68.010 189.300 68.060 ;
        RECT 151.320 67.990 161.430 68.010 ;
        POLYGON 144.100 67.990 144.115 67.860 144.100 67.860 ;
        RECT 118.290 67.765 144.115 67.860 ;
        POLYGON 151.170 67.990 151.170 67.850 150.695 67.850 ;
        RECT 151.170 67.900 161.430 67.990 ;
        POLYGON 161.430 68.010 161.805 67.900 161.430 67.900 ;
        POLYGON 173.330 68.010 173.390 68.010 173.390 67.960 ;
        RECT 173.390 67.960 189.300 68.010 ;
        POLYGON 173.390 67.960 173.455 67.960 173.455 67.900 ;
        RECT 173.455 67.905 189.300 67.960 ;
        POLYGON 189.300 68.670 189.875 67.905 189.300 67.905 ;
        POLYGON 207.260 68.670 207.260 67.925 207.130 67.925 ;
        RECT 207.260 68.345 226.360 68.680 ;
        POLYGON 226.360 68.680 226.570 68.680 226.360 68.345 ;
        POLYGON 237.285 68.680 237.285 68.350 236.875 68.350 ;
        RECT 237.285 68.640 267.505 68.680 ;
        RECT 237.285 68.630 250.930 68.640 ;
        POLYGON 250.930 68.640 251.245 68.640 250.930 68.630 ;
        POLYGON 251.245 68.640 251.410 68.640 251.410 68.635 ;
        RECT 251.410 68.635 267.505 68.640 ;
        POLYGON 251.655 68.635 251.985 68.635 251.985 68.630 ;
        RECT 251.985 68.630 267.505 68.635 ;
        RECT 237.285 68.625 250.510 68.630 ;
        POLYGON 250.510 68.630 250.925 68.630 250.510 68.625 ;
        POLYGON 251.985 68.630 252.070 68.630 252.070 68.625 ;
        RECT 252.070 68.625 267.505 68.630 ;
        POLYGON 267.505 68.680 267.575 68.625 267.505 68.625 ;
        POLYGON 284.215 68.680 284.260 68.680 284.260 68.625 ;
        RECT 284.260 68.625 303.120 68.680 ;
        RECT 237.285 68.620 250.500 68.625 ;
        POLYGON 250.500 68.625 250.510 68.625 250.500 68.620 ;
        POLYGON 252.075 68.625 252.205 68.625 252.205 68.620 ;
        RECT 252.205 68.620 267.575 68.625 ;
        RECT 237.285 68.590 249.925 68.620 ;
        POLYGON 249.925 68.620 250.495 68.620 249.925 68.590 ;
        POLYGON 252.205 68.620 252.340 68.620 252.340 68.615 ;
        RECT 252.340 68.615 267.575 68.620 ;
        POLYGON 252.340 68.615 252.715 68.615 252.715 68.595 ;
        RECT 252.715 68.595 267.575 68.615 ;
        POLYGON 252.715 68.595 252.805 68.595 252.805 68.590 ;
        RECT 252.805 68.590 267.575 68.595 ;
        RECT 237.285 68.585 249.780 68.590 ;
        POLYGON 249.780 68.590 249.925 68.590 249.780 68.585 ;
        POLYGON 252.820 68.590 252.875 68.590 252.875 68.585 ;
        RECT 252.875 68.585 267.575 68.590 ;
        RECT 237.285 68.580 249.760 68.585 ;
        POLYGON 249.760 68.585 249.780 68.585 249.760 68.580 ;
        POLYGON 252.875 68.585 252.930 68.585 252.930 68.580 ;
        RECT 252.930 68.580 267.575 68.585 ;
        RECT 237.285 68.545 249.345 68.580 ;
        POLYGON 249.345 68.580 249.760 68.580 249.345 68.545 ;
        POLYGON 252.930 68.580 253.155 68.580 253.155 68.560 ;
        RECT 253.155 68.560 267.575 68.580 ;
        POLYGON 253.195 68.560 253.375 68.560 253.375 68.545 ;
        RECT 253.375 68.545 267.575 68.560 ;
        RECT 237.285 68.520 249.060 68.545 ;
        POLYGON 249.060 68.545 249.345 68.545 249.060 68.520 ;
        POLYGON 253.375 68.545 253.440 68.545 253.440 68.540 ;
        RECT 253.440 68.540 267.575 68.545 ;
        POLYGON 253.440 68.540 253.605 68.540 253.605 68.520 ;
        RECT 253.605 68.520 267.575 68.540 ;
        RECT 237.285 68.500 248.905 68.520 ;
        POLYGON 248.905 68.520 249.060 68.520 248.905 68.500 ;
        POLYGON 253.605 68.520 253.770 68.520 253.770 68.500 ;
        RECT 253.770 68.500 267.575 68.520 ;
        RECT 237.285 68.490 248.845 68.500 ;
        POLYGON 248.845 68.500 248.905 68.500 248.845 68.490 ;
        POLYGON 253.770 68.500 253.855 68.500 253.855 68.490 ;
        RECT 253.855 68.490 267.575 68.500 ;
        RECT 237.285 68.430 248.350 68.490 ;
        POLYGON 248.350 68.490 248.840 68.490 248.350 68.430 ;
        POLYGON 253.855 68.490 253.980 68.490 253.980 68.475 ;
        RECT 253.980 68.475 267.575 68.490 ;
        POLYGON 253.990 68.475 254.040 68.475 254.040 68.470 ;
        RECT 254.040 68.470 267.575 68.475 ;
        POLYGON 254.045 68.470 254.220 68.470 254.220 68.445 ;
        RECT 254.220 68.445 267.575 68.470 ;
        POLYGON 267.575 68.625 267.780 68.445 267.575 68.445 ;
        POLYGON 284.260 68.625 284.280 68.625 284.280 68.600 ;
        RECT 284.280 68.600 303.120 68.625 ;
        POLYGON 284.280 68.600 284.395 68.600 284.395 68.450 ;
        RECT 284.395 68.445 303.120 68.600 ;
        POLYGON 254.220 68.445 254.315 68.445 254.315 68.430 ;
        RECT 254.315 68.430 267.780 68.445 ;
        RECT 237.285 68.405 248.205 68.430 ;
        POLYGON 248.205 68.430 248.350 68.430 248.205 68.405 ;
        POLYGON 254.315 68.430 254.485 68.430 254.485 68.405 ;
        RECT 254.485 68.405 267.780 68.430 ;
        RECT 237.285 68.380 248.055 68.405 ;
        POLYGON 248.055 68.405 248.205 68.405 248.055 68.380 ;
        POLYGON 254.485 68.405 254.650 68.405 254.650 68.380 ;
        RECT 254.650 68.380 267.780 68.405 ;
        RECT 237.285 68.350 247.765 68.380 ;
        POLYGON 236.870 68.350 236.870 68.345 236.865 68.345 ;
        RECT 236.870 68.345 247.765 68.350 ;
        RECT 207.260 68.245 226.300 68.345 ;
        POLYGON 226.300 68.345 226.360 68.345 226.300 68.245 ;
        POLYGON 236.865 68.345 236.865 68.245 236.755 68.245 ;
        RECT 236.865 68.335 247.765 68.345 ;
        POLYGON 247.765 68.380 248.055 68.380 247.765 68.335 ;
        POLYGON 254.650 68.380 254.850 68.380 254.850 68.350 ;
        RECT 254.850 68.350 267.780 68.380 ;
        POLYGON 254.850 68.350 254.880 68.350 254.880 68.345 ;
        RECT 254.880 68.345 267.780 68.350 ;
        POLYGON 254.885 68.345 254.930 68.345 254.930 68.335 ;
        RECT 254.930 68.335 267.780 68.345 ;
        RECT 236.865 68.315 247.655 68.335 ;
        POLYGON 247.655 68.335 247.760 68.335 247.655 68.315 ;
        POLYGON 254.930 68.335 255.030 68.335 255.030 68.315 ;
        RECT 255.030 68.315 267.780 68.335 ;
        RECT 236.865 68.245 247.210 68.315 ;
        RECT 207.260 68.085 226.200 68.245 ;
        POLYGON 226.200 68.245 226.300 68.245 226.200 68.085 ;
        POLYGON 236.755 68.245 236.755 68.115 236.610 68.115 ;
        RECT 236.755 68.225 247.210 68.245 ;
        POLYGON 247.210 68.315 247.655 68.315 247.210 68.225 ;
        POLYGON 255.030 68.315 255.155 68.315 255.155 68.290 ;
        RECT 255.155 68.290 267.780 68.315 ;
        POLYGON 255.160 68.290 255.290 68.290 255.290 68.265 ;
        RECT 255.290 68.265 267.780 68.290 ;
        POLYGON 255.295 68.265 255.495 68.265 255.495 68.225 ;
        RECT 255.495 68.225 267.780 68.265 ;
        RECT 236.755 68.200 247.080 68.225 ;
        POLYGON 247.080 68.225 247.210 68.225 247.080 68.200 ;
        POLYGON 255.495 68.225 255.525 68.225 255.525 68.220 ;
        RECT 255.525 68.220 267.780 68.225 ;
        POLYGON 255.525 68.220 255.605 68.220 255.605 68.200 ;
        RECT 255.605 68.200 267.780 68.220 ;
        RECT 236.755 68.195 247.075 68.200 ;
        RECT 236.755 68.180 246.980 68.195 ;
        POLYGON 246.980 68.195 247.075 68.195 246.980 68.180 ;
        POLYGON 255.605 68.200 255.690 68.200 255.690 68.180 ;
        RECT 255.690 68.180 267.780 68.200 ;
        RECT 236.755 68.115 246.685 68.180 ;
        POLYGON 236.610 68.115 236.610 68.085 236.575 68.085 ;
        RECT 236.610 68.105 246.685 68.115 ;
        POLYGON 246.685 68.180 246.980 68.180 246.685 68.105 ;
        POLYGON 255.690 68.180 255.715 68.180 255.715 68.175 ;
        RECT 255.715 68.175 267.780 68.180 ;
        POLYGON 255.720 68.175 256.010 68.175 256.010 68.105 ;
        RECT 256.010 68.105 267.780 68.175 ;
        RECT 236.610 68.085 246.380 68.105 ;
        RECT 207.260 67.925 226.100 68.085 ;
        POLYGON 207.130 67.915 207.130 67.905 207.125 67.905 ;
        RECT 207.130 67.910 226.100 67.925 ;
        POLYGON 226.100 68.085 226.200 68.085 226.100 67.915 ;
        POLYGON 236.575 68.085 236.575 67.935 236.410 67.935 ;
        RECT 236.575 68.025 246.380 68.085 ;
        POLYGON 246.380 68.105 246.685 68.105 246.380 68.025 ;
        POLYGON 256.010 68.105 256.180 68.105 256.180 68.065 ;
        RECT 256.180 68.065 267.780 68.105 ;
        POLYGON 256.180 68.065 256.325 68.065 256.325 68.025 ;
        RECT 256.325 68.025 267.780 68.065 ;
        RECT 236.575 68.015 246.330 68.025 ;
        POLYGON 246.330 68.025 246.375 68.025 246.330 68.015 ;
        POLYGON 256.325 68.025 256.330 68.025 256.330 68.020 ;
        RECT 256.330 68.020 267.780 68.025 ;
        POLYGON 256.330 68.020 256.355 68.020 256.355 68.015 ;
        RECT 256.355 68.015 267.780 68.020 ;
        RECT 236.575 67.935 245.995 68.015 ;
        POLYGON 236.410 67.935 236.410 67.915 236.390 67.915 ;
        RECT 236.410 67.915 245.995 67.935 ;
        POLYGON 245.995 68.015 246.330 68.015 245.995 67.915 ;
        POLYGON 256.360 68.015 256.535 68.015 256.535 67.960 ;
        RECT 256.535 67.960 267.780 68.015 ;
        POLYGON 256.540 67.960 256.695 67.960 256.695 67.915 ;
        RECT 256.695 67.915 267.780 67.960 ;
        POLYGON 267.780 68.445 268.385 67.915 267.780 67.915 ;
        POLYGON 284.395 68.445 284.690 68.445 284.690 68.070 ;
        RECT 284.690 68.070 303.120 68.445 ;
        POLYGON 284.690 68.070 284.795 68.070 284.795 67.920 ;
        RECT 284.795 67.915 303.120 68.070 ;
        RECT 207.130 67.905 226.070 67.910 ;
        RECT 173.455 67.900 189.875 67.905 ;
        RECT 151.170 67.850 161.805 67.900 ;
        POLYGON 150.695 67.850 150.695 67.825 150.635 67.825 ;
        RECT 150.695 67.825 161.805 67.850 ;
        POLYGON 144.115 67.825 144.125 67.765 144.115 67.765 ;
        RECT 118.290 67.720 144.125 67.765 ;
        POLYGON 150.630 67.825 150.630 67.745 150.415 67.745 ;
        RECT 150.630 67.815 161.805 67.825 ;
        POLYGON 161.805 67.900 162.050 67.815 161.805 67.815 ;
        POLYGON 173.455 67.900 173.505 67.900 173.505 67.860 ;
        RECT 173.505 67.860 189.875 67.900 ;
        POLYGON 173.505 67.860 173.555 67.860 173.555 67.815 ;
        RECT 173.555 67.830 189.875 67.860 ;
        POLYGON 189.875 67.905 189.930 67.830 189.875 67.830 ;
        POLYGON 207.125 67.895 207.125 67.870 207.120 67.870 ;
        RECT 207.125 67.870 226.070 67.905 ;
        RECT 207.120 67.855 226.070 67.870 ;
        POLYGON 226.070 67.910 226.100 67.910 226.070 67.860 ;
        POLYGON 236.390 67.915 236.390 67.860 236.330 67.860 ;
        RECT 236.390 67.905 245.960 67.915 ;
        POLYGON 245.960 67.915 245.995 67.915 245.960 67.905 ;
        POLYGON 256.695 67.915 256.730 67.915 256.730 67.905 ;
        RECT 256.730 67.905 268.385 67.915 ;
        RECT 236.390 67.860 245.795 67.905 ;
        POLYGON 236.330 67.860 236.330 67.855 236.325 67.855 ;
        RECT 236.330 67.855 245.795 67.860 ;
        POLYGON 245.795 67.905 245.960 67.905 245.795 67.855 ;
        POLYGON 256.730 67.905 256.805 67.905 256.805 67.885 ;
        RECT 256.805 67.885 268.385 67.905 ;
        POLYGON 256.805 67.885 256.890 67.885 256.890 67.855 ;
        RECT 256.890 67.855 268.385 67.885 ;
        POLYGON 268.385 67.915 268.450 67.855 268.385 67.855 ;
        POLYGON 284.795 67.915 284.840 67.915 284.840 67.855 ;
        RECT 284.840 67.855 303.120 67.915 ;
        POLYGON 207.120 67.855 207.120 67.840 207.115 67.840 ;
        RECT 207.120 67.840 226.000 67.855 ;
        RECT 173.555 67.815 189.930 67.830 ;
        RECT 150.630 67.760 162.055 67.815 ;
        POLYGON 162.055 67.815 162.220 67.760 162.055 67.760 ;
        POLYGON 173.555 67.815 173.615 67.815 173.615 67.760 ;
        RECT 173.615 67.760 189.930 67.815 ;
        RECT 150.630 67.745 162.220 67.760 ;
        POLYGON 150.410 67.745 150.410 67.735 150.380 67.735 ;
        RECT 150.410 67.735 162.220 67.745 ;
        POLYGON 144.125 67.735 144.130 67.720 144.125 67.720 ;
        RECT 118.290 67.570 144.130 67.720 ;
        POLYGON 150.380 67.735 150.380 67.675 150.210 67.675 ;
        RECT 150.380 67.675 162.220 67.735 ;
        RECT 49.125 66.950 111.745 67.565 ;
        POLYGON 49.125 66.950 49.195 66.950 49.195 66.515 ;
        RECT 49.195 66.515 111.745 66.950 ;
        POLYGON 49.195 66.515 49.525 66.515 49.525 64.435 ;
        RECT 49.525 66.020 111.745 66.515 ;
        POLYGON 111.745 67.565 112.015 67.565 111.745 66.020 ;
        POLYGON 118.215 67.565 118.215 67.315 118.180 67.315 ;
        RECT 118.215 67.530 144.130 67.570 ;
        POLYGON 144.130 67.675 144.150 67.530 144.130 67.530 ;
        RECT 118.215 67.485 144.150 67.530 ;
        POLYGON 150.210 67.675 150.210 67.510 149.750 67.510 ;
        RECT 150.210 67.640 162.220 67.675 ;
        POLYGON 162.220 67.760 162.565 67.640 162.220 67.640 ;
        POLYGON 173.615 67.760 173.745 67.760 173.745 67.640 ;
        RECT 173.745 67.640 189.930 67.760 ;
        RECT 150.210 67.515 162.565 67.640 ;
        POLYGON 162.565 67.640 162.920 67.515 162.565 67.515 ;
        POLYGON 173.745 67.640 173.850 67.640 173.850 67.550 ;
        RECT 173.850 67.595 189.930 67.640 ;
        POLYGON 189.930 67.830 190.090 67.595 189.930 67.595 ;
        POLYGON 207.115 67.830 207.115 67.735 207.095 67.735 ;
        RECT 207.115 67.735 226.000 67.840 ;
        POLYGON 226.000 67.855 226.070 67.855 226.000 67.735 ;
        POLYGON 236.325 67.855 236.325 67.825 236.290 67.825 ;
        RECT 236.325 67.830 245.710 67.855 ;
        POLYGON 245.710 67.855 245.795 67.855 245.710 67.830 ;
        POLYGON 256.890 67.855 256.965 67.855 256.965 67.830 ;
        RECT 256.965 67.830 268.450 67.855 ;
        RECT 236.325 67.825 245.605 67.830 ;
        POLYGON 236.290 67.825 236.290 67.735 236.190 67.735 ;
        RECT 236.290 67.790 245.605 67.825 ;
        POLYGON 245.605 67.830 245.710 67.830 245.605 67.790 ;
        POLYGON 256.965 67.830 257.080 67.830 257.080 67.790 ;
        RECT 257.080 67.790 268.450 67.830 ;
        RECT 236.290 67.775 245.560 67.790 ;
        POLYGON 245.560 67.790 245.605 67.790 245.560 67.775 ;
        POLYGON 257.080 67.790 257.125 67.790 257.125 67.775 ;
        RECT 257.125 67.775 268.450 67.790 ;
        RECT 236.290 67.735 245.445 67.775 ;
        POLYGON 245.445 67.775 245.555 67.775 245.445 67.735 ;
        POLYGON 257.125 67.775 257.240 67.775 257.240 67.735 ;
        RECT 257.240 67.735 268.450 67.775 ;
        POLYGON 268.450 67.855 268.590 67.735 268.450 67.735 ;
        POLYGON 284.840 67.855 284.925 67.855 284.925 67.735 ;
        RECT 284.925 67.735 303.120 67.855 ;
        POLYGON 207.095 67.725 207.095 67.610 207.075 67.610 ;
        RECT 207.095 67.610 225.920 67.735 ;
        RECT 207.075 67.595 225.920 67.610 ;
        POLYGON 225.920 67.735 226.000 67.735 225.920 67.600 ;
        POLYGON 236.190 67.735 236.190 67.600 236.040 67.600 ;
        RECT 236.190 67.600 244.860 67.735 ;
        POLYGON 236.040 67.600 236.040 67.595 236.035 67.595 ;
        RECT 236.040 67.595 244.860 67.600 ;
        RECT 173.850 67.590 190.090 67.595 ;
        POLYGON 190.090 67.595 190.095 67.590 190.090 67.590 ;
        POLYGON 207.075 67.595 207.075 67.590 207.070 67.590 ;
        RECT 207.075 67.590 225.835 67.595 ;
        RECT 173.850 67.550 190.095 67.590 ;
        POLYGON 173.850 67.550 173.885 67.550 173.885 67.515 ;
        RECT 173.885 67.515 190.095 67.550 ;
        RECT 150.210 67.510 162.920 67.515 ;
        POLYGON 149.745 67.510 149.745 67.495 149.710 67.495 ;
        RECT 149.745 67.495 162.920 67.510 ;
        POLYGON 144.150 67.495 144.155 67.485 144.150 67.485 ;
        RECT 118.215 67.440 144.155 67.485 ;
        POLYGON 149.710 67.495 149.710 67.475 149.665 67.475 ;
        RECT 149.710 67.475 162.920 67.495 ;
        POLYGON 144.155 67.475 144.160 67.440 144.155 67.440 ;
        RECT 118.215 67.345 144.160 67.440 ;
        POLYGON 149.665 67.475 149.665 67.400 149.485 67.400 ;
        RECT 149.665 67.440 162.920 67.475 ;
        POLYGON 162.920 67.515 163.105 67.440 162.920 67.440 ;
        POLYGON 173.885 67.515 173.920 67.515 173.920 67.485 ;
        RECT 173.920 67.485 190.095 67.515 ;
        POLYGON 173.920 67.485 173.965 67.485 173.965 67.440 ;
        RECT 173.965 67.440 190.095 67.485 ;
        RECT 149.665 67.425 163.105 67.440 ;
        POLYGON 163.105 67.440 163.145 67.425 163.105 67.425 ;
        POLYGON 173.965 67.440 173.985 67.440 173.985 67.425 ;
        RECT 173.985 67.425 190.095 67.440 ;
        RECT 149.665 67.400 163.145 67.425 ;
        POLYGON 144.160 67.400 144.170 67.345 144.160 67.345 ;
        POLYGON 149.485 67.400 149.485 67.345 149.350 67.345 ;
        RECT 149.485 67.345 163.145 67.400 ;
        RECT 118.215 67.315 144.170 67.345 ;
        POLYGON 118.180 67.310 118.180 67.245 118.170 67.245 ;
        RECT 118.180 67.300 144.170 67.315 ;
        POLYGON 144.170 67.345 144.175 67.300 144.170 67.300 ;
        RECT 118.180 67.245 144.175 67.300 ;
        POLYGON 149.350 67.345 149.350 67.295 149.230 67.295 ;
        RECT 149.350 67.295 163.145 67.345 ;
        POLYGON 118.170 67.235 118.170 66.345 118.045 66.345 ;
        RECT 118.170 67.205 144.175 67.245 ;
        POLYGON 144.175 67.295 144.185 67.205 144.175 67.205 ;
        POLYGON 149.230 67.295 149.230 67.205 149.015 67.205 ;
        RECT 149.230 67.205 163.145 67.295 ;
        RECT 118.170 67.160 144.185 67.205 ;
        POLYGON 149.015 67.205 149.015 67.175 148.945 67.175 ;
        RECT 149.015 67.175 163.145 67.205 ;
        POLYGON 148.945 67.175 148.945 67.165 148.920 67.165 ;
        RECT 148.945 67.165 163.145 67.175 ;
        POLYGON 144.185 67.165 144.190 67.160 144.185 67.160 ;
        RECT 118.170 66.925 144.190 67.160 ;
        POLYGON 148.920 67.165 148.920 67.125 148.830 67.125 ;
        RECT 148.920 67.125 163.145 67.165 ;
        POLYGON 144.190 67.125 144.215 66.925 144.190 66.925 ;
        RECT 118.170 66.830 144.215 66.925 ;
        POLYGON 148.830 67.125 148.830 66.900 148.355 66.900 ;
        RECT 148.830 67.070 163.145 67.125 ;
        POLYGON 163.145 67.425 164.000 67.070 163.145 67.070 ;
        POLYGON 173.985 67.425 174.025 67.425 174.025 67.390 ;
        RECT 174.025 67.390 190.095 67.425 ;
        POLYGON 174.025 67.390 174.220 67.390 174.220 67.215 ;
        RECT 174.220 67.215 190.095 67.390 ;
        POLYGON 174.220 67.215 174.365 67.215 174.365 67.070 ;
        RECT 174.365 67.070 190.095 67.215 ;
        RECT 148.830 67.045 164.000 67.070 ;
        POLYGON 164.000 67.070 164.050 67.045 164.000 67.045 ;
        POLYGON 174.365 67.070 174.390 67.070 174.390 67.045 ;
        RECT 174.390 67.045 190.095 67.070 ;
        RECT 148.830 67.010 164.050 67.045 ;
        POLYGON 164.050 67.045 164.125 67.010 164.050 67.010 ;
        POLYGON 174.390 67.045 174.425 67.045 174.425 67.015 ;
        RECT 174.425 67.015 190.095 67.045 ;
        POLYGON 174.425 67.015 174.430 67.015 174.430 67.010 ;
        RECT 174.430 67.010 190.095 67.015 ;
        RECT 148.830 67.000 164.130 67.010 ;
        POLYGON 164.130 67.010 164.145 67.000 164.130 67.000 ;
        POLYGON 174.430 67.010 174.440 67.010 174.440 67.000 ;
        RECT 174.440 67.000 190.095 67.010 ;
        RECT 148.830 66.900 164.145 67.000 ;
        POLYGON 144.215 66.900 144.225 66.830 144.215 66.830 ;
        RECT 118.170 66.785 144.225 66.830 ;
        POLYGON 148.355 66.900 148.355 66.820 148.190 66.820 ;
        RECT 148.355 66.820 164.145 66.900 ;
        POLYGON 144.225 66.820 144.230 66.785 144.225 66.785 ;
        RECT 118.170 66.740 144.230 66.785 ;
        POLYGON 148.190 66.820 148.190 66.780 148.100 66.780 ;
        RECT 148.190 66.780 164.145 66.820 ;
        POLYGON 148.100 66.780 148.100 66.745 148.030 66.745 ;
        RECT 148.100 66.745 164.145 66.780 ;
        POLYGON 144.230 66.745 144.235 66.740 144.230 66.740 ;
        RECT 118.170 66.645 144.235 66.740 ;
        POLYGON 148.030 66.745 148.030 66.705 147.945 66.705 ;
        RECT 148.030 66.705 164.145 66.745 ;
        POLYGON 144.235 66.705 144.245 66.645 144.235 66.645 ;
        RECT 118.170 66.600 144.245 66.645 ;
        POLYGON 147.945 66.705 147.945 66.625 147.800 66.625 ;
        RECT 147.945 66.625 164.145 66.705 ;
        POLYGON 144.245 66.625 144.250 66.600 144.245 66.600 ;
        RECT 118.170 66.550 144.250 66.600 ;
        POLYGON 147.800 66.625 147.800 66.560 147.680 66.560 ;
        RECT 147.800 66.620 164.145 66.625 ;
        POLYGON 164.145 67.000 164.930 66.620 164.145 66.620 ;
        POLYGON 174.440 67.000 174.825 67.000 174.825 66.620 ;
        RECT 174.825 66.675 190.095 67.000 ;
        POLYGON 190.095 67.590 190.735 66.675 190.095 66.675 ;
        POLYGON 207.070 67.580 207.070 67.550 207.065 67.550 ;
        RECT 207.070 67.550 225.835 67.590 ;
        POLYGON 207.065 67.550 207.065 66.720 206.920 66.720 ;
        RECT 207.065 67.450 225.835 67.550 ;
        POLYGON 225.835 67.595 225.920 67.595 225.835 67.450 ;
        POLYGON 236.035 67.595 236.035 67.570 236.005 67.570 ;
        RECT 236.035 67.570 244.860 67.595 ;
        POLYGON 236.005 67.570 236.005 67.450 235.885 67.450 ;
        RECT 236.005 67.525 244.860 67.570 ;
        POLYGON 244.860 67.735 245.445 67.735 244.860 67.525 ;
        POLYGON 257.240 67.735 257.345 67.735 257.345 67.700 ;
        RECT 257.345 67.700 268.590 67.735 ;
        POLYGON 257.345 67.700 257.415 67.700 257.415 67.675 ;
        RECT 257.415 67.675 268.590 67.700 ;
        POLYGON 257.415 67.675 257.495 67.675 257.495 67.645 ;
        RECT 257.495 67.645 268.590 67.675 ;
        POLYGON 257.495 67.645 257.640 67.645 257.640 67.595 ;
        RECT 257.640 67.635 268.590 67.645 ;
        POLYGON 268.590 67.735 268.705 67.635 268.590 67.635 ;
        POLYGON 284.925 67.735 284.995 67.735 284.995 67.635 ;
        RECT 284.995 67.635 303.120 67.735 ;
        RECT 257.640 67.620 268.705 67.635 ;
        POLYGON 268.705 67.635 268.730 67.620 268.705 67.620 ;
        POLYGON 284.995 67.635 285.005 67.635 285.005 67.620 ;
        RECT 285.005 67.620 303.120 67.635 ;
        RECT 257.640 67.595 268.730 67.620 ;
        POLYGON 268.730 67.620 268.755 67.595 268.730 67.595 ;
        POLYGON 285.005 67.620 285.020 67.620 285.020 67.600 ;
        RECT 285.020 67.595 303.120 67.620 ;
        POLYGON 257.640 67.595 257.845 67.595 257.845 67.525 ;
        RECT 257.845 67.525 268.755 67.595 ;
        RECT 236.005 67.490 244.765 67.525 ;
        POLYGON 244.765 67.525 244.860 67.525 244.765 67.490 ;
        POLYGON 257.850 67.525 257.920 67.525 257.920 67.500 ;
        RECT 257.920 67.500 268.755 67.525 ;
        POLYGON 257.920 67.500 257.940 67.500 257.940 67.490 ;
        RECT 257.940 67.490 268.755 67.500 ;
        RECT 236.005 67.485 244.750 67.490 ;
        POLYGON 244.750 67.490 244.765 67.490 244.750 67.485 ;
        POLYGON 257.940 67.490 257.955 67.490 257.955 67.485 ;
        RECT 257.955 67.485 268.755 67.490 ;
        RECT 236.005 67.450 244.530 67.485 ;
        RECT 207.065 67.220 225.700 67.450 ;
        POLYGON 225.700 67.450 225.835 67.450 225.700 67.220 ;
        POLYGON 235.885 67.450 235.885 67.220 235.655 67.220 ;
        RECT 235.885 67.395 244.530 67.450 ;
        POLYGON 244.530 67.485 244.750 67.485 244.530 67.395 ;
        POLYGON 257.955 67.485 258.135 67.485 258.135 67.410 ;
        RECT 258.135 67.410 268.755 67.485 ;
        POLYGON 258.135 67.410 258.170 67.410 258.170 67.395 ;
        RECT 258.170 67.395 268.755 67.410 ;
        RECT 235.885 67.220 243.960 67.395 ;
        RECT 207.065 66.720 225.430 67.220 ;
        POLYGON 206.920 66.710 206.920 66.675 206.910 66.675 ;
        RECT 206.920 66.705 225.430 66.720 ;
        POLYGON 225.430 67.220 225.700 67.220 225.430 66.710 ;
        POLYGON 235.655 67.220 235.655 66.840 235.275 66.840 ;
        RECT 235.655 67.155 243.960 67.220 ;
        POLYGON 243.960 67.395 244.525 67.395 243.960 67.155 ;
        POLYGON 258.170 67.395 258.290 67.395 258.290 67.345 ;
        RECT 258.290 67.350 268.755 67.395 ;
        POLYGON 268.755 67.595 269.010 67.350 268.755 67.350 ;
        POLYGON 285.020 67.595 285.195 67.595 285.195 67.350 ;
        RECT 285.195 67.350 303.120 67.595 ;
        RECT 258.290 67.345 269.010 67.350 ;
        POLYGON 258.290 67.345 258.660 67.345 258.660 67.195 ;
        RECT 258.660 67.195 269.010 67.345 ;
        POLYGON 258.660 67.195 258.750 67.195 258.750 67.155 ;
        RECT 258.750 67.155 269.010 67.195 ;
        RECT 235.655 67.110 243.845 67.155 ;
        POLYGON 243.845 67.155 243.960 67.155 243.845 67.110 ;
        POLYGON 258.750 67.155 258.855 67.155 258.855 67.110 ;
        RECT 258.855 67.110 269.010 67.155 ;
        RECT 235.655 67.080 243.780 67.110 ;
        POLYGON 243.780 67.110 243.845 67.110 243.780 67.080 ;
        POLYGON 258.855 67.110 258.930 67.110 258.930 67.080 ;
        RECT 258.930 67.080 269.010 67.110 ;
        RECT 235.655 66.920 243.455 67.080 ;
        POLYGON 243.455 67.080 243.780 67.080 243.455 66.920 ;
        POLYGON 258.930 67.080 259.000 67.080 259.000 67.055 ;
        RECT 259.000 67.055 269.010 67.080 ;
        POLYGON 259.000 67.055 259.270 67.055 259.270 66.920 ;
        RECT 259.270 66.920 269.010 67.055 ;
        RECT 235.655 66.840 243.190 66.920 ;
        POLYGON 235.275 66.840 235.275 66.745 235.175 66.745 ;
        RECT 235.275 66.795 243.190 66.840 ;
        POLYGON 243.190 66.920 243.455 66.920 243.190 66.795 ;
        POLYGON 259.270 66.920 259.530 66.920 259.530 66.795 ;
        RECT 259.530 66.795 269.010 66.920 ;
        RECT 235.275 66.745 243.010 66.795 ;
        POLYGON 235.175 66.745 235.175 66.710 235.145 66.710 ;
        RECT 235.175 66.710 243.010 66.745 ;
        POLYGON 243.010 66.795 243.190 66.795 243.010 66.710 ;
        POLYGON 259.530 66.795 259.655 66.795 259.655 66.735 ;
        RECT 259.655 66.780 269.010 66.795 ;
        POLYGON 269.010 67.350 269.610 66.780 269.010 66.780 ;
        POLYGON 285.195 67.350 285.595 67.350 285.595 66.785 ;
        RECT 285.595 66.780 303.120 67.350 ;
        RECT 259.655 66.735 269.610 66.780 ;
        POLYGON 259.655 66.735 259.710 66.735 259.710 66.710 ;
        RECT 259.710 66.710 269.610 66.735 ;
        POLYGON 269.610 66.780 269.680 66.710 269.610 66.710 ;
        POLYGON 285.595 66.780 285.645 66.780 285.645 66.710 ;
        RECT 285.645 66.710 303.120 66.780 ;
        RECT 206.920 66.675 225.230 66.705 ;
        RECT 174.825 66.620 190.735 66.675 ;
        RECT 147.800 66.565 164.930 66.620 ;
        POLYGON 164.930 66.620 165.045 66.565 164.930 66.565 ;
        POLYGON 174.825 66.620 174.845 66.620 174.845 66.605 ;
        RECT 174.845 66.605 190.735 66.620 ;
        POLYGON 174.845 66.605 174.855 66.605 174.855 66.600 ;
        RECT 174.855 66.600 190.735 66.605 ;
        POLYGON 174.855 66.600 174.890 66.600 174.890 66.565 ;
        RECT 174.890 66.565 190.735 66.600 ;
        RECT 147.800 66.560 165.045 66.565 ;
        POLYGON 144.250 66.560 144.255 66.550 144.250 66.550 ;
        RECT 118.170 66.345 144.255 66.550 ;
        POLYGON 147.680 66.560 147.680 66.520 147.605 66.520 ;
        RECT 147.680 66.530 165.045 66.560 ;
        POLYGON 165.045 66.565 165.115 66.530 165.045 66.530 ;
        POLYGON 174.890 66.565 174.925 66.565 174.925 66.530 ;
        RECT 174.925 66.530 190.735 66.565 ;
        RECT 147.680 66.520 165.115 66.530 ;
        POLYGON 118.045 66.345 118.045 66.020 118.000 66.020 ;
        RECT 118.045 66.320 144.255 66.345 ;
        POLYGON 144.255 66.520 144.280 66.320 144.255 66.320 ;
        POLYGON 147.605 66.520 147.605 66.320 147.245 66.320 ;
        RECT 147.605 66.320 165.115 66.520 ;
        RECT 118.045 66.270 144.280 66.320 ;
        POLYGON 147.245 66.320 147.245 66.305 147.215 66.305 ;
        RECT 147.245 66.305 165.115 66.320 ;
        POLYGON 144.280 66.305 144.285 66.270 144.280 66.270 ;
        RECT 118.045 66.180 144.285 66.270 ;
        POLYGON 147.215 66.305 147.215 66.240 147.090 66.240 ;
        RECT 147.215 66.300 165.115 66.305 ;
        POLYGON 165.115 66.530 165.520 66.300 165.115 66.300 ;
        POLYGON 174.925 66.530 175.105 66.530 175.105 66.345 ;
        RECT 175.105 66.345 190.735 66.530 ;
        POLYGON 175.105 66.345 175.110 66.345 175.110 66.335 ;
        RECT 175.110 66.335 190.735 66.345 ;
        POLYGON 175.110 66.335 175.140 66.335 175.140 66.300 ;
        RECT 175.140 66.300 190.735 66.335 ;
        RECT 147.215 66.270 165.525 66.300 ;
        POLYGON 165.525 66.300 165.575 66.270 165.525 66.270 ;
        POLYGON 175.140 66.300 175.170 66.300 175.170 66.270 ;
        RECT 175.170 66.270 190.735 66.300 ;
        RECT 147.215 66.240 165.575 66.270 ;
        POLYGON 144.285 66.240 144.295 66.180 144.285 66.180 ;
        POLYGON 147.090 66.240 147.090 66.180 146.995 66.180 ;
        RECT 147.090 66.180 165.575 66.240 ;
        RECT 118.045 66.085 144.295 66.180 ;
        POLYGON 144.295 66.180 144.305 66.085 144.295 66.085 ;
        RECT 118.045 66.040 144.305 66.085 ;
        POLYGON 146.995 66.180 146.995 66.055 146.795 66.055 ;
        RECT 146.995 66.150 165.575 66.180 ;
        POLYGON 165.575 66.270 165.790 66.150 165.575 66.150 ;
        POLYGON 175.170 66.270 175.290 66.270 175.290 66.150 ;
        RECT 175.290 66.150 190.735 66.270 ;
        RECT 146.995 66.055 165.790 66.150 ;
        POLYGON 144.305 66.055 144.310 66.040 144.305 66.040 ;
        RECT 118.045 66.020 144.310 66.040 ;
        POLYGON 146.795 66.055 146.795 66.035 146.765 66.035 ;
        RECT 146.795 66.035 165.790 66.055 ;
        RECT 49.525 65.185 111.645 66.020 ;
        POLYGON 111.645 66.020 111.745 66.020 111.645 65.185 ;
        POLYGON 118.000 66.020 118.000 65.445 117.920 65.445 ;
        RECT 118.000 65.900 144.310 66.020 ;
        POLYGON 144.310 66.035 144.325 65.900 144.310 65.900 ;
        RECT 118.000 65.855 144.325 65.900 ;
        POLYGON 146.765 66.035 146.765 65.890 146.525 65.890 ;
        RECT 146.765 66.005 165.790 66.035 ;
        POLYGON 165.790 66.150 166.050 66.005 165.790 66.005 ;
        POLYGON 175.290 66.150 175.315 66.150 175.315 66.125 ;
        RECT 175.315 66.125 190.735 66.150 ;
        POLYGON 175.315 66.125 175.360 66.125 175.360 66.075 ;
        RECT 175.360 66.075 190.735 66.125 ;
        POLYGON 175.360 66.075 175.385 66.075 175.385 66.055 ;
        RECT 175.385 66.055 190.735 66.075 ;
        POLYGON 175.385 66.055 175.400 66.055 175.400 66.035 ;
        RECT 175.400 66.035 190.735 66.055 ;
        POLYGON 175.400 66.035 175.430 66.035 175.430 66.005 ;
        RECT 175.430 66.005 190.735 66.035 ;
        RECT 146.765 65.995 166.050 66.005 ;
        POLYGON 166.050 66.005 166.070 65.995 166.050 65.995 ;
        POLYGON 175.430 66.005 175.440 66.005 175.440 65.995 ;
        RECT 175.440 65.995 190.735 66.005 ;
        RECT 146.765 65.890 166.070 65.995 ;
        POLYGON 144.325 65.890 144.330 65.855 144.325 65.855 ;
        POLYGON 146.525 65.890 146.525 65.855 146.470 65.855 ;
        RECT 146.525 65.855 166.070 65.890 ;
        RECT 118.000 65.825 144.330 65.855 ;
        POLYGON 144.330 65.855 144.335 65.825 144.330 65.825 ;
        RECT 118.000 65.735 144.335 65.825 ;
        POLYGON 146.470 65.855 146.470 65.800 146.380 65.800 ;
        RECT 146.470 65.800 166.070 65.855 ;
        POLYGON 144.335 65.800 144.350 65.735 144.335 65.735 ;
        POLYGON 146.380 65.800 146.380 65.735 146.270 65.735 ;
        RECT 146.380 65.735 166.070 65.800 ;
        RECT 118.000 65.705 144.350 65.735 ;
        POLYGON 144.350 65.735 144.355 65.705 144.350 65.705 ;
        RECT 118.000 65.620 144.355 65.705 ;
        POLYGON 146.270 65.735 146.270 65.695 146.215 65.695 ;
        RECT 146.270 65.695 166.070 65.735 ;
        POLYGON 144.355 65.695 144.370 65.620 144.355 65.620 ;
        RECT 118.000 65.530 144.370 65.620 ;
        POLYGON 146.215 65.695 146.215 65.595 146.070 65.595 ;
        RECT 146.215 65.665 166.070 65.695 ;
        POLYGON 166.070 65.995 166.595 65.665 166.070 65.665 ;
        POLYGON 175.440 65.995 175.470 65.995 175.470 65.965 ;
        RECT 175.470 65.965 190.735 65.995 ;
        POLYGON 175.470 65.965 175.510 65.965 175.510 65.920 ;
        RECT 175.510 65.920 190.735 65.965 ;
        POLYGON 175.510 65.920 175.530 65.920 175.530 65.905 ;
        RECT 175.530 65.905 190.735 65.920 ;
        POLYGON 175.530 65.905 175.555 65.905 175.555 65.870 ;
        RECT 175.555 65.870 190.735 65.905 ;
        POLYGON 175.555 65.870 175.575 65.870 175.575 65.855 ;
        RECT 175.575 65.855 190.735 65.870 ;
        POLYGON 175.575 65.855 175.670 65.855 175.670 65.755 ;
        RECT 175.670 65.780 190.735 65.855 ;
        POLYGON 190.735 66.675 191.315 65.780 190.735 65.780 ;
        POLYGON 206.910 66.665 206.910 66.005 206.795 66.005 ;
        RECT 206.910 66.330 225.230 66.675 ;
        POLYGON 225.230 66.705 225.430 66.705 225.230 66.330 ;
        POLYGON 235.145 66.710 235.145 66.565 235.015 66.565 ;
        RECT 235.145 66.685 242.960 66.710 ;
        POLYGON 242.960 66.710 243.010 66.710 242.960 66.685 ;
        POLYGON 259.710 66.710 259.765 66.710 259.765 66.685 ;
        RECT 259.765 66.685 269.680 66.710 ;
        RECT 235.145 66.565 242.720 66.685 ;
        POLYGON 235.015 66.565 235.015 66.330 234.800 66.330 ;
        RECT 235.015 66.555 242.720 66.565 ;
        POLYGON 242.720 66.685 242.960 66.685 242.720 66.555 ;
        POLYGON 259.765 66.685 259.820 66.685 259.820 66.660 ;
        RECT 259.820 66.660 269.680 66.685 ;
        POLYGON 259.820 66.660 260.030 66.660 260.030 66.555 ;
        RECT 260.030 66.555 269.680 66.660 ;
        RECT 235.015 66.400 242.440 66.555 ;
        POLYGON 242.440 66.555 242.715 66.555 242.440 66.400 ;
        POLYGON 260.030 66.555 260.045 66.555 260.045 66.550 ;
        RECT 260.045 66.550 269.680 66.555 ;
        POLYGON 260.045 66.550 260.145 66.550 260.145 66.495 ;
        RECT 260.145 66.515 269.680 66.550 ;
        POLYGON 269.680 66.710 269.885 66.515 269.680 66.515 ;
        POLYGON 285.645 66.710 285.680 66.710 285.680 66.665 ;
        RECT 285.680 66.665 303.120 66.710 ;
        POLYGON 285.680 66.665 285.775 66.665 285.775 66.515 ;
        RECT 285.775 66.515 303.120 66.665 ;
        RECT 260.145 66.495 269.885 66.515 ;
        POLYGON 260.145 66.495 260.310 66.495 260.310 66.400 ;
        RECT 260.310 66.400 269.885 66.495 ;
        RECT 235.015 66.370 242.385 66.400 ;
        POLYGON 242.385 66.400 242.440 66.400 242.385 66.370 ;
        POLYGON 260.310 66.400 260.365 66.400 260.365 66.370 ;
        RECT 260.365 66.370 269.885 66.400 ;
        RECT 235.015 66.330 242.110 66.370 ;
        RECT 206.910 66.325 225.225 66.330 ;
        POLYGON 225.225 66.330 225.230 66.330 225.225 66.325 ;
        POLYGON 234.800 66.330 234.800 66.325 234.795 66.325 ;
        RECT 234.800 66.325 242.110 66.330 ;
        RECT 206.910 66.005 224.970 66.325 ;
        POLYGON 206.795 66.005 206.795 65.795 206.770 65.795 ;
        RECT 206.795 65.795 224.970 66.005 ;
        POLYGON 224.970 66.325 225.225 66.325 224.970 65.795 ;
        POLYGON 234.795 66.320 234.795 65.865 234.380 65.865 ;
        RECT 234.795 66.220 242.110 66.325 ;
        POLYGON 242.110 66.370 242.380 66.370 242.110 66.220 ;
        POLYGON 260.365 66.370 260.385 66.370 260.385 66.360 ;
        RECT 260.385 66.360 269.885 66.370 ;
        POLYGON 260.385 66.360 260.635 66.360 260.635 66.220 ;
        RECT 260.635 66.220 269.885 66.360 ;
        RECT 234.795 65.980 241.710 66.220 ;
        POLYGON 241.710 66.220 242.110 66.220 241.710 65.980 ;
        POLYGON 260.635 66.220 260.970 66.220 260.970 66.035 ;
        RECT 260.970 66.035 269.885 66.220 ;
        POLYGON 260.970 66.035 261.050 66.035 261.050 65.990 ;
        RECT 261.050 65.990 269.885 66.035 ;
        POLYGON 261.050 65.990 261.065 65.990 261.065 65.980 ;
        RECT 261.065 65.980 269.885 65.990 ;
        RECT 234.795 65.960 241.680 65.980 ;
        POLYGON 241.680 65.980 241.710 65.980 241.680 65.960 ;
        POLYGON 261.070 65.980 261.100 65.980 261.100 65.960 ;
        RECT 261.100 65.960 269.885 65.980 ;
        RECT 234.795 65.865 241.390 65.960 ;
        POLYGON 234.380 65.865 234.380 65.795 234.320 65.795 ;
        RECT 234.380 65.795 241.390 65.865 ;
        RECT 206.770 65.780 224.965 65.795 ;
        POLYGON 224.965 65.795 224.970 65.795 224.965 65.785 ;
        POLYGON 234.320 65.790 234.320 65.785 234.315 65.785 ;
        RECT 234.320 65.785 241.390 65.795 ;
        POLYGON 234.315 65.785 234.315 65.780 234.310 65.780 ;
        RECT 234.315 65.780 241.390 65.785 ;
        POLYGON 241.390 65.960 241.680 65.960 241.390 65.780 ;
        POLYGON 261.100 65.960 261.380 65.960 261.380 65.780 ;
        RECT 261.380 65.825 269.885 65.960 ;
        POLYGON 269.885 66.515 270.555 65.825 269.885 65.825 ;
        POLYGON 285.775 66.515 286.220 66.515 286.220 65.825 ;
        RECT 286.220 65.825 303.120 66.515 ;
        RECT 261.380 65.795 270.555 65.825 ;
        POLYGON 270.555 65.825 270.585 65.795 270.555 65.795 ;
        POLYGON 286.220 65.825 286.235 65.825 286.235 65.800 ;
        RECT 286.235 65.795 303.120 65.825 ;
        RECT 261.380 65.780 270.585 65.795 ;
        POLYGON 270.585 65.795 270.595 65.780 270.585 65.780 ;
        POLYGON 286.235 65.795 286.245 65.795 286.245 65.785 ;
        RECT 286.245 65.780 303.120 65.795 ;
        RECT 175.670 65.755 191.315 65.780 ;
        POLYGON 175.670 65.755 175.685 65.755 175.685 65.740 ;
        RECT 175.685 65.740 191.315 65.755 ;
        POLYGON 175.685 65.740 175.700 65.740 175.700 65.720 ;
        RECT 175.700 65.720 191.315 65.740 ;
        POLYGON 175.700 65.720 175.750 65.720 175.750 65.665 ;
        RECT 175.750 65.665 191.315 65.720 ;
        RECT 146.215 65.640 166.595 65.665 ;
        POLYGON 166.595 65.665 166.630 65.640 166.595 65.640 ;
        POLYGON 175.750 65.665 175.775 65.665 175.775 65.640 ;
        RECT 175.775 65.640 191.315 65.665 ;
        RECT 146.215 65.595 166.630 65.640 ;
        POLYGON 144.370 65.595 144.385 65.530 144.370 65.530 ;
        RECT 118.000 65.500 144.385 65.530 ;
        POLYGON 146.065 65.595 146.065 65.515 145.945 65.515 ;
        RECT 146.065 65.515 166.630 65.595 ;
        POLYGON 144.385 65.515 144.390 65.500 144.385 65.500 ;
        RECT 118.000 65.445 144.390 65.500 ;
        POLYGON 145.945 65.515 145.945 65.490 145.910 65.490 ;
        RECT 145.945 65.490 166.630 65.515 ;
        POLYGON 144.390 65.490 144.400 65.445 144.390 65.445 ;
        POLYGON 117.920 65.435 117.920 65.190 117.885 65.190 ;
        RECT 117.920 65.295 144.400 65.445 ;
        POLYGON 145.910 65.490 145.910 65.435 145.830 65.435 ;
        RECT 145.910 65.435 166.630 65.490 ;
        POLYGON 144.400 65.435 144.425 65.295 144.400 65.295 ;
        RECT 117.920 65.240 144.425 65.295 ;
        POLYGON 145.830 65.435 145.830 65.290 145.625 65.290 ;
        RECT 145.830 65.410 166.630 65.435 ;
        POLYGON 166.630 65.640 166.995 65.410 166.630 65.410 ;
        POLYGON 175.775 65.640 175.970 65.640 175.970 65.440 ;
        RECT 175.970 65.440 191.315 65.640 ;
        POLYGON 175.970 65.440 175.995 65.440 175.995 65.410 ;
        RECT 175.995 65.415 191.315 65.440 ;
        POLYGON 191.315 65.780 191.550 65.415 191.315 65.415 ;
        POLYGON 206.770 65.780 206.770 65.455 206.730 65.455 ;
        RECT 206.770 65.455 224.785 65.780 ;
        POLYGON 206.730 65.450 206.730 65.415 206.725 65.415 ;
        RECT 206.730 65.420 224.785 65.455 ;
        POLYGON 224.785 65.780 224.965 65.780 224.785 65.420 ;
        POLYGON 234.310 65.780 234.310 65.420 234.010 65.420 ;
        RECT 234.310 65.720 241.290 65.780 ;
        POLYGON 241.290 65.780 241.390 65.780 241.290 65.720 ;
        POLYGON 261.380 65.780 261.475 65.780 261.475 65.720 ;
        RECT 261.475 65.720 270.595 65.780 ;
        RECT 234.310 65.525 241.010 65.720 ;
        POLYGON 241.010 65.720 241.290 65.720 241.010 65.525 ;
        POLYGON 261.475 65.720 261.760 65.720 261.760 65.540 ;
        RECT 261.760 65.540 270.595 65.720 ;
        POLYGON 261.760 65.540 261.780 65.540 261.780 65.525 ;
        RECT 261.780 65.525 270.595 65.540 ;
        RECT 234.310 65.450 240.900 65.525 ;
        POLYGON 240.900 65.525 241.010 65.525 240.900 65.450 ;
        POLYGON 261.780 65.525 261.900 65.525 261.900 65.450 ;
        RECT 261.900 65.450 270.595 65.525 ;
        POLYGON 270.595 65.780 270.915 65.450 270.595 65.450 ;
        POLYGON 286.245 65.780 286.460 65.780 286.460 65.450 ;
        RECT 286.460 65.450 303.120 65.780 ;
        RECT 234.310 65.420 240.660 65.450 ;
        RECT 206.730 65.415 224.575 65.420 ;
        RECT 175.995 65.410 191.550 65.415 ;
        POLYGON 191.550 65.415 191.555 65.410 191.550 65.410 ;
        RECT 145.830 65.390 166.995 65.410 ;
        POLYGON 166.995 65.410 167.020 65.390 166.995 65.390 ;
        POLYGON 175.995 65.410 176.010 65.410 176.010 65.390 ;
        RECT 176.010 65.390 191.555 65.410 ;
        RECT 145.830 65.310 167.020 65.390 ;
        POLYGON 167.020 65.390 167.135 65.310 167.020 65.310 ;
        POLYGON 176.010 65.390 176.080 65.390 176.080 65.310 ;
        RECT 176.080 65.310 191.555 65.390 ;
        RECT 145.830 65.290 167.135 65.310 ;
        POLYGON 144.425 65.290 144.435 65.240 144.425 65.240 ;
        RECT 117.920 65.210 144.435 65.240 ;
        POLYGON 145.625 65.290 145.625 65.225 145.530 65.225 ;
        RECT 145.625 65.230 167.135 65.290 ;
        RECT 145.625 65.225 155.500 65.230 ;
        POLYGON 155.500 65.230 155.635 65.230 155.500 65.225 ;
        POLYGON 155.995 65.230 156.160 65.230 156.160 65.225 ;
        RECT 156.160 65.225 167.135 65.230 ;
        POLYGON 144.435 65.225 144.440 65.210 144.435 65.210 ;
        RECT 117.920 65.190 144.440 65.210 ;
        RECT 49.525 64.415 111.460 65.185 ;
        POLYGON 49.525 64.415 49.800 64.415 49.800 62.710 ;
        RECT 49.800 63.625 111.460 64.415 ;
        POLYGON 111.460 65.185 111.645 65.185 111.460 63.625 ;
        POLYGON 117.885 65.185 117.885 64.800 117.830 64.800 ;
        RECT 117.885 65.120 144.440 65.190 ;
        POLYGON 145.530 65.225 145.530 65.185 145.470 65.185 ;
        RECT 145.530 65.200 154.920 65.225 ;
        POLYGON 154.920 65.225 155.475 65.225 154.920 65.200 ;
        POLYGON 156.480 65.225 156.505 65.225 156.505 65.220 ;
        RECT 156.505 65.220 167.135 65.225 ;
        POLYGON 156.555 65.220 156.815 65.220 156.815 65.200 ;
        RECT 156.815 65.200 167.135 65.220 ;
        RECT 145.530 65.195 154.780 65.200 ;
        POLYGON 154.780 65.200 154.865 65.200 154.780 65.195 ;
        POLYGON 156.815 65.200 156.880 65.200 156.880 65.195 ;
        RECT 156.880 65.195 167.135 65.200 ;
        RECT 145.530 65.185 154.410 65.195 ;
        POLYGON 144.440 65.185 144.455 65.120 144.440 65.120 ;
        POLYGON 145.470 65.185 145.470 65.120 145.385 65.120 ;
        RECT 145.470 65.160 154.410 65.185 ;
        POLYGON 154.410 65.195 154.770 65.195 154.410 65.160 ;
        POLYGON 156.880 65.195 156.950 65.195 156.950 65.190 ;
        RECT 156.950 65.190 167.135 65.195 ;
        POLYGON 156.975 65.190 157.100 65.190 157.100 65.180 ;
        RECT 157.100 65.180 167.135 65.190 ;
        POLYGON 157.105 65.180 157.265 65.180 157.265 65.170 ;
        RECT 157.265 65.170 167.135 65.180 ;
        POLYGON 157.270 65.170 157.370 65.170 157.370 65.165 ;
        RECT 157.370 65.165 167.135 65.170 ;
        POLYGON 157.370 65.165 157.405 65.165 157.405 65.160 ;
        RECT 157.405 65.160 167.135 65.165 ;
        RECT 145.470 65.125 154.045 65.160 ;
        POLYGON 154.045 65.160 154.405 65.160 154.045 65.125 ;
        POLYGON 157.405 65.160 157.640 65.160 157.640 65.130 ;
        RECT 157.640 65.130 167.135 65.160 ;
        POLYGON 157.640 65.130 157.700 65.130 157.700 65.125 ;
        RECT 157.700 65.125 167.135 65.130 ;
        RECT 145.470 65.120 154.000 65.125 ;
        POLYGON 154.000 65.125 154.045 65.125 154.000 65.120 ;
        POLYGON 157.710 65.125 157.745 65.125 157.745 65.120 ;
        RECT 157.745 65.120 167.135 65.125 ;
        RECT 117.885 64.915 144.455 65.120 ;
        POLYGON 144.455 65.120 144.490 64.915 144.455 64.915 ;
        RECT 117.885 64.890 144.490 64.915 ;
        POLYGON 145.385 65.120 145.385 64.900 145.100 64.900 ;
        RECT 145.385 65.115 153.925 65.120 ;
        POLYGON 153.925 65.120 153.995 65.120 153.925 65.115 ;
        POLYGON 157.745 65.120 157.785 65.120 157.785 65.115 ;
        RECT 157.785 65.115 167.135 65.120 ;
        RECT 145.385 65.110 153.900 65.115 ;
        POLYGON 153.900 65.115 153.925 65.115 153.900 65.110 ;
        POLYGON 157.785 65.115 157.825 65.115 157.825 65.110 ;
        RECT 157.825 65.110 167.135 65.115 ;
        RECT 145.385 65.035 153.425 65.110 ;
        POLYGON 153.425 65.110 153.895 65.110 153.425 65.035 ;
        POLYGON 157.825 65.110 158.020 65.110 158.020 65.085 ;
        RECT 158.020 65.085 167.135 65.110 ;
        POLYGON 158.020 65.085 158.170 65.085 158.170 65.065 ;
        RECT 158.170 65.080 167.135 65.085 ;
        POLYGON 167.135 65.310 167.455 65.080 167.135 65.080 ;
        POLYGON 176.080 65.310 176.285 65.310 176.285 65.080 ;
        RECT 176.285 65.080 191.555 65.310 ;
        RECT 158.170 65.065 167.455 65.080 ;
        POLYGON 158.170 65.065 158.235 65.065 158.235 65.060 ;
        RECT 158.235 65.060 167.455 65.065 ;
        POLYGON 158.235 65.060 158.370 65.060 158.370 65.035 ;
        RECT 158.370 65.035 167.455 65.060 ;
        RECT 145.385 65.025 153.340 65.035 ;
        POLYGON 153.340 65.035 153.395 65.035 153.340 65.025 ;
        POLYGON 158.370 65.035 158.430 65.035 158.430 65.025 ;
        RECT 158.430 65.025 167.455 65.035 ;
        RECT 145.385 64.985 153.075 65.025 ;
        POLYGON 153.075 65.025 153.335 65.025 153.075 64.985 ;
        POLYGON 158.435 65.025 158.660 65.025 158.660 64.985 ;
        RECT 158.660 64.985 167.455 65.025 ;
        RECT 145.385 64.950 152.905 64.985 ;
        POLYGON 152.905 64.985 153.075 64.985 152.905 64.950 ;
        POLYGON 158.660 64.985 158.690 64.985 158.690 64.980 ;
        RECT 158.690 64.980 167.455 64.985 ;
        POLYGON 158.690 64.980 158.750 64.980 158.750 64.965 ;
        RECT 158.750 64.965 167.455 64.980 ;
        POLYGON 158.755 64.965 158.840 64.965 158.840 64.950 ;
        RECT 158.840 64.950 167.455 64.965 ;
        RECT 145.385 64.940 152.860 64.950 ;
        POLYGON 152.860 64.950 152.900 64.950 152.860 64.940 ;
        POLYGON 158.840 64.950 158.895 64.950 158.895 64.940 ;
        RECT 158.895 64.940 167.455 64.950 ;
        RECT 145.385 64.900 152.645 64.940 ;
        POLYGON 144.490 64.900 144.495 64.890 144.490 64.890 ;
        POLYGON 145.100 64.900 145.100 64.890 145.085 64.890 ;
        RECT 145.100 64.895 152.645 64.900 ;
        POLYGON 152.645 64.940 152.855 64.940 152.645 64.895 ;
        POLYGON 158.895 64.940 159.095 64.940 159.095 64.905 ;
        RECT 159.095 64.905 167.455 64.940 ;
        POLYGON 159.095 64.905 159.140 64.905 159.140 64.895 ;
        RECT 159.140 64.895 167.455 64.905 ;
        RECT 145.100 64.890 152.415 64.895 ;
        RECT 117.885 64.800 144.495 64.890 ;
        POLYGON 144.495 64.890 144.510 64.800 144.495 64.800 ;
        POLYGON 117.830 64.795 117.830 64.510 117.790 64.510 ;
        RECT 117.830 64.710 144.510 64.800 ;
        POLYGON 145.085 64.890 145.085 64.775 144.935 64.775 ;
        RECT 145.085 64.845 152.415 64.890 ;
        POLYGON 152.415 64.895 152.640 64.895 152.415 64.845 ;
        POLYGON 159.145 64.895 159.195 64.895 159.195 64.880 ;
        RECT 159.195 64.880 167.455 64.895 ;
        POLYGON 159.200 64.880 159.355 64.880 159.355 64.845 ;
        RECT 159.355 64.845 167.455 64.880 ;
        RECT 145.085 64.820 152.290 64.845 ;
        POLYGON 152.290 64.845 152.415 64.845 152.290 64.820 ;
        POLYGON 159.355 64.845 159.470 64.845 159.470 64.820 ;
        RECT 159.470 64.820 167.455 64.845 ;
        RECT 145.085 64.810 152.235 64.820 ;
        POLYGON 152.235 64.820 152.290 64.820 152.235 64.810 ;
        POLYGON 159.470 64.820 159.510 64.820 159.510 64.810 ;
        RECT 159.510 64.810 167.455 64.820 ;
        RECT 145.085 64.775 151.970 64.810 ;
        POLYGON 144.510 64.775 144.525 64.710 144.510 64.710 ;
        POLYGON 144.935 64.775 144.935 64.710 144.850 64.710 ;
        RECT 144.935 64.740 151.970 64.775 ;
        POLYGON 151.970 64.810 152.235 64.810 151.970 64.740 ;
        POLYGON 159.510 64.810 159.695 64.810 159.695 64.765 ;
        RECT 159.695 64.765 167.455 64.810 ;
        POLYGON 159.700 64.765 159.800 64.765 159.800 64.740 ;
        RECT 159.800 64.740 167.455 64.765 ;
        RECT 144.935 64.730 151.935 64.740 ;
        POLYGON 151.935 64.740 151.965 64.740 151.935 64.730 ;
        POLYGON 159.800 64.740 159.840 64.740 159.840 64.730 ;
        RECT 159.840 64.730 167.455 64.740 ;
        RECT 144.935 64.710 151.735 64.730 ;
        RECT 117.830 64.680 144.525 64.710 ;
        POLYGON 144.525 64.710 144.530 64.680 144.525 64.680 ;
        RECT 117.830 64.620 144.530 64.680 ;
        POLYGON 144.850 64.710 144.850 64.675 144.805 64.675 ;
        RECT 144.850 64.675 151.735 64.710 ;
        POLYGON 151.735 64.730 151.935 64.730 151.735 64.675 ;
        POLYGON 159.845 64.730 159.950 64.730 159.950 64.705 ;
        RECT 159.950 64.720 167.455 64.730 ;
        POLYGON 167.455 65.080 167.950 64.720 167.455 64.720 ;
        POLYGON 176.285 65.080 176.600 65.080 176.600 64.720 ;
        RECT 176.600 64.720 191.555 65.080 ;
        RECT 159.950 64.705 167.950 64.720 ;
        POLYGON 159.950 64.705 160.050 64.705 160.050 64.675 ;
        RECT 160.050 64.675 167.950 64.705 ;
        POLYGON 144.805 64.675 144.805 64.670 144.800 64.670 ;
        RECT 144.805 64.670 151.465 64.675 ;
        POLYGON 144.530 64.670 144.540 64.620 144.530 64.620 ;
        POLYGON 144.800 64.670 144.800 64.620 144.740 64.620 ;
        RECT 144.800 64.620 151.465 64.670 ;
        RECT 117.830 64.590 144.540 64.620 ;
        POLYGON 144.740 64.620 144.740 64.605 144.720 64.605 ;
        RECT 144.740 64.605 151.465 64.620 ;
        POLYGON 151.465 64.675 151.735 64.675 151.465 64.605 ;
        POLYGON 160.050 64.675 160.155 64.675 160.155 64.645 ;
        RECT 160.155 64.645 167.950 64.675 ;
        POLYGON 160.155 64.645 160.185 64.645 160.185 64.635 ;
        RECT 160.185 64.635 167.950 64.645 ;
        POLYGON 160.185 64.635 160.285 64.635 160.285 64.605 ;
        RECT 160.285 64.605 167.950 64.635 ;
        POLYGON 144.540 64.605 144.545 64.590 144.540 64.590 ;
        RECT 117.830 64.535 144.545 64.590 ;
        POLYGON 144.720 64.605 144.720 64.580 144.690 64.580 ;
        RECT 144.720 64.590 151.410 64.605 ;
        POLYGON 151.410 64.605 151.465 64.605 151.410 64.590 ;
        POLYGON 160.285 64.605 160.335 64.605 160.335 64.590 ;
        RECT 160.335 64.590 167.950 64.605 ;
        RECT 144.720 64.580 151.320 64.590 ;
        POLYGON 144.545 64.580 144.555 64.535 144.545 64.535 ;
        RECT 117.830 64.510 144.555 64.535 ;
        POLYGON 144.685 64.580 144.685 64.530 144.625 64.530 ;
        RECT 144.685 64.560 151.320 64.580 ;
        POLYGON 151.320 64.590 151.410 64.590 151.320 64.560 ;
        POLYGON 160.335 64.590 160.435 64.590 160.435 64.560 ;
        RECT 160.435 64.560 167.950 64.590 ;
        RECT 144.685 64.530 151.180 64.560 ;
        POLYGON 144.625 64.530 144.625 64.510 144.605 64.510 ;
        RECT 144.625 64.515 151.180 64.530 ;
        POLYGON 151.180 64.560 151.320 64.560 151.180 64.515 ;
        POLYGON 160.435 64.560 160.520 64.560 160.520 64.535 ;
        RECT 160.520 64.535 167.950 64.560 ;
        POLYGON 160.520 64.535 160.590 64.535 160.590 64.515 ;
        RECT 160.590 64.515 167.950 64.535 ;
        RECT 144.625 64.510 150.995 64.515 ;
        POLYGON 117.790 64.500 117.790 64.400 117.775 64.400 ;
        RECT 117.790 64.485 144.555 64.510 ;
        POLYGON 144.555 64.510 144.560 64.485 144.555 64.485 ;
        POLYGON 144.605 64.510 144.605 64.485 144.575 64.485 ;
        RECT 144.605 64.485 150.995 64.510 ;
        RECT 117.790 64.470 144.560 64.485 ;
        POLYGON 144.575 64.485 144.575 64.470 144.560 64.470 ;
        RECT 144.575 64.470 150.995 64.485 ;
        RECT 117.790 64.455 150.995 64.470 ;
        POLYGON 150.995 64.515 151.180 64.515 150.995 64.455 ;
        POLYGON 160.590 64.515 160.665 64.515 160.665 64.495 ;
        RECT 160.665 64.495 167.950 64.515 ;
        POLYGON 160.665 64.495 160.795 64.495 160.795 64.455 ;
        RECT 160.795 64.475 167.950 64.495 ;
        POLYGON 167.950 64.720 168.255 64.475 167.950 64.475 ;
        POLYGON 176.600 64.720 176.670 64.720 176.670 64.640 ;
        RECT 176.670 64.640 191.555 64.720 ;
        RECT 160.795 64.455 168.255 64.475 ;
        POLYGON 176.670 64.640 176.815 64.640 176.815 64.470 ;
        RECT 176.815 64.470 191.555 64.640 ;
        RECT 117.790 64.400 150.635 64.455 ;
        POLYGON 117.775 64.400 117.775 63.625 117.720 63.625 ;
        RECT 117.775 64.335 150.635 64.400 ;
        POLYGON 150.635 64.455 150.995 64.455 150.635 64.335 ;
        POLYGON 160.795 64.455 160.830 64.455 160.830 64.440 ;
        RECT 160.830 64.440 168.255 64.455 ;
        POLYGON 160.830 64.440 161.130 64.440 161.130 64.335 ;
        RECT 161.130 64.335 168.255 64.440 ;
        RECT 117.775 64.325 150.600 64.335 ;
        POLYGON 150.600 64.335 150.635 64.335 150.600 64.325 ;
        POLYGON 161.130 64.335 161.150 64.335 161.150 64.325 ;
        RECT 161.150 64.325 168.255 64.335 ;
        RECT 117.775 64.300 150.540 64.325 ;
        POLYGON 150.540 64.325 150.600 64.325 150.540 64.300 ;
        POLYGON 161.150 64.325 161.175 64.325 161.175 64.315 ;
        RECT 161.175 64.320 168.255 64.325 ;
        POLYGON 168.255 64.470 168.445 64.320 168.255 64.320 ;
        POLYGON 176.815 64.470 176.940 64.470 176.940 64.325 ;
        RECT 176.940 64.320 191.555 64.470 ;
        RECT 161.175 64.315 168.445 64.320 ;
        POLYGON 161.175 64.315 161.215 64.315 161.215 64.300 ;
        RECT 161.215 64.300 168.445 64.315 ;
        RECT 117.775 64.130 150.095 64.300 ;
        POLYGON 150.095 64.300 150.540 64.300 150.095 64.130 ;
        POLYGON 161.215 64.300 161.485 64.300 161.485 64.205 ;
        RECT 161.485 64.205 168.445 64.300 ;
        POLYGON 161.485 64.205 161.585 64.205 161.585 64.170 ;
        RECT 161.585 64.170 168.445 64.205 ;
        POLYGON 161.585 64.170 161.635 64.170 161.635 64.150 ;
        RECT 161.635 64.150 168.445 64.170 ;
        POLYGON 161.635 64.150 161.680 64.150 161.680 64.130 ;
        RECT 161.680 64.130 168.445 64.150 ;
        RECT 117.775 64.125 150.090 64.130 ;
        POLYGON 150.090 64.130 150.095 64.130 150.090 64.125 ;
        POLYGON 161.680 64.130 161.695 64.130 161.695 64.125 ;
        RECT 161.695 64.125 168.445 64.130 ;
        RECT 117.775 64.015 149.805 64.125 ;
        POLYGON 149.805 64.125 150.090 64.125 149.805 64.015 ;
        POLYGON 161.695 64.125 161.805 64.125 161.805 64.080 ;
        RECT 161.805 64.080 168.445 64.125 ;
        POLYGON 161.805 64.080 161.955 64.080 161.955 64.015 ;
        RECT 161.955 64.015 168.445 64.080 ;
        RECT 117.775 63.990 149.750 64.015 ;
        POLYGON 149.750 64.015 149.805 64.015 149.750 63.990 ;
        POLYGON 161.955 64.015 162.010 64.015 162.010 63.990 ;
        RECT 162.010 63.995 168.445 64.015 ;
        POLYGON 168.445 64.320 168.840 63.995 168.445 63.995 ;
        POLYGON 176.940 64.320 177.200 64.320 177.200 63.995 ;
        RECT 177.200 64.105 191.555 64.320 ;
        POLYGON 191.555 65.410 192.330 64.105 191.555 64.105 ;
        POLYGON 206.725 65.410 206.725 64.150 206.575 64.150 ;
        RECT 206.725 64.940 224.575 65.415 ;
        POLYGON 224.575 65.420 224.785 65.420 224.575 64.940 ;
        POLYGON 234.010 65.415 234.010 65.260 233.880 65.260 ;
        RECT 234.010 65.290 240.660 65.420 ;
        POLYGON 240.660 65.450 240.900 65.450 240.660 65.290 ;
        POLYGON 261.900 65.450 261.950 65.450 261.950 65.420 ;
        RECT 261.950 65.420 270.915 65.450 ;
        POLYGON 261.950 65.420 262.020 65.420 262.020 65.375 ;
        RECT 262.020 65.375 270.915 65.420 ;
        POLYGON 262.020 65.375 262.115 65.375 262.115 65.310 ;
        RECT 262.115 65.360 270.915 65.375 ;
        POLYGON 270.915 65.450 271.005 65.360 270.915 65.360 ;
        POLYGON 286.460 65.450 286.515 65.450 286.515 65.365 ;
        RECT 286.515 65.360 303.120 65.450 ;
        RECT 262.115 65.310 271.005 65.360 ;
        POLYGON 262.115 65.310 262.140 65.310 262.140 65.290 ;
        RECT 262.140 65.290 271.005 65.310 ;
        RECT 234.010 65.260 240.505 65.290 ;
        POLYGON 233.880 65.260 233.880 65.130 233.775 65.130 ;
        RECT 233.880 65.180 240.505 65.260 ;
        POLYGON 240.505 65.290 240.660 65.290 240.505 65.180 ;
        POLYGON 262.140 65.290 262.195 65.290 262.195 65.250 ;
        RECT 262.195 65.250 271.005 65.290 ;
        POLYGON 250.620 65.250 250.620 65.245 250.525 65.245 ;
        POLYGON 250.620 65.250 250.855 65.245 250.620 65.245 ;
        POLYGON 262.195 65.250 262.200 65.250 262.200 65.245 ;
        RECT 262.200 65.245 271.005 65.250 ;
        POLYGON 250.495 65.245 250.495 65.220 249.925 65.220 ;
        RECT 250.495 65.240 251.245 65.245 ;
        POLYGON 251.245 65.245 251.480 65.240 251.245 65.240 ;
        POLYGON 262.200 65.245 262.205 65.245 262.205 65.240 ;
        RECT 262.205 65.240 271.005 65.245 ;
        RECT 250.495 65.225 251.480 65.240 ;
        POLYGON 251.480 65.240 251.655 65.225 251.480 65.225 ;
        POLYGON 262.205 65.240 262.225 65.240 262.225 65.225 ;
        RECT 262.225 65.225 271.005 65.240 ;
        RECT 250.495 65.220 251.655 65.225 ;
        POLYGON 249.920 65.220 249.920 65.215 249.785 65.215 ;
        RECT 249.920 65.215 251.655 65.220 ;
        POLYGON 249.760 65.215 249.760 65.180 249.395 65.180 ;
        RECT 249.760 65.205 251.655 65.215 ;
        POLYGON 251.655 65.225 251.975 65.205 251.655 65.205 ;
        POLYGON 262.225 65.225 262.255 65.225 262.255 65.205 ;
        RECT 262.255 65.205 271.005 65.225 ;
        RECT 249.760 65.200 251.985 65.205 ;
        POLYGON 251.985 65.205 252.075 65.200 251.985 65.200 ;
        POLYGON 262.255 65.205 262.260 65.205 262.260 65.200 ;
        RECT 262.260 65.200 271.005 65.205 ;
        RECT 249.760 65.180 252.080 65.200 ;
        POLYGON 252.080 65.200 252.340 65.180 252.080 65.180 ;
        POLYGON 262.260 65.200 262.290 65.200 262.290 65.180 ;
        RECT 262.290 65.180 271.005 65.200 ;
        RECT 233.880 65.130 240.335 65.180 ;
        POLYGON 233.775 65.130 233.775 64.945 233.620 64.945 ;
        RECT 233.775 65.050 240.335 65.130 ;
        POLYGON 240.335 65.180 240.505 65.180 240.335 65.050 ;
        POLYGON 249.395 65.180 249.395 65.175 249.345 65.175 ;
        RECT 249.395 65.175 252.340 65.180 ;
        POLYGON 249.345 65.175 249.345 65.145 249.060 65.145 ;
        RECT 249.345 65.145 252.340 65.175 ;
        POLYGON 249.055 65.145 249.055 65.130 248.905 65.130 ;
        RECT 249.055 65.135 252.340 65.145 ;
        POLYGON 252.340 65.180 252.710 65.135 252.340 65.135 ;
        POLYGON 262.290 65.180 262.350 65.180 262.350 65.135 ;
        RECT 262.350 65.135 271.005 65.180 ;
        RECT 249.055 65.130 252.715 65.135 ;
        POLYGON 248.905 65.130 248.905 65.120 248.840 65.120 ;
        RECT 248.905 65.120 252.715 65.130 ;
        POLYGON 252.715 65.135 252.815 65.120 252.715 65.120 ;
        POLYGON 262.350 65.135 262.370 65.135 262.370 65.120 ;
        RECT 262.370 65.120 271.005 65.135 ;
        POLYGON 248.840 65.120 248.840 65.050 248.410 65.050 ;
        RECT 248.840 65.080 252.820 65.120 ;
        POLYGON 252.820 65.120 253.155 65.080 252.820 65.080 ;
        POLYGON 262.370 65.120 262.405 65.120 262.405 65.095 ;
        RECT 262.405 65.095 271.005 65.120 ;
        POLYGON 262.405 65.095 262.425 65.095 262.425 65.080 ;
        RECT 262.425 65.080 271.005 65.095 ;
        RECT 248.840 65.075 253.155 65.080 ;
        POLYGON 253.155 65.080 253.195 65.075 253.155 65.075 ;
        POLYGON 262.425 65.080 262.430 65.080 262.430 65.075 ;
        RECT 262.430 65.075 271.005 65.080 ;
        RECT 248.840 65.050 253.195 65.075 ;
        RECT 233.775 64.990 240.255 65.050 ;
        POLYGON 240.255 65.050 240.335 65.050 240.255 64.990 ;
        POLYGON 248.410 65.050 248.410 65.040 248.350 65.040 ;
        RECT 248.410 65.040 253.195 65.050 ;
        POLYGON 248.345 65.040 248.345 65.020 248.205 65.020 ;
        RECT 248.345 65.030 253.195 65.040 ;
        POLYGON 253.195 65.075 253.440 65.030 253.195 65.030 ;
        POLYGON 262.430 65.075 262.495 65.075 262.495 65.030 ;
        RECT 262.495 65.030 271.005 65.075 ;
        RECT 248.345 65.020 253.440 65.030 ;
        POLYGON 248.200 65.020 248.200 64.995 248.055 64.995 ;
        RECT 248.200 64.995 253.440 65.020 ;
        POLYGON 248.055 64.995 248.055 64.990 248.030 64.990 ;
        RECT 248.055 64.990 253.440 64.995 ;
        RECT 233.775 64.945 239.760 64.990 ;
        POLYGON 233.620 64.945 233.620 64.940 233.615 64.940 ;
        RECT 233.620 64.940 239.760 64.945 ;
        RECT 206.725 64.490 224.375 64.940 ;
        POLYGON 224.375 64.940 224.575 64.940 224.375 64.490 ;
        POLYGON 233.615 64.940 233.615 64.490 233.285 64.490 ;
        RECT 233.615 64.605 239.760 64.940 ;
        POLYGON 239.760 64.990 240.255 64.990 239.760 64.605 ;
        POLYGON 248.030 64.990 248.030 64.935 247.760 64.935 ;
        RECT 248.030 64.935 253.440 64.990 ;
        POLYGON 247.760 64.935 247.760 64.910 247.655 64.910 ;
        RECT 247.760 64.930 253.440 64.935 ;
        POLYGON 253.440 65.030 253.985 64.930 253.440 64.930 ;
        POLYGON 262.495 65.030 262.635 65.030 262.635 64.930 ;
        RECT 262.635 64.930 271.005 65.030 ;
        RECT 247.760 64.920 253.990 64.930 ;
        POLYGON 253.990 64.930 254.045 64.920 253.990 64.920 ;
        POLYGON 262.635 64.930 262.650 64.930 262.650 64.920 ;
        RECT 262.650 64.920 271.005 64.930 ;
        RECT 247.760 64.910 254.045 64.920 ;
        POLYGON 247.655 64.910 247.655 64.815 247.210 64.815 ;
        RECT 247.655 64.895 254.045 64.910 ;
        POLYGON 254.045 64.920 254.150 64.895 254.045 64.895 ;
        POLYGON 262.650 64.920 262.685 64.920 262.685 64.895 ;
        RECT 262.685 64.895 271.005 64.920 ;
        RECT 247.655 64.880 254.150 64.895 ;
        POLYGON 254.150 64.895 254.220 64.880 254.150 64.880 ;
        POLYGON 262.685 64.895 262.705 64.895 262.705 64.880 ;
        RECT 262.705 64.880 271.005 64.895 ;
        RECT 247.655 64.815 254.225 64.880 ;
        POLYGON 247.210 64.815 247.210 64.780 247.075 64.780 ;
        RECT 247.210 64.780 254.225 64.815 ;
        POLYGON 247.070 64.780 247.070 64.755 246.980 64.755 ;
        RECT 247.070 64.755 254.225 64.780 ;
        POLYGON 246.980 64.755 246.980 64.670 246.685 64.670 ;
        RECT 246.980 64.730 254.225 64.755 ;
        POLYGON 254.225 64.880 254.850 64.730 254.225 64.730 ;
        POLYGON 262.705 64.880 262.770 64.880 262.770 64.835 ;
        RECT 262.770 64.835 271.005 64.880 ;
        POLYGON 262.770 64.835 262.915 64.835 262.915 64.730 ;
        RECT 262.915 64.810 271.005 64.835 ;
        POLYGON 271.005 65.360 271.490 64.810 271.005 64.810 ;
        POLYGON 286.515 65.360 286.610 65.360 286.610 65.220 ;
        RECT 286.610 65.220 303.120 65.360 ;
        POLYGON 286.610 65.220 286.850 65.220 286.850 64.815 ;
        RECT 286.850 64.810 303.120 65.220 ;
        RECT 262.915 64.730 271.490 64.810 ;
        RECT 246.980 64.720 254.850 64.730 ;
        POLYGON 254.850 64.730 254.885 64.720 254.850 64.720 ;
        POLYGON 262.915 64.730 262.925 64.730 262.925 64.720 ;
        RECT 262.925 64.720 271.490 64.730 ;
        RECT 246.980 64.670 254.885 64.720 ;
        POLYGON 246.680 64.670 246.680 64.605 246.450 64.605 ;
        RECT 246.680 64.640 254.885 64.670 ;
        POLYGON 254.885 64.720 255.155 64.640 254.885 64.640 ;
        POLYGON 262.925 64.720 262.950 64.720 262.950 64.705 ;
        RECT 262.950 64.705 271.490 64.720 ;
        POLYGON 262.950 64.705 263.020 64.705 263.020 64.650 ;
        RECT 263.020 64.650 271.490 64.705 ;
        POLYGON 263.020 64.650 263.030 64.650 263.030 64.640 ;
        RECT 263.030 64.640 271.490 64.650 ;
        RECT 246.680 64.605 255.160 64.640 ;
        RECT 233.615 64.550 239.690 64.605 ;
        POLYGON 239.690 64.605 239.760 64.605 239.690 64.550 ;
        POLYGON 246.450 64.605 246.450 64.585 246.380 64.585 ;
        RECT 246.450 64.600 255.160 64.605 ;
        POLYGON 255.160 64.640 255.295 64.600 255.160 64.600 ;
        POLYGON 263.030 64.640 263.075 64.640 263.075 64.600 ;
        RECT 263.075 64.600 271.490 64.640 ;
        RECT 246.450 64.585 255.295 64.600 ;
        POLYGON 246.375 64.585 246.375 64.550 246.270 64.550 ;
        RECT 246.375 64.550 255.295 64.585 ;
        RECT 233.615 64.535 239.670 64.550 ;
        POLYGON 239.670 64.550 239.690 64.550 239.670 64.535 ;
        POLYGON 246.270 64.550 246.270 64.535 246.225 64.535 ;
        RECT 246.270 64.535 255.295 64.550 ;
        RECT 233.615 64.490 239.615 64.535 ;
        RECT 206.725 64.290 224.295 64.490 ;
        POLYGON 224.295 64.490 224.375 64.490 224.295 64.290 ;
        POLYGON 233.285 64.490 233.285 64.290 233.140 64.290 ;
        RECT 233.285 64.485 239.615 64.490 ;
        POLYGON 239.615 64.535 239.670 64.535 239.615 64.485 ;
        POLYGON 246.225 64.535 246.225 64.485 246.080 64.485 ;
        RECT 246.225 64.530 255.295 64.535 ;
        POLYGON 255.295 64.600 255.525 64.530 255.295 64.530 ;
        POLYGON 263.075 64.600 263.145 64.600 263.145 64.545 ;
        RECT 263.145 64.545 271.490 64.600 ;
        POLYGON 263.145 64.545 263.160 64.545 263.160 64.530 ;
        RECT 263.160 64.530 271.490 64.545 ;
        RECT 246.225 64.485 255.525 64.530 ;
        RECT 233.285 64.290 239.225 64.485 ;
        RECT 206.725 64.150 224.240 64.290 ;
        POLYGON 224.240 64.290 224.295 64.290 224.240 64.150 ;
        POLYGON 233.140 64.290 233.140 64.150 233.040 64.150 ;
        RECT 233.140 64.150 239.225 64.290 ;
        POLYGON 239.225 64.485 239.615 64.485 239.225 64.150 ;
        POLYGON 246.080 64.485 246.080 64.445 245.960 64.445 ;
        RECT 246.080 64.475 255.525 64.485 ;
        POLYGON 255.525 64.530 255.720 64.475 255.525 64.475 ;
        POLYGON 263.160 64.530 263.230 64.530 263.230 64.475 ;
        RECT 263.230 64.475 271.490 64.530 ;
        RECT 246.080 64.445 255.720 64.475 ;
        POLYGON 245.960 64.445 245.960 64.360 245.710 64.360 ;
        RECT 245.960 64.360 255.720 64.445 ;
        POLYGON 245.710 64.360 245.710 64.310 245.560 64.310 ;
        RECT 245.710 64.310 255.720 64.360 ;
        POLYGON 255.720 64.475 256.180 64.310 255.720 64.310 ;
        POLYGON 263.230 64.475 263.240 64.475 263.240 64.470 ;
        RECT 263.240 64.470 271.490 64.475 ;
        POLYGON 263.240 64.470 263.430 64.470 263.430 64.310 ;
        RECT 263.430 64.310 271.490 64.470 ;
        POLYGON 245.555 64.310 245.555 64.150 245.165 64.150 ;
        RECT 245.555 64.260 256.180 64.310 ;
        POLYGON 256.180 64.310 256.325 64.260 256.180 64.260 ;
        POLYGON 263.430 64.310 263.495 64.310 263.495 64.260 ;
        RECT 263.495 64.260 271.490 64.310 ;
        RECT 245.555 64.245 256.330 64.260 ;
        POLYGON 256.330 64.260 256.360 64.245 256.330 64.245 ;
        POLYGON 263.495 64.260 263.510 64.260 263.510 64.245 ;
        RECT 263.510 64.245 271.490 64.260 ;
        RECT 245.555 64.180 256.360 64.245 ;
        POLYGON 256.360 64.245 256.540 64.180 256.360 64.180 ;
        POLYGON 263.510 64.245 263.600 64.245 263.600 64.180 ;
        RECT 263.600 64.190 271.490 64.245 ;
        POLYGON 271.490 64.810 272.045 64.190 271.490 64.190 ;
        POLYGON 286.850 64.810 287.165 64.810 287.165 64.280 ;
        RECT 287.165 64.280 303.120 64.810 ;
        POLYGON 287.165 64.280 287.215 64.280 287.215 64.195 ;
        RECT 287.215 64.190 303.120 64.280 ;
        RECT 263.600 64.180 272.045 64.190 ;
        RECT 245.555 64.150 256.540 64.180 ;
        POLYGON 256.540 64.180 256.610 64.150 256.540 64.150 ;
        POLYGON 263.600 64.180 263.635 64.180 263.635 64.150 ;
        RECT 263.635 64.150 272.045 64.180 ;
        POLYGON 272.045 64.190 272.075 64.150 272.045 64.150 ;
        POLYGON 287.215 64.190 287.240 64.190 287.240 64.155 ;
        RECT 287.240 64.150 303.120 64.190 ;
        POLYGON 206.575 64.145 206.575 64.105 206.570 64.105 ;
        RECT 206.575 64.105 224.200 64.150 ;
        RECT 177.200 63.995 192.330 64.105 ;
        RECT 162.010 63.990 168.840 63.995 ;
        RECT 117.775 63.945 149.650 63.990 ;
        POLYGON 149.650 63.990 149.750 63.990 149.650 63.945 ;
        POLYGON 162.010 63.990 162.025 63.990 162.025 63.985 ;
        RECT 162.025 63.985 168.840 63.990 ;
        POLYGON 162.025 63.985 162.120 63.985 162.120 63.945 ;
        RECT 162.120 63.945 168.840 63.985 ;
        RECT 117.775 63.905 149.565 63.945 ;
        POLYGON 149.565 63.945 149.650 63.945 149.565 63.905 ;
        POLYGON 162.120 63.945 162.210 63.945 162.210 63.905 ;
        RECT 162.210 63.905 168.840 63.945 ;
        RECT 117.775 63.750 149.220 63.905 ;
        POLYGON 149.220 63.905 149.565 63.905 149.220 63.750 ;
        POLYGON 162.210 63.905 162.455 63.905 162.455 63.800 ;
        RECT 162.455 63.810 168.840 63.905 ;
        POLYGON 168.840 63.995 169.045 63.810 168.840 63.810 ;
        POLYGON 177.200 63.995 177.210 63.995 177.210 63.985 ;
        RECT 177.210 63.985 192.330 63.995 ;
        POLYGON 177.210 63.985 177.345 63.985 177.345 63.810 ;
        RECT 177.345 63.920 192.330 63.985 ;
        POLYGON 192.330 64.105 192.435 63.920 192.330 63.920 ;
        POLYGON 206.570 64.105 206.570 63.975 206.555 63.975 ;
        RECT 206.570 64.045 224.200 64.105 ;
        POLYGON 224.200 64.150 224.240 64.150 224.200 64.045 ;
        POLYGON 233.040 64.150 233.040 64.045 232.965 64.045 ;
        RECT 233.040 64.065 239.125 64.150 ;
        POLYGON 239.125 64.150 239.225 64.150 239.125 64.065 ;
        POLYGON 245.165 64.150 245.165 64.065 244.960 64.065 ;
        RECT 245.165 64.070 256.610 64.150 ;
        POLYGON 256.610 64.150 256.805 64.070 256.610 64.070 ;
        POLYGON 263.635 64.150 263.730 64.150 263.730 64.070 ;
        RECT 263.730 64.070 272.075 64.150 ;
        RECT 245.165 64.065 256.805 64.070 ;
        RECT 233.040 64.045 239.045 64.065 ;
        RECT 206.570 63.975 224.170 64.045 ;
        RECT 206.555 63.960 224.170 63.975 ;
        POLYGON 224.170 64.045 224.200 64.045 224.170 63.965 ;
        POLYGON 232.965 64.045 232.965 63.970 232.910 63.970 ;
        RECT 232.965 64.000 239.045 64.045 ;
        POLYGON 239.045 64.065 239.125 64.065 239.045 64.000 ;
        POLYGON 244.960 64.065 244.960 64.025 244.860 64.025 ;
        RECT 244.960 64.025 256.805 64.065 ;
        POLYGON 244.860 64.025 244.860 64.000 244.800 64.000 ;
        RECT 244.860 64.000 256.805 64.025 ;
        RECT 232.965 63.970 239.000 64.000 ;
        POLYGON 232.910 63.970 232.910 63.965 232.905 63.965 ;
        RECT 232.910 63.965 239.000 63.970 ;
        RECT 232.905 63.960 239.000 63.965 ;
        POLYGON 239.000 64.000 239.045 64.000 239.000 63.960 ;
        POLYGON 244.800 64.000 244.800 63.985 244.765 63.985 ;
        RECT 244.800 63.985 256.805 64.000 ;
        POLYGON 244.765 63.985 244.765 63.980 244.750 63.980 ;
        RECT 244.765 63.980 256.805 63.985 ;
        POLYGON 244.750 63.980 244.750 63.960 244.710 63.960 ;
        RECT 244.750 63.960 256.805 63.980 ;
        POLYGON 256.805 64.070 257.065 63.960 256.805 63.960 ;
        POLYGON 263.730 64.070 263.820 64.070 263.820 64.000 ;
        RECT 263.820 64.000 272.075 64.070 ;
        POLYGON 263.820 64.000 263.860 64.000 263.860 63.960 ;
        RECT 263.860 63.960 272.075 64.000 ;
        POLYGON 272.075 64.150 272.235 63.960 272.075 63.960 ;
        POLYGON 287.240 64.150 287.285 64.150 287.285 64.080 ;
        RECT 287.285 64.080 303.120 64.150 ;
        POLYGON 287.285 64.080 287.290 64.080 287.290 64.070 ;
        RECT 287.290 64.060 303.120 64.080 ;
        POLYGON 287.290 64.060 287.295 64.060 287.295 64.045 ;
        RECT 287.295 64.045 303.120 64.060 ;
        POLYGON 287.295 64.045 287.305 64.045 287.305 63.960 ;
        POLYGON 206.555 63.960 206.555 63.935 206.550 63.935 ;
        RECT 206.555 63.935 224.150 63.960 ;
        RECT 177.345 63.910 192.435 63.920 ;
        POLYGON 192.435 63.920 192.440 63.910 192.435 63.910 ;
        POLYGON 206.550 63.915 206.550 63.910 206.545 63.910 ;
        RECT 206.550 63.910 224.150 63.935 ;
        POLYGON 224.150 63.960 224.170 63.960 224.150 63.915 ;
        POLYGON 232.905 63.960 232.905 63.920 232.875 63.920 ;
        RECT 232.905 63.920 238.955 63.960 ;
        RECT 232.875 63.915 238.955 63.920 ;
        POLYGON 238.955 63.960 239.000 63.960 238.955 63.915 ;
        POLYGON 244.710 63.960 244.710 63.915 244.615 63.915 ;
        RECT 244.710 63.915 257.065 63.960 ;
        POLYGON 257.065 63.960 257.175 63.915 257.065 63.915 ;
        POLYGON 263.860 63.960 263.910 63.960 263.910 63.915 ;
        RECT 263.910 63.915 272.235 63.960 ;
        POLYGON 272.235 63.960 272.270 63.915 272.235 63.915 ;
        RECT 287.305 63.920 303.120 64.045 ;
        POLYGON 287.305 63.920 287.310 63.920 287.310 63.915 ;
        RECT 177.345 63.810 192.440 63.910 ;
        RECT 162.455 63.800 169.045 63.810 ;
        POLYGON 162.460 63.800 162.560 63.800 162.560 63.750 ;
        RECT 162.560 63.750 169.045 63.800 ;
        RECT 117.775 63.665 149.040 63.750 ;
        POLYGON 149.040 63.750 149.220 63.750 149.040 63.665 ;
        POLYGON 162.560 63.750 162.730 63.750 162.730 63.665 ;
        RECT 162.730 63.665 169.045 63.750 ;
        RECT 117.775 63.625 148.830 63.665 ;
        RECT 49.800 63.015 111.390 63.625 ;
        POLYGON 111.390 63.625 111.460 63.625 111.390 63.015 ;
        POLYGON 117.720 63.625 117.720 63.015 117.675 63.015 ;
        RECT 117.720 63.555 148.830 63.625 ;
        POLYGON 148.830 63.665 149.030 63.665 148.830 63.555 ;
        POLYGON 162.730 63.665 162.740 63.665 162.740 63.660 ;
        RECT 162.740 63.660 169.045 63.665 ;
        POLYGON 162.740 63.660 162.880 63.660 162.880 63.595 ;
        RECT 162.880 63.595 169.045 63.660 ;
        POLYGON 162.880 63.595 162.915 63.595 162.915 63.575 ;
        RECT 162.915 63.575 169.045 63.595 ;
        POLYGON 162.920 63.575 162.955 63.575 162.955 63.555 ;
        RECT 162.955 63.555 169.045 63.575 ;
        RECT 117.720 63.540 148.800 63.555 ;
        POLYGON 148.800 63.555 148.830 63.555 148.800 63.540 ;
        POLYGON 162.955 63.555 162.985 63.555 162.985 63.540 ;
        RECT 162.985 63.540 169.045 63.555 ;
        RECT 117.720 63.395 148.520 63.540 ;
        POLYGON 148.520 63.540 148.800 63.540 148.520 63.395 ;
        POLYGON 162.985 63.540 163.275 63.540 163.275 63.395 ;
        RECT 163.275 63.510 169.045 63.540 ;
        POLYGON 169.045 63.810 169.375 63.510 169.045 63.510 ;
        POLYGON 177.345 63.810 177.580 63.810 177.580 63.515 ;
        RECT 177.580 63.655 192.440 63.810 ;
        POLYGON 192.440 63.910 192.580 63.655 192.440 63.655 ;
        POLYGON 206.545 63.890 206.545 63.685 206.520 63.685 ;
        RECT 206.545 63.830 224.120 63.910 ;
        POLYGON 224.120 63.910 224.150 63.910 224.120 63.830 ;
        POLYGON 232.875 63.915 232.875 63.830 232.815 63.830 ;
        RECT 232.875 63.830 238.715 63.915 ;
        RECT 206.545 63.685 224.065 63.830 ;
        POLYGON 224.065 63.830 224.120 63.830 224.065 63.690 ;
        POLYGON 232.815 63.830 232.815 63.695 232.725 63.695 ;
        RECT 232.815 63.695 238.715 63.830 ;
        POLYGON 232.725 63.690 232.725 63.685 232.720 63.685 ;
        RECT 232.725 63.685 238.715 63.695 ;
        POLYGON 238.715 63.915 238.955 63.915 238.715 63.685 ;
        POLYGON 244.615 63.915 244.615 63.875 244.530 63.875 ;
        RECT 244.615 63.875 257.175 63.915 ;
        POLYGON 244.525 63.875 244.525 63.685 244.125 63.685 ;
        RECT 244.525 63.845 257.175 63.875 ;
        POLYGON 257.175 63.915 257.345 63.845 257.175 63.845 ;
        POLYGON 263.910 63.915 263.985 63.915 263.985 63.845 ;
        RECT 263.985 63.845 272.270 63.915 ;
        RECT 244.525 63.770 257.345 63.845 ;
        POLYGON 257.345 63.845 257.495 63.770 257.345 63.770 ;
        POLYGON 263.985 63.845 264.070 63.845 264.070 63.770 ;
        RECT 264.070 63.835 272.270 63.845 ;
        POLYGON 272.270 63.915 272.340 63.835 272.270 63.835 ;
        RECT 287.310 63.910 303.120 63.920 ;
        POLYGON 287.310 63.910 287.315 63.910 287.315 63.865 ;
        RECT 287.315 63.835 303.120 63.910 ;
        RECT 264.070 63.770 272.340 63.835 ;
        RECT 244.525 63.685 257.495 63.770 ;
        POLYGON 257.495 63.770 257.670 63.685 257.495 63.685 ;
        POLYGON 264.070 63.770 264.105 63.770 264.105 63.740 ;
        RECT 264.105 63.740 272.340 63.770 ;
        POLYGON 264.105 63.740 264.160 63.740 264.160 63.685 ;
        RECT 264.160 63.685 272.340 63.740 ;
        POLYGON 272.340 63.835 272.460 63.685 272.340 63.685 ;
        POLYGON 287.315 63.835 287.330 63.835 287.330 63.735 ;
        RECT 287.330 63.735 303.120 63.835 ;
        POLYGON 287.330 63.735 287.335 63.735 287.335 63.685 ;
        POLYGON 206.520 63.680 206.520 63.655 206.515 63.655 ;
        RECT 206.520 63.655 223.855 63.685 ;
        RECT 177.580 63.510 192.580 63.655 ;
        RECT 163.275 63.395 169.375 63.510 ;
        RECT 117.720 63.325 148.390 63.395 ;
        POLYGON 148.390 63.395 148.520 63.395 148.390 63.325 ;
        POLYGON 163.275 63.395 163.285 63.395 163.285 63.390 ;
        RECT 163.285 63.390 169.375 63.395 ;
        POLYGON 163.285 63.390 163.345 63.390 163.345 63.355 ;
        RECT 163.345 63.355 169.375 63.390 ;
        POLYGON 163.350 63.355 163.400 63.355 163.400 63.325 ;
        RECT 163.400 63.325 169.375 63.355 ;
        RECT 117.720 63.265 148.280 63.325 ;
        POLYGON 148.280 63.325 148.390 63.325 148.280 63.265 ;
        POLYGON 163.400 63.325 163.505 63.325 163.505 63.265 ;
        RECT 163.505 63.265 169.375 63.325 ;
        RECT 117.720 63.105 148.010 63.265 ;
        POLYGON 148.010 63.265 148.280 63.265 148.010 63.105 ;
        POLYGON 163.505 63.265 163.680 63.265 163.680 63.165 ;
        RECT 163.680 63.220 169.375 63.265 ;
        POLYGON 169.375 63.510 169.690 63.220 169.375 63.220 ;
        POLYGON 177.580 63.510 177.810 63.510 177.810 63.220 ;
        RECT 177.810 63.220 192.580 63.510 ;
        RECT 163.680 63.165 169.690 63.220 ;
        POLYGON 163.685 63.165 163.790 63.165 163.790 63.105 ;
        RECT 163.790 63.105 169.690 63.165 ;
        RECT 117.720 63.095 147.995 63.105 ;
        POLYGON 147.995 63.105 148.010 63.105 147.995 63.095 ;
        POLYGON 163.790 63.105 163.805 63.105 163.805 63.095 ;
        RECT 163.805 63.095 169.690 63.105 ;
        RECT 117.720 63.065 147.945 63.095 ;
        POLYGON 147.945 63.095 147.995 63.095 147.945 63.065 ;
        POLYGON 163.805 63.095 163.860 63.095 163.860 63.065 ;
        RECT 163.860 63.090 169.690 63.095 ;
        POLYGON 169.690 63.220 169.820 63.090 169.690 63.090 ;
        POLYGON 177.810 63.220 177.840 63.220 177.840 63.185 ;
        RECT 177.840 63.185 192.580 63.220 ;
        POLYGON 177.840 63.185 177.900 63.185 177.900 63.095 ;
        RECT 177.900 63.090 192.580 63.185 ;
        RECT 163.860 63.065 169.820 63.090 ;
        RECT 117.720 63.015 147.605 63.065 ;
        RECT 49.800 62.710 111.320 63.015 ;
        POLYGON 49.800 62.710 49.890 62.710 49.890 62.290 ;
        RECT 49.890 62.290 111.320 62.710 ;
        RECT 23.000 60.000 45.000 62.000 ;
        POLYGON 49.890 62.290 50.380 62.290 50.380 60.015 ;
        RECT 50.380 61.950 111.320 62.290 ;
        POLYGON 111.320 63.015 111.390 63.015 111.320 61.950 ;
        POLYGON 117.675 62.990 117.675 62.570 117.645 62.570 ;
        RECT 117.675 62.860 147.605 63.015 ;
        POLYGON 147.605 63.065 147.945 63.065 147.605 62.860 ;
        POLYGON 163.860 63.065 163.940 63.065 163.940 63.020 ;
        RECT 163.940 63.030 169.820 63.065 ;
        POLYGON 169.820 63.090 169.875 63.030 169.820 63.030 ;
        POLYGON 177.900 63.090 177.945 63.090 177.945 63.030 ;
        RECT 177.945 63.030 192.580 63.090 ;
        RECT 163.940 63.020 169.875 63.030 ;
        POLYGON 163.940 63.020 163.995 63.020 163.995 62.985 ;
        RECT 163.995 62.985 169.875 63.020 ;
        POLYGON 164.000 62.985 164.050 62.985 164.050 62.955 ;
        RECT 164.050 62.955 169.875 62.985 ;
        POLYGON 155.430 62.955 155.430 62.945 154.915 62.945 ;
        RECT 155.430 62.945 155.685 62.955 ;
        POLYGON 155.685 62.955 155.995 62.945 155.685 62.945 ;
        POLYGON 164.050 62.955 164.060 62.955 164.060 62.950 ;
        RECT 164.060 62.950 169.875 62.955 ;
        POLYGON 164.060 62.950 164.065 62.950 164.065 62.945 ;
        RECT 164.065 62.945 169.875 62.950 ;
        POLYGON 154.855 62.945 154.855 62.940 154.785 62.940 ;
        RECT 154.855 62.940 155.995 62.945 ;
        POLYGON 154.780 62.940 154.780 62.935 154.770 62.935 ;
        RECT 154.780 62.935 155.995 62.940 ;
        POLYGON 155.995 62.945 156.230 62.935 155.995 62.935 ;
        POLYGON 164.065 62.945 164.080 62.945 164.080 62.935 ;
        RECT 164.080 62.935 169.875 62.945 ;
        POLYGON 154.765 62.935 154.765 62.915 154.405 62.915 ;
        RECT 154.765 62.920 156.240 62.935 ;
        POLYGON 156.240 62.935 156.480 62.920 156.240 62.920 ;
        POLYGON 164.080 62.935 164.100 62.935 164.100 62.920 ;
        RECT 164.100 62.920 169.875 62.935 ;
        RECT 154.765 62.915 156.505 62.920 ;
        POLYGON 156.505 62.920 156.555 62.915 156.505 62.915 ;
        POLYGON 164.100 62.920 164.110 62.920 164.110 62.915 ;
        RECT 164.110 62.915 169.875 62.920 ;
        POLYGON 154.405 62.915 154.405 62.880 154.045 62.880 ;
        RECT 154.405 62.880 156.555 62.915 ;
        POLYGON 154.045 62.880 154.045 62.875 154.000 62.875 ;
        RECT 154.045 62.875 156.555 62.880 ;
        POLYGON 156.555 62.915 156.965 62.875 156.555 62.875 ;
        POLYGON 164.110 62.915 164.170 62.915 164.170 62.875 ;
        RECT 164.170 62.875 169.875 62.915 ;
        POLYGON 153.995 62.875 153.995 62.865 153.930 62.865 ;
        RECT 153.995 62.865 156.975 62.875 ;
        POLYGON 156.975 62.875 157.105 62.865 156.975 62.865 ;
        POLYGON 164.170 62.875 164.185 62.875 164.185 62.865 ;
        RECT 164.185 62.865 169.875 62.875 ;
        POLYGON 153.895 62.865 153.895 62.860 153.860 62.860 ;
        RECT 153.895 62.860 157.105 62.865 ;
        RECT 117.675 62.825 147.550 62.860 ;
        POLYGON 147.550 62.860 147.605 62.860 147.550 62.825 ;
        POLYGON 153.860 62.860 153.860 62.825 153.625 62.825 ;
        RECT 153.860 62.840 157.105 62.860 ;
        POLYGON 157.105 62.865 157.270 62.840 157.105 62.840 ;
        POLYGON 164.185 62.865 164.225 62.865 164.225 62.840 ;
        RECT 164.225 62.840 169.875 62.865 ;
        RECT 153.860 62.830 157.270 62.840 ;
        POLYGON 157.270 62.840 157.365 62.830 157.270 62.830 ;
        POLYGON 164.225 62.840 164.240 62.840 164.240 62.830 ;
        RECT 164.240 62.830 169.875 62.840 ;
        RECT 153.860 62.825 157.370 62.830 ;
        RECT 117.675 62.800 147.510 62.825 ;
        POLYGON 147.510 62.825 147.550 62.825 147.510 62.800 ;
        POLYGON 153.625 62.825 153.625 62.800 153.460 62.800 ;
        RECT 153.625 62.800 157.370 62.825 ;
        RECT 117.675 62.610 147.230 62.800 ;
        POLYGON 147.230 62.800 147.510 62.800 147.230 62.610 ;
        POLYGON 153.460 62.800 153.460 62.795 153.425 62.795 ;
        RECT 153.460 62.795 157.370 62.800 ;
        POLYGON 153.395 62.795 153.395 62.780 153.340 62.780 ;
        RECT 153.395 62.790 157.370 62.795 ;
        POLYGON 157.370 62.830 157.640 62.790 157.370 62.790 ;
        POLYGON 164.240 62.830 164.300 62.830 164.300 62.790 ;
        RECT 164.300 62.790 169.875 62.830 ;
        RECT 153.395 62.780 157.640 62.790 ;
        POLYGON 157.640 62.790 157.705 62.780 157.640 62.780 ;
        POLYGON 164.300 62.790 164.315 62.790 164.315 62.780 ;
        RECT 164.315 62.780 169.875 62.790 ;
        POLYGON 153.335 62.780 153.335 62.735 153.075 62.735 ;
        RECT 153.335 62.735 157.710 62.780 ;
        POLYGON 153.075 62.735 153.075 62.700 152.905 62.700 ;
        RECT 153.075 62.725 157.710 62.735 ;
        POLYGON 157.710 62.780 158.020 62.725 157.710 62.725 ;
        POLYGON 164.315 62.780 164.400 62.780 164.400 62.725 ;
        RECT 164.400 62.725 169.875 62.780 ;
        RECT 153.075 62.700 158.025 62.725 ;
        POLYGON 158.025 62.725 158.170 62.700 158.025 62.700 ;
        POLYGON 164.400 62.725 164.435 62.725 164.435 62.705 ;
        RECT 164.435 62.705 169.875 62.725 ;
        POLYGON 164.435 62.705 164.440 62.705 164.440 62.700 ;
        RECT 164.440 62.700 169.875 62.705 ;
        POLYGON 152.900 62.700 152.900 62.690 152.855 62.690 ;
        RECT 152.900 62.690 158.170 62.700 ;
        POLYGON 152.855 62.690 152.855 62.645 152.645 62.645 ;
        RECT 152.855 62.685 158.170 62.690 ;
        POLYGON 158.170 62.700 158.235 62.685 158.170 62.685 ;
        POLYGON 164.440 62.700 164.465 62.700 164.465 62.685 ;
        RECT 164.465 62.685 169.875 62.700 ;
        RECT 152.855 62.645 158.235 62.685 ;
        POLYGON 158.235 62.685 158.430 62.645 158.235 62.645 ;
        POLYGON 164.465 62.685 164.520 62.685 164.520 62.650 ;
        RECT 164.520 62.650 169.875 62.685 ;
        POLYGON 164.520 62.650 164.525 62.650 164.525 62.645 ;
        RECT 164.525 62.645 169.875 62.650 ;
        POLYGON 152.640 62.645 152.640 62.610 152.495 62.610 ;
        RECT 152.640 62.610 158.435 62.645 ;
        RECT 117.675 62.570 147.020 62.610 ;
        POLYGON 117.645 62.555 117.645 61.950 117.600 61.950 ;
        RECT 117.645 62.460 147.020 62.570 ;
        POLYGON 147.020 62.610 147.230 62.610 147.020 62.460 ;
        POLYGON 152.495 62.610 152.495 62.590 152.415 62.590 ;
        RECT 152.495 62.590 158.435 62.610 ;
        POLYGON 158.435 62.645 158.690 62.590 158.435 62.590 ;
        POLYGON 164.525 62.645 164.610 62.645 164.610 62.590 ;
        RECT 164.610 62.590 169.875 62.645 ;
        POLYGON 152.415 62.590 152.415 62.560 152.290 62.560 ;
        RECT 152.415 62.575 158.690 62.590 ;
        POLYGON 158.690 62.590 158.755 62.575 158.690 62.575 ;
        POLYGON 164.610 62.590 164.635 62.590 164.635 62.575 ;
        RECT 164.635 62.575 169.875 62.590 ;
        RECT 152.415 62.560 158.755 62.575 ;
        POLYGON 152.290 62.560 152.290 62.545 152.240 62.545 ;
        RECT 152.290 62.545 158.755 62.560 ;
        POLYGON 152.235 62.545 152.235 62.470 151.970 62.470 ;
        RECT 152.235 62.490 158.755 62.545 ;
        POLYGON 158.755 62.575 159.095 62.490 158.755 62.490 ;
        POLYGON 164.635 62.575 164.770 62.575 164.770 62.490 ;
        RECT 164.770 62.490 169.875 62.575 ;
        RECT 152.235 62.475 159.095 62.490 ;
        POLYGON 159.095 62.490 159.145 62.475 159.095 62.475 ;
        POLYGON 164.770 62.490 164.795 62.490 164.795 62.475 ;
        RECT 164.795 62.475 169.875 62.490 ;
        RECT 152.235 62.470 159.145 62.475 ;
        POLYGON 151.965 62.470 151.965 62.465 151.935 62.465 ;
        RECT 151.965 62.465 159.145 62.470 ;
        POLYGON 151.935 62.465 151.935 62.460 151.920 62.460 ;
        RECT 151.935 62.460 159.145 62.465 ;
        POLYGON 159.145 62.475 159.200 62.460 159.145 62.460 ;
        POLYGON 164.795 62.475 164.815 62.475 164.815 62.460 ;
        RECT 164.815 62.460 169.875 62.475 ;
        RECT 117.645 62.360 146.865 62.460 ;
        POLYGON 146.865 62.460 147.020 62.460 146.865 62.360 ;
        POLYGON 151.920 62.460 151.920 62.400 151.735 62.400 ;
        RECT 151.920 62.400 159.200 62.460 ;
        POLYGON 151.735 62.400 151.735 62.360 151.610 62.360 ;
        RECT 151.735 62.380 159.200 62.400 ;
        POLYGON 159.200 62.460 159.470 62.380 159.200 62.380 ;
        POLYGON 164.815 62.460 164.830 62.460 164.830 62.450 ;
        RECT 164.830 62.450 169.875 62.460 ;
        POLYGON 164.830 62.450 164.925 62.450 164.925 62.380 ;
        RECT 164.925 62.435 169.875 62.450 ;
        POLYGON 169.875 63.030 170.455 62.435 169.875 62.435 ;
        POLYGON 177.945 63.030 178.365 63.030 178.365 62.435 ;
        RECT 178.365 62.775 192.580 63.030 ;
        POLYGON 192.580 63.655 193.060 62.775 192.580 62.775 ;
        POLYGON 206.515 63.640 206.515 63.005 206.440 63.005 ;
        RECT 206.515 63.145 223.855 63.655 ;
        POLYGON 223.855 63.685 224.065 63.685 223.855 63.145 ;
        POLYGON 232.720 63.685 232.720 63.145 232.360 63.145 ;
        RECT 232.720 63.680 238.710 63.685 ;
        POLYGON 238.710 63.685 238.715 63.685 238.710 63.680 ;
        POLYGON 244.125 63.685 244.125 63.680 244.115 63.680 ;
        RECT 244.125 63.680 257.670 63.685 ;
        RECT 232.720 63.585 238.605 63.680 ;
        POLYGON 238.605 63.680 238.705 63.680 238.605 63.585 ;
        POLYGON 244.115 63.680 244.115 63.605 243.960 63.605 ;
        RECT 244.115 63.605 257.670 63.680 ;
        POLYGON 243.960 63.605 243.960 63.585 243.925 63.585 ;
        RECT 243.960 63.600 257.670 63.605 ;
        POLYGON 257.670 63.685 257.850 63.600 257.670 63.600 ;
        POLYGON 264.160 63.685 264.255 63.685 264.255 63.600 ;
        RECT 264.255 63.610 272.460 63.685 ;
        POLYGON 272.460 63.685 272.525 63.610 272.460 63.610 ;
        RECT 287.335 63.655 303.120 63.735 ;
        POLYGON 287.335 63.655 287.340 63.655 287.340 63.610 ;
        RECT 287.340 63.610 303.120 63.655 ;
        RECT 264.255 63.600 272.525 63.610 ;
        RECT 243.960 63.585 257.850 63.600 ;
        RECT 232.720 63.360 238.370 63.585 ;
        POLYGON 238.370 63.585 238.605 63.585 238.370 63.360 ;
        POLYGON 243.925 63.585 243.925 63.540 243.845 63.540 ;
        RECT 243.925 63.565 257.850 63.585 ;
        POLYGON 257.850 63.600 257.920 63.565 257.850 63.565 ;
        POLYGON 264.255 63.600 264.290 63.600 264.290 63.565 ;
        RECT 264.290 63.565 272.525 63.600 ;
        RECT 243.925 63.540 257.920 63.565 ;
        POLYGON 243.845 63.540 243.845 63.505 243.780 63.505 ;
        RECT 243.845 63.505 257.920 63.540 ;
        POLYGON 243.780 63.505 243.780 63.360 243.520 63.360 ;
        RECT 243.780 63.455 257.920 63.505 ;
        POLYGON 257.920 63.565 258.135 63.455 257.920 63.455 ;
        POLYGON 264.290 63.565 264.355 63.565 264.355 63.510 ;
        RECT 264.355 63.510 272.525 63.565 ;
        POLYGON 264.355 63.510 264.410 63.510 264.410 63.455 ;
        RECT 264.410 63.455 272.525 63.510 ;
        RECT 243.780 63.370 258.135 63.455 ;
        POLYGON 258.135 63.455 258.290 63.370 258.135 63.370 ;
        POLYGON 264.410 63.455 264.420 63.455 264.420 63.450 ;
        RECT 264.420 63.450 272.525 63.455 ;
        POLYGON 264.420 63.450 264.455 63.450 264.455 63.420 ;
        RECT 264.455 63.420 272.525 63.450 ;
        POLYGON 264.455 63.420 264.505 63.420 264.505 63.370 ;
        RECT 264.505 63.370 272.525 63.420 ;
        RECT 243.780 63.360 258.295 63.370 ;
        RECT 232.720 63.310 238.320 63.360 ;
        POLYGON 238.320 63.360 238.370 63.360 238.320 63.310 ;
        POLYGON 243.520 63.360 243.520 63.325 243.455 63.325 ;
        RECT 243.520 63.325 258.295 63.360 ;
        POLYGON 243.455 63.325 243.455 63.310 243.430 63.310 ;
        RECT 243.455 63.310 258.295 63.325 ;
        RECT 232.720 63.145 238.135 63.310 ;
        RECT 206.515 63.005 223.720 63.145 ;
        POLYGON 206.440 63.005 206.440 62.800 206.425 62.800 ;
        RECT 206.440 62.800 223.720 63.005 ;
        POLYGON 223.720 63.145 223.855 63.145 223.720 62.800 ;
        POLYGON 232.360 63.145 232.360 62.955 232.240 62.955 ;
        RECT 232.360 63.115 238.135 63.145 ;
        POLYGON 238.135 63.310 238.320 63.310 238.135 63.115 ;
        POLYGON 243.430 63.310 243.430 63.180 243.190 63.180 ;
        RECT 243.430 63.180 258.295 63.310 ;
        POLYGON 243.190 63.180 243.190 63.115 243.085 63.115 ;
        RECT 243.190 63.165 258.295 63.180 ;
        POLYGON 258.295 63.370 258.660 63.165 258.295 63.165 ;
        POLYGON 264.505 63.370 264.690 63.370 264.690 63.205 ;
        RECT 264.690 63.205 272.525 63.370 ;
        POLYGON 264.690 63.205 264.730 63.205 264.730 63.165 ;
        RECT 264.730 63.165 272.525 63.205 ;
        RECT 243.190 63.115 258.660 63.165 ;
        POLYGON 258.660 63.165 258.750 63.115 258.660 63.115 ;
        POLYGON 264.730 63.165 264.755 63.165 264.755 63.140 ;
        RECT 264.755 63.140 272.525 63.165 ;
        POLYGON 264.755 63.140 264.775 63.140 264.775 63.115 ;
        RECT 264.775 63.115 272.525 63.140 ;
        RECT 232.360 62.955 237.835 63.115 ;
        POLYGON 232.240 62.955 232.240 62.800 232.145 62.800 ;
        RECT 232.240 62.800 237.835 62.955 ;
        POLYGON 237.835 63.115 238.135 63.115 237.835 62.805 ;
        POLYGON 243.085 63.115 243.085 63.035 242.960 63.035 ;
        RECT 243.085 63.035 258.750 63.115 ;
        POLYGON 242.960 63.035 242.960 62.880 242.720 62.880 ;
        RECT 242.960 63.025 258.750 63.035 ;
        POLYGON 258.750 63.115 258.905 63.025 258.750 63.025 ;
        POLYGON 264.775 63.115 264.865 63.115 264.865 63.025 ;
        RECT 264.865 63.045 272.525 63.115 ;
        POLYGON 272.525 63.610 272.965 63.045 272.525 63.045 ;
        POLYGON 287.340 63.610 287.400 63.610 287.400 63.070 ;
        RECT 287.400 63.045 303.120 63.610 ;
        RECT 264.865 63.025 272.965 63.045 ;
        RECT 242.960 62.970 258.905 63.025 ;
        POLYGON 258.905 63.025 259.000 62.970 258.905 62.970 ;
        POLYGON 264.865 63.025 264.915 63.025 264.915 62.970 ;
        RECT 264.915 62.970 272.965 63.025 ;
        RECT 242.960 62.955 259.000 62.970 ;
        RECT 242.960 62.925 249.790 62.955 ;
        POLYGON 249.790 62.955 250.375 62.955 249.790 62.925 ;
        POLYGON 250.620 62.955 251.075 62.955 251.075 62.945 ;
        RECT 251.075 62.945 259.000 62.955 ;
        POLYGON 251.265 62.945 251.330 62.945 251.330 62.940 ;
        RECT 251.330 62.940 259.000 62.945 ;
        POLYGON 251.345 62.940 251.440 62.940 251.440 62.935 ;
        RECT 251.440 62.935 259.000 62.940 ;
        POLYGON 251.455 62.935 251.475 62.935 251.475 62.930 ;
        RECT 251.475 62.930 259.000 62.935 ;
        POLYGON 251.505 62.930 251.590 62.930 251.590 62.925 ;
        RECT 251.590 62.925 259.000 62.930 ;
        RECT 242.960 62.920 249.665 62.925 ;
        POLYGON 249.665 62.925 249.760 62.925 249.665 62.920 ;
        POLYGON 251.590 62.925 251.680 62.925 251.680 62.920 ;
        RECT 251.680 62.920 259.000 62.925 ;
        RECT 242.960 62.890 249.370 62.920 ;
        POLYGON 249.370 62.920 249.620 62.920 249.370 62.890 ;
        POLYGON 251.680 62.920 251.850 62.920 251.850 62.900 ;
        RECT 251.850 62.900 259.000 62.920 ;
        POLYGON 251.855 62.900 251.975 62.900 251.975 62.890 ;
        RECT 251.975 62.890 259.000 62.900 ;
        RECT 242.960 62.880 248.970 62.890 ;
        POLYGON 242.715 62.880 242.715 62.805 242.595 62.805 ;
        RECT 242.715 62.850 248.970 62.880 ;
        POLYGON 248.970 62.890 249.370 62.890 248.970 62.850 ;
        POLYGON 251.975 62.890 252.040 62.890 252.040 62.885 ;
        RECT 252.040 62.885 259.000 62.890 ;
        POLYGON 252.040 62.885 252.090 62.885 252.090 62.880 ;
        RECT 252.090 62.880 259.000 62.885 ;
        POLYGON 252.090 62.880 252.150 62.880 252.150 62.870 ;
        RECT 252.150 62.870 259.000 62.880 ;
        POLYGON 252.155 62.870 252.330 62.870 252.330 62.850 ;
        RECT 252.330 62.850 259.000 62.870 ;
        RECT 242.715 62.840 248.910 62.850 ;
        POLYGON 248.910 62.850 248.965 62.850 248.910 62.840 ;
        POLYGON 252.340 62.850 252.345 62.850 252.345 62.845 ;
        RECT 252.345 62.845 259.000 62.850 ;
        POLYGON 252.350 62.845 252.390 62.845 252.390 62.840 ;
        RECT 252.390 62.840 259.000 62.845 ;
        RECT 242.715 62.830 248.805 62.840 ;
        POLYGON 248.805 62.840 248.905 62.840 248.805 62.830 ;
        POLYGON 252.390 62.840 252.435 62.840 252.435 62.835 ;
        RECT 252.435 62.835 259.000 62.840 ;
        POLYGON 259.000 62.970 259.210 62.835 259.000 62.835 ;
        POLYGON 264.915 62.970 265.025 62.970 265.025 62.860 ;
        RECT 265.025 62.860 272.965 62.970 ;
        POLYGON 265.025 62.860 265.045 62.860 265.045 62.835 ;
        RECT 265.045 62.835 272.965 62.860 ;
        POLYGON 272.965 63.045 273.120 62.835 272.965 62.835 ;
        POLYGON 287.400 63.045 287.425 63.045 287.425 62.845 ;
        RECT 287.425 62.835 303.120 63.045 ;
        POLYGON 252.435 62.835 252.470 62.835 252.470 62.830 ;
        RECT 252.470 62.830 259.210 62.835 ;
        RECT 242.715 62.805 248.660 62.830 ;
        POLYGON 248.660 62.830 248.805 62.830 248.660 62.805 ;
        POLYGON 252.470 62.830 252.505 62.830 252.505 62.825 ;
        RECT 252.505 62.825 259.210 62.830 ;
        POLYGON 252.505 62.825 252.630 62.825 252.630 62.805 ;
        RECT 252.630 62.805 259.210 62.825 ;
        POLYGON 242.595 62.805 242.595 62.800 242.590 62.800 ;
        RECT 242.595 62.800 248.630 62.805 ;
        POLYGON 248.630 62.805 248.660 62.805 248.630 62.800 ;
        POLYGON 252.635 62.805 252.665 62.805 252.665 62.800 ;
        RECT 252.665 62.800 259.210 62.805 ;
        POLYGON 259.210 62.835 259.260 62.800 259.210 62.800 ;
        POLYGON 265.045 62.835 265.080 62.835 265.080 62.800 ;
        RECT 265.080 62.800 273.120 62.835 ;
        POLYGON 273.120 62.835 273.145 62.800 273.120 62.800 ;
        POLYGON 287.425 62.835 287.430 62.835 287.430 62.800 ;
        RECT 178.365 62.770 193.060 62.775 ;
        POLYGON 193.060 62.775 193.065 62.770 193.060 62.770 ;
        RECT 178.365 62.435 193.065 62.770 ;
        RECT 164.925 62.380 170.455 62.435 ;
        RECT 151.735 62.360 159.470 62.380 ;
        RECT 117.645 62.345 146.845 62.360 ;
        POLYGON 146.845 62.360 146.865 62.360 146.845 62.345 ;
        POLYGON 151.610 62.360 151.610 62.345 151.560 62.345 ;
        RECT 151.610 62.345 159.470 62.360 ;
        RECT 117.645 62.100 146.535 62.345 ;
        POLYGON 146.535 62.345 146.845 62.345 146.535 62.100 ;
        POLYGON 151.560 62.345 151.560 62.315 151.465 62.315 ;
        RECT 151.560 62.315 159.470 62.345 ;
        POLYGON 159.470 62.380 159.700 62.315 159.470 62.315 ;
        POLYGON 164.925 62.380 165.015 62.380 165.015 62.315 ;
        RECT 165.015 62.315 170.455 62.380 ;
        POLYGON 151.465 62.315 151.465 62.300 151.415 62.300 ;
        RECT 151.465 62.300 159.700 62.315 ;
        POLYGON 151.410 62.300 151.410 62.265 151.320 62.265 ;
        RECT 151.410 62.265 159.700 62.300 ;
        POLYGON 159.700 62.315 159.845 62.265 159.700 62.265 ;
        POLYGON 165.015 62.315 165.045 62.315 165.045 62.295 ;
        RECT 165.045 62.300 170.455 62.315 ;
        POLYGON 170.455 62.435 170.575 62.300 170.455 62.300 ;
        POLYGON 178.365 62.435 178.460 62.435 178.460 62.300 ;
        RECT 178.460 62.300 193.065 62.435 ;
        RECT 165.045 62.295 170.575 62.300 ;
        POLYGON 165.045 62.295 165.080 62.295 165.080 62.265 ;
        RECT 165.080 62.265 170.575 62.295 ;
        POLYGON 151.320 62.265 151.320 62.215 151.180 62.215 ;
        RECT 151.320 62.230 159.845 62.265 ;
        POLYGON 159.845 62.265 159.950 62.230 159.845 62.230 ;
        POLYGON 165.080 62.265 165.090 62.265 165.090 62.260 ;
        RECT 165.090 62.260 170.575 62.265 ;
        POLYGON 165.090 62.260 165.125 62.260 165.125 62.230 ;
        RECT 165.125 62.230 170.575 62.260 ;
        RECT 151.320 62.215 159.950 62.230 ;
        POLYGON 151.180 62.215 151.180 62.150 150.995 62.150 ;
        RECT 151.180 62.160 159.950 62.215 ;
        POLYGON 159.950 62.230 160.155 62.160 159.950 62.160 ;
        POLYGON 165.125 62.230 165.140 62.230 165.140 62.220 ;
        RECT 165.140 62.220 170.575 62.230 ;
        POLYGON 165.140 62.220 165.220 62.220 165.220 62.160 ;
        RECT 165.220 62.160 170.575 62.220 ;
        RECT 151.180 62.150 160.160 62.160 ;
        POLYGON 160.160 62.160 160.185 62.150 160.160 62.150 ;
        POLYGON 165.220 62.160 165.235 62.160 165.235 62.150 ;
        RECT 165.235 62.150 170.575 62.160 ;
        POLYGON 150.995 62.150 150.995 62.100 150.870 62.100 ;
        RECT 150.995 62.100 160.185 62.150 ;
        RECT 117.645 62.085 146.515 62.100 ;
        POLYGON 146.515 62.100 146.535 62.100 146.515 62.085 ;
        POLYGON 150.870 62.100 150.870 62.085 150.835 62.085 ;
        RECT 150.870 62.085 160.185 62.100 ;
        RECT 117.645 61.950 146.270 62.085 ;
        RECT 50.380 60.450 111.225 61.950 ;
        POLYGON 111.225 61.950 111.320 61.950 111.225 60.450 ;
        POLYGON 117.600 61.935 117.600 61.520 117.570 61.520 ;
        RECT 117.600 61.900 146.270 61.950 ;
        POLYGON 146.270 62.085 146.515 62.085 146.270 61.900 ;
        POLYGON 150.835 62.085 150.835 62.030 150.695 62.030 ;
        RECT 150.835 62.030 160.185 62.085 ;
        POLYGON 150.695 62.030 150.695 62.005 150.635 62.005 ;
        RECT 150.695 62.020 160.185 62.030 ;
        POLYGON 160.185 62.150 160.520 62.020 160.185 62.020 ;
        POLYGON 165.235 62.150 165.415 62.150 165.415 62.020 ;
        RECT 165.415 62.020 170.575 62.150 ;
        RECT 150.695 62.005 160.520 62.020 ;
        POLYGON 150.635 62.005 150.635 61.990 150.600 61.990 ;
        RECT 150.635 61.990 160.520 62.005 ;
        POLYGON 150.600 61.990 150.600 61.965 150.540 61.965 ;
        RECT 150.600 61.965 160.520 61.990 ;
        POLYGON 160.520 62.020 160.665 61.965 160.520 61.965 ;
        POLYGON 165.415 62.020 165.470 62.020 165.470 61.980 ;
        RECT 165.470 61.980 170.575 62.020 ;
        RECT 165.475 61.975 170.575 61.980 ;
        POLYGON 165.475 61.975 165.485 61.975 165.485 61.965 ;
        RECT 165.485 61.965 170.575 61.975 ;
        POLYGON 150.540 61.965 150.540 61.900 150.395 61.900 ;
        RECT 150.540 61.910 160.665 61.965 ;
        POLYGON 160.665 61.965 160.795 61.910 160.665 61.910 ;
        POLYGON 165.485 61.965 165.560 61.965 165.560 61.910 ;
        RECT 165.560 61.910 170.575 61.965 ;
        RECT 150.540 61.900 160.795 61.910 ;
        RECT 117.600 61.825 146.180 61.900 ;
        POLYGON 146.180 61.900 146.270 61.900 146.180 61.825 ;
        POLYGON 150.395 61.900 150.395 61.825 150.230 61.825 ;
        RECT 150.395 61.895 160.795 61.900 ;
        POLYGON 160.795 61.910 160.830 61.895 160.795 61.895 ;
        POLYGON 165.560 61.910 165.580 61.910 165.580 61.895 ;
        RECT 165.580 61.895 170.575 61.910 ;
        RECT 150.395 61.825 160.830 61.895 ;
        RECT 117.600 61.820 146.170 61.825 ;
        POLYGON 146.170 61.825 146.180 61.825 146.170 61.820 ;
        POLYGON 150.230 61.825 150.230 61.820 150.215 61.820 ;
        RECT 150.230 61.820 160.830 61.825 ;
        RECT 117.600 61.725 146.060 61.820 ;
        POLYGON 146.060 61.820 146.170 61.820 146.060 61.725 ;
        POLYGON 150.215 61.820 150.215 61.765 150.095 61.765 ;
        RECT 150.215 61.770 160.830 61.820 ;
        POLYGON 160.830 61.895 161.130 61.770 160.830 61.770 ;
        POLYGON 165.580 61.895 165.730 61.895 165.730 61.770 ;
        RECT 165.730 61.770 170.575 61.895 ;
        RECT 150.215 61.765 161.130 61.770 ;
        POLYGON 150.090 61.765 150.090 61.725 150.010 61.725 ;
        RECT 150.090 61.745 161.130 61.765 ;
        POLYGON 161.130 61.770 161.175 61.745 161.130 61.745 ;
        POLYGON 165.730 61.770 165.765 61.770 165.765 61.745 ;
        RECT 165.765 61.745 170.575 61.770 ;
        RECT 150.090 61.725 161.175 61.745 ;
        RECT 117.600 61.545 145.855 61.725 ;
        POLYGON 145.855 61.725 146.060 61.725 145.855 61.545 ;
        POLYGON 150.010 61.725 150.010 61.625 149.805 61.625 ;
        RECT 150.010 61.625 161.175 61.725 ;
        POLYGON 149.805 61.625 149.805 61.595 149.750 61.595 ;
        RECT 149.805 61.600 161.175 61.625 ;
        POLYGON 161.175 61.745 161.485 61.600 161.175 61.600 ;
        POLYGON 165.765 61.745 165.790 61.745 165.790 61.725 ;
        RECT 165.790 61.725 170.575 61.745 ;
        POLYGON 165.790 61.725 165.845 61.725 165.845 61.680 ;
        RECT 165.845 61.680 170.575 61.725 ;
        POLYGON 165.845 61.680 165.940 61.680 165.940 61.600 ;
        RECT 165.940 61.600 170.575 61.680 ;
        RECT 149.805 61.595 161.485 61.600 ;
        POLYGON 149.750 61.595 149.750 61.545 149.650 61.545 ;
        RECT 149.750 61.555 161.485 61.595 ;
        POLYGON 161.485 61.600 161.585 61.555 161.485 61.555 ;
        POLYGON 165.940 61.600 165.995 61.600 165.995 61.555 ;
        RECT 165.995 61.555 170.575 61.600 ;
        RECT 149.750 61.545 161.585 61.555 ;
        RECT 117.600 61.520 145.595 61.545 ;
        POLYGON 117.570 61.510 117.570 60.525 117.500 60.525 ;
        RECT 117.570 61.315 145.595 61.520 ;
        POLYGON 145.595 61.545 145.855 61.545 145.595 61.315 ;
        POLYGON 149.650 61.545 149.650 61.500 149.565 61.500 ;
        RECT 149.650 61.530 161.585 61.545 ;
        POLYGON 161.585 61.555 161.635 61.530 161.585 61.530 ;
        POLYGON 165.995 61.555 166.025 61.555 166.025 61.530 ;
        RECT 166.025 61.530 170.575 61.555 ;
        RECT 149.650 61.500 161.635 61.530 ;
        POLYGON 149.565 61.500 149.565 61.315 149.230 61.315 ;
        RECT 149.565 61.440 161.635 61.500 ;
        POLYGON 161.635 61.530 161.805 61.440 161.635 61.440 ;
        POLYGON 166.025 61.530 166.050 61.530 166.050 61.510 ;
        RECT 166.050 61.515 170.575 61.530 ;
        POLYGON 170.575 62.300 171.260 61.515 170.575 61.515 ;
        POLYGON 178.460 62.300 178.660 62.300 178.660 62.020 ;
        RECT 178.660 62.020 193.065 62.300 ;
        POLYGON 178.660 62.020 178.975 62.020 178.975 61.515 ;
        RECT 178.975 61.975 193.065 62.020 ;
        POLYGON 193.065 62.770 193.465 61.975 193.065 61.975 ;
        RECT 178.975 61.515 193.465 61.975 ;
        POLYGON 206.425 62.770 206.425 62.005 206.375 62.005 ;
        RECT 206.425 62.545 223.620 62.800 ;
        POLYGON 223.620 62.800 223.720 62.800 223.620 62.545 ;
        POLYGON 232.145 62.795 232.145 62.550 231.995 62.550 ;
        RECT 232.145 62.695 237.730 62.800 ;
        POLYGON 237.730 62.800 237.835 62.800 237.730 62.695 ;
        POLYGON 242.590 62.800 242.590 62.705 242.440 62.705 ;
        RECT 242.590 62.755 248.370 62.800 ;
        POLYGON 248.370 62.800 248.630 62.800 248.370 62.755 ;
        POLYGON 252.665 62.800 252.700 62.800 252.700 62.795 ;
        RECT 252.700 62.795 259.260 62.800 ;
        POLYGON 252.705 62.795 252.905 62.795 252.905 62.765 ;
        RECT 252.905 62.765 259.260 62.795 ;
        POLYGON 252.905 62.765 252.915 62.765 252.915 62.760 ;
        RECT 252.915 62.760 259.260 62.765 ;
        POLYGON 252.915 62.760 252.940 62.760 252.940 62.755 ;
        RECT 252.940 62.755 259.260 62.760 ;
        RECT 242.590 62.745 248.320 62.755 ;
        POLYGON 248.320 62.755 248.370 62.755 248.320 62.745 ;
        POLYGON 252.940 62.755 252.970 62.755 252.970 62.750 ;
        RECT 252.970 62.750 259.260 62.755 ;
        POLYGON 252.970 62.750 252.995 62.750 252.995 62.745 ;
        RECT 252.995 62.745 259.260 62.750 ;
        RECT 242.590 62.710 248.100 62.745 ;
        POLYGON 248.100 62.745 248.315 62.745 248.100 62.710 ;
        POLYGON 252.995 62.745 253.165 62.745 253.165 62.715 ;
        RECT 253.165 62.715 259.260 62.745 ;
        POLYGON 253.165 62.715 253.185 62.715 253.185 62.710 ;
        RECT 253.185 62.710 259.260 62.715 ;
        RECT 242.590 62.705 248.055 62.710 ;
        POLYGON 242.440 62.705 242.440 62.695 242.425 62.695 ;
        RECT 242.440 62.700 248.055 62.705 ;
        POLYGON 248.055 62.710 248.100 62.710 248.055 62.700 ;
        POLYGON 253.195 62.710 253.230 62.710 253.230 62.705 ;
        RECT 253.230 62.705 259.260 62.710 ;
        POLYGON 253.230 62.705 253.250 62.705 253.250 62.700 ;
        RECT 253.250 62.700 259.260 62.705 ;
        RECT 242.440 62.695 247.995 62.700 ;
        RECT 232.145 62.670 237.715 62.695 ;
        POLYGON 237.715 62.695 237.730 62.695 237.715 62.670 ;
        POLYGON 242.425 62.695 242.425 62.670 242.390 62.670 ;
        RECT 242.425 62.690 247.995 62.695 ;
        POLYGON 247.995 62.700 248.055 62.700 247.995 62.690 ;
        POLYGON 253.250 62.700 253.300 62.700 253.300 62.690 ;
        RECT 253.300 62.690 259.260 62.700 ;
        RECT 242.425 62.670 247.840 62.690 ;
        RECT 232.145 62.620 237.670 62.670 ;
        POLYGON 237.670 62.670 237.715 62.670 237.670 62.620 ;
        POLYGON 242.390 62.670 242.390 62.660 242.380 62.660 ;
        RECT 242.390 62.660 247.840 62.670 ;
        POLYGON 242.380 62.660 242.380 62.620 242.325 62.620 ;
        RECT 242.380 62.655 247.840 62.660 ;
        POLYGON 247.840 62.690 247.995 62.690 247.840 62.655 ;
        POLYGON 253.300 62.690 253.325 62.690 253.325 62.685 ;
        RECT 253.325 62.685 259.260 62.690 ;
        POLYGON 253.325 62.685 253.415 62.685 253.415 62.665 ;
        RECT 253.415 62.665 259.260 62.685 ;
        POLYGON 253.415 62.665 253.455 62.665 253.455 62.655 ;
        RECT 253.455 62.655 259.260 62.665 ;
        RECT 242.380 62.620 247.590 62.655 ;
        RECT 232.145 62.550 237.335 62.620 ;
        RECT 206.425 62.265 223.530 62.545 ;
        POLYGON 223.530 62.545 223.620 62.545 223.530 62.265 ;
        POLYGON 231.995 62.545 231.995 62.390 231.900 62.390 ;
        RECT 231.995 62.390 237.335 62.550 ;
        POLYGON 231.900 62.390 231.900 62.265 231.830 62.265 ;
        RECT 231.900 62.265 237.335 62.390 ;
        RECT 206.425 62.005 223.450 62.265 ;
        POLYGON 223.450 62.265 223.530 62.265 223.450 62.015 ;
        POLYGON 231.830 62.265 231.830 62.020 231.695 62.020 ;
        RECT 231.830 62.235 237.335 62.265 ;
        POLYGON 237.335 62.620 237.670 62.620 237.335 62.235 ;
        POLYGON 242.325 62.620 242.325 62.465 242.110 62.465 ;
        RECT 242.325 62.595 247.590 62.620 ;
        POLYGON 247.590 62.655 247.840 62.655 247.590 62.595 ;
        POLYGON 253.455 62.655 253.500 62.655 253.500 62.645 ;
        RECT 253.500 62.645 259.260 62.655 ;
        POLYGON 253.505 62.645 253.665 62.645 253.665 62.610 ;
        RECT 253.665 62.610 259.260 62.645 ;
        POLYGON 253.670 62.610 253.715 62.610 253.715 62.595 ;
        RECT 253.715 62.595 259.260 62.610 ;
        RECT 242.325 62.570 247.485 62.595 ;
        POLYGON 247.485 62.595 247.590 62.595 247.485 62.570 ;
        POLYGON 253.715 62.595 253.815 62.595 253.815 62.570 ;
        RECT 253.815 62.570 259.260 62.595 ;
        RECT 242.325 62.535 247.340 62.570 ;
        POLYGON 247.340 62.570 247.485 62.570 247.340 62.535 ;
        POLYGON 253.815 62.570 253.920 62.570 253.920 62.545 ;
        RECT 253.920 62.550 259.260 62.570 ;
        POLYGON 259.260 62.800 259.655 62.550 259.260 62.550 ;
        POLYGON 265.080 62.800 265.280 62.800 265.280 62.600 ;
        RECT 265.280 62.600 273.145 62.800 ;
        POLYGON 265.280 62.600 265.325 62.600 265.325 62.550 ;
        RECT 265.325 62.550 273.145 62.600 ;
        RECT 253.920 62.545 259.655 62.550 ;
        POLYGON 253.925 62.545 253.960 62.545 253.960 62.535 ;
        RECT 253.960 62.535 259.655 62.545 ;
        RECT 242.325 62.505 247.210 62.535 ;
        POLYGON 247.210 62.535 247.335 62.535 247.210 62.505 ;
        POLYGON 253.960 62.535 254.040 62.535 254.040 62.515 ;
        RECT 254.040 62.515 259.655 62.535 ;
        POLYGON 254.045 62.515 254.075 62.515 254.075 62.505 ;
        RECT 254.075 62.505 259.655 62.515 ;
        RECT 242.325 62.500 247.200 62.505 ;
        POLYGON 247.200 62.505 247.210 62.505 247.200 62.500 ;
        POLYGON 254.075 62.505 254.090 62.505 254.090 62.500 ;
        RECT 254.090 62.500 259.655 62.505 ;
        RECT 242.325 62.480 247.130 62.500 ;
        POLYGON 247.130 62.500 247.200 62.500 247.130 62.480 ;
        POLYGON 254.090 62.500 254.145 62.500 254.145 62.485 ;
        RECT 254.145 62.485 259.655 62.500 ;
        POLYGON 254.145 62.485 254.165 62.485 254.165 62.480 ;
        RECT 254.165 62.480 259.655 62.485 ;
        RECT 242.325 62.465 247.085 62.480 ;
        POLYGON 247.085 62.480 247.130 62.480 247.085 62.465 ;
        POLYGON 254.165 62.480 254.185 62.480 254.185 62.475 ;
        RECT 254.185 62.475 259.655 62.480 ;
        POLYGON 254.185 62.475 254.215 62.475 254.215 62.465 ;
        RECT 254.215 62.465 259.655 62.475 ;
        POLYGON 242.110 62.465 242.110 62.235 241.785 62.235 ;
        RECT 242.110 62.385 246.820 62.465 ;
        POLYGON 246.820 62.465 247.085 62.465 246.820 62.385 ;
        POLYGON 254.215 62.465 254.495 62.465 254.495 62.385 ;
        RECT 254.495 62.435 259.655 62.465 ;
        POLYGON 259.655 62.550 259.820 62.435 259.655 62.435 ;
        POLYGON 265.325 62.550 265.440 62.550 265.440 62.435 ;
        RECT 265.440 62.500 273.145 62.550 ;
        POLYGON 273.145 62.800 273.365 62.500 273.145 62.500 ;
        RECT 287.430 62.770 303.120 62.835 ;
        POLYGON 287.430 62.770 287.455 62.770 287.455 62.535 ;
        RECT 287.455 62.500 303.120 62.770 ;
        RECT 265.440 62.435 273.365 62.500 ;
        RECT 254.495 62.385 259.820 62.435 ;
        RECT 242.110 62.380 246.805 62.385 ;
        POLYGON 246.805 62.385 246.820 62.385 246.805 62.380 ;
        POLYGON 254.495 62.385 254.515 62.385 254.515 62.380 ;
        RECT 254.515 62.380 259.820 62.385 ;
        RECT 242.110 62.290 246.505 62.380 ;
        POLYGON 246.505 62.380 246.805 62.380 246.505 62.290 ;
        POLYGON 254.515 62.380 254.550 62.380 254.550 62.370 ;
        RECT 254.550 62.370 259.820 62.380 ;
        POLYGON 254.550 62.370 254.755 62.370 254.755 62.300 ;
        RECT 254.755 62.300 259.820 62.370 ;
        POLYGON 254.755 62.300 254.785 62.300 254.785 62.290 ;
        RECT 254.785 62.290 259.820 62.300 ;
        RECT 242.110 62.265 246.420 62.290 ;
        POLYGON 246.420 62.290 246.505 62.290 246.420 62.265 ;
        POLYGON 254.785 62.290 254.865 62.290 254.865 62.265 ;
        RECT 254.865 62.275 259.820 62.290 ;
        POLYGON 259.820 62.435 260.045 62.275 259.820 62.275 ;
        POLYGON 265.440 62.435 265.495 62.435 265.495 62.380 ;
        RECT 265.495 62.380 273.365 62.435 ;
        POLYGON 265.495 62.380 265.515 62.380 265.515 62.355 ;
        RECT 265.515 62.355 273.365 62.380 ;
        POLYGON 265.515 62.355 265.585 62.355 265.585 62.275 ;
        RECT 265.585 62.275 273.365 62.355 ;
        RECT 254.865 62.265 260.045 62.275 ;
        RECT 242.110 62.250 246.380 62.265 ;
        POLYGON 246.380 62.265 246.420 62.265 246.380 62.250 ;
        POLYGON 254.865 62.265 254.885 62.265 254.885 62.260 ;
        RECT 254.885 62.260 260.045 62.265 ;
        POLYGON 254.885 62.260 254.910 62.260 254.910 62.250 ;
        RECT 254.910 62.250 260.045 62.260 ;
        RECT 242.110 62.235 246.245 62.250 ;
        RECT 231.830 62.020 237.140 62.235 ;
        POLYGON 231.695 62.015 231.695 62.010 231.690 62.010 ;
        RECT 231.695 62.010 237.140 62.020 ;
        RECT 231.690 62.005 237.140 62.010 ;
        POLYGON 237.140 62.235 237.335 62.235 237.140 62.005 ;
        POLYGON 241.785 62.235 241.785 62.180 241.710 62.180 ;
        RECT 241.785 62.200 246.245 62.235 ;
        POLYGON 246.245 62.250 246.375 62.250 246.245 62.200 ;
        POLYGON 254.910 62.250 254.955 62.250 254.955 62.235 ;
        RECT 254.955 62.235 260.045 62.250 ;
        POLYGON 254.955 62.235 255.050 62.235 255.050 62.200 ;
        RECT 255.050 62.200 260.045 62.235 ;
        POLYGON 260.045 62.275 260.145 62.200 260.045 62.200 ;
        POLYGON 265.585 62.275 265.650 62.275 265.650 62.200 ;
        RECT 265.650 62.265 273.365 62.275 ;
        POLYGON 273.365 62.500 273.525 62.265 273.365 62.265 ;
        POLYGON 287.455 62.500 287.480 62.500 287.480 62.300 ;
        RECT 287.480 62.265 303.120 62.500 ;
        RECT 265.650 62.200 273.525 62.265 ;
        RECT 241.785 62.190 246.220 62.200 ;
        POLYGON 246.220 62.200 246.245 62.200 246.220 62.190 ;
        POLYGON 255.050 62.200 255.080 62.200 255.080 62.190 ;
        RECT 255.080 62.190 260.145 62.200 ;
        RECT 241.785 62.180 246.040 62.190 ;
        POLYGON 241.710 62.175 241.710 62.150 241.680 62.150 ;
        RECT 241.710 62.150 246.040 62.180 ;
        POLYGON 241.680 62.150 241.680 62.005 241.500 62.005 ;
        RECT 241.680 62.125 246.040 62.150 ;
        POLYGON 246.040 62.190 246.220 62.190 246.040 62.125 ;
        POLYGON 255.080 62.190 255.265 62.190 255.265 62.125 ;
        RECT 255.265 62.125 260.145 62.190 ;
        RECT 241.680 62.090 245.945 62.125 ;
        POLYGON 245.945 62.125 246.040 62.125 245.945 62.090 ;
        POLYGON 255.265 62.125 255.280 62.125 255.280 62.120 ;
        RECT 255.280 62.120 260.145 62.125 ;
        POLYGON 255.280 62.120 255.355 62.120 255.355 62.090 ;
        RECT 255.355 62.090 260.145 62.120 ;
        RECT 241.680 62.005 245.735 62.090 ;
        POLYGON 245.735 62.090 245.945 62.090 245.735 62.005 ;
        POLYGON 255.355 62.090 255.420 62.090 255.420 62.065 ;
        RECT 255.420 62.065 260.145 62.090 ;
        POLYGON 255.420 62.065 255.570 62.065 255.570 62.005 ;
        RECT 255.570 62.030 260.145 62.065 ;
        POLYGON 260.145 62.200 260.385 62.030 260.145 62.030 ;
        POLYGON 265.650 62.200 265.705 62.200 265.705 62.140 ;
        RECT 265.705 62.140 273.525 62.200 ;
        POLYGON 265.705 62.140 265.730 62.140 265.730 62.110 ;
        RECT 265.730 62.110 273.525 62.140 ;
        POLYGON 265.730 62.110 265.795 62.110 265.795 62.035 ;
        RECT 265.795 62.030 273.525 62.110 ;
        RECT 255.570 62.005 260.385 62.030 ;
        POLYGON 260.385 62.030 260.415 62.005 260.385 62.005 ;
        POLYGON 265.795 62.030 265.820 62.030 265.820 62.005 ;
        RECT 265.820 62.010 273.525 62.030 ;
        POLYGON 273.525 62.265 273.695 62.010 273.525 62.010 ;
        POLYGON 287.480 62.265 287.490 62.265 287.490 62.210 ;
        RECT 287.490 62.210 303.120 62.265 ;
        RECT 265.820 62.005 273.695 62.010 ;
        POLYGON 287.490 62.210 287.515 62.210 287.515 62.005 ;
        RECT 166.050 61.510 171.260 61.515 ;
        POLYGON 166.050 61.510 166.095 61.510 166.095 61.470 ;
        RECT 166.095 61.485 171.260 61.510 ;
        POLYGON 171.260 61.515 171.285 61.485 171.260 61.485 ;
        POLYGON 178.975 61.515 178.995 61.515 178.995 61.485 ;
        RECT 178.995 61.485 193.465 61.515 ;
        RECT 166.095 61.470 171.285 61.485 ;
        POLYGON 166.095 61.470 166.130 61.470 166.130 61.440 ;
        RECT 166.130 61.440 171.285 61.470 ;
        RECT 149.565 61.325 161.805 61.440 ;
        POLYGON 161.805 61.440 162.025 61.325 161.805 61.325 ;
        POLYGON 166.130 61.440 166.190 61.440 166.190 61.390 ;
        RECT 166.190 61.430 171.285 61.440 ;
        POLYGON 171.285 61.485 171.325 61.430 171.285 61.430 ;
        POLYGON 178.995 61.485 179.025 61.485 179.025 61.435 ;
        RECT 179.025 61.430 193.465 61.485 ;
        RECT 166.190 61.390 171.325 61.430 ;
        POLYGON 166.190 61.390 166.270 61.390 166.270 61.325 ;
        RECT 166.270 61.325 171.325 61.390 ;
        RECT 149.565 61.315 162.025 61.325 ;
        RECT 117.570 61.270 145.545 61.315 ;
        POLYGON 145.545 61.315 145.595 61.315 145.545 61.270 ;
        POLYGON 149.230 61.315 149.230 61.310 149.220 61.310 ;
        RECT 149.230 61.310 162.025 61.315 ;
        POLYGON 149.220 61.310 149.220 61.270 149.155 61.270 ;
        RECT 149.220 61.270 162.025 61.310 ;
        POLYGON 162.025 61.325 162.120 61.270 162.025 61.270 ;
        POLYGON 166.270 61.325 166.310 61.325 166.310 61.295 ;
        RECT 166.310 61.295 171.325 61.325 ;
        POLYGON 166.310 61.295 166.335 61.295 166.335 61.270 ;
        RECT 166.335 61.285 171.325 61.295 ;
        POLYGON 171.325 61.430 171.435 61.285 171.325 61.285 ;
        POLYGON 179.025 61.430 179.105 61.430 179.105 61.310 ;
        RECT 179.105 61.405 193.465 61.430 ;
        POLYGON 193.465 61.970 193.750 61.405 193.465 61.405 ;
        POLYGON 206.375 61.970 206.375 61.465 206.340 61.465 ;
        RECT 206.375 61.465 223.270 62.005 ;
        POLYGON 206.340 61.450 206.340 61.405 206.335 61.405 ;
        RECT 206.340 61.445 223.270 61.465 ;
        POLYGON 223.270 62.005 223.450 62.005 223.270 61.450 ;
        POLYGON 231.690 62.005 231.690 61.810 231.580 61.810 ;
        RECT 231.690 62.000 237.135 62.005 ;
        POLYGON 237.135 62.005 237.140 62.005 237.135 62.000 ;
        POLYGON 241.500 62.005 241.500 62.000 241.495 62.000 ;
        RECT 241.500 62.000 245.670 62.005 ;
        RECT 231.690 61.860 237.025 62.000 ;
        POLYGON 237.025 62.000 237.135 62.000 237.025 61.860 ;
        POLYGON 241.495 62.000 241.495 61.860 241.320 61.860 ;
        RECT 241.495 61.980 245.670 62.000 ;
        POLYGON 245.670 62.005 245.735 62.005 245.670 61.980 ;
        POLYGON 255.570 62.005 255.630 62.005 255.630 61.980 ;
        RECT 255.630 61.980 260.415 62.005 ;
        RECT 241.495 61.975 245.660 61.980 ;
        POLYGON 245.660 61.980 245.665 61.980 245.660 61.975 ;
        POLYGON 255.630 61.980 255.645 61.980 255.645 61.975 ;
        RECT 255.645 61.975 260.415 61.980 ;
        RECT 241.495 61.945 245.580 61.975 ;
        POLYGON 245.580 61.975 245.660 61.975 245.580 61.945 ;
        POLYGON 255.645 61.975 255.720 61.975 255.720 61.945 ;
        RECT 255.720 61.945 260.415 61.975 ;
        RECT 241.495 61.935 245.560 61.945 ;
        POLYGON 245.560 61.945 245.580 61.945 245.560 61.935 ;
        POLYGON 255.720 61.945 255.740 61.945 255.740 61.935 ;
        RECT 255.740 61.935 260.415 61.945 ;
        RECT 241.495 61.860 245.385 61.935 ;
        POLYGON 245.385 61.935 245.560 61.935 245.385 61.860 ;
        POLYGON 255.740 61.935 255.750 61.935 255.750 61.930 ;
        RECT 255.750 61.930 260.415 61.935 ;
        POLYGON 255.750 61.930 255.775 61.930 255.775 61.920 ;
        RECT 255.775 61.920 260.415 61.930 ;
        POLYGON 255.775 61.920 255.815 61.920 255.815 61.905 ;
        RECT 255.815 61.905 260.415 61.920 ;
        POLYGON 255.815 61.905 255.915 61.905 255.915 61.860 ;
        RECT 255.915 61.860 260.415 61.905 ;
        RECT 231.690 61.835 237.005 61.860 ;
        POLYGON 237.005 61.860 237.025 61.860 237.005 61.835 ;
        POLYGON 241.320 61.860 241.320 61.855 241.315 61.855 ;
        RECT 241.320 61.855 245.285 61.860 ;
        POLYGON 241.315 61.855 241.315 61.835 241.290 61.835 ;
        RECT 241.315 61.835 245.285 61.855 ;
        RECT 231.690 61.810 236.875 61.835 ;
        POLYGON 231.580 61.810 231.580 61.450 231.400 61.450 ;
        RECT 231.580 61.660 236.875 61.810 ;
        POLYGON 236.875 61.835 237.005 61.835 236.875 61.660 ;
        POLYGON 241.290 61.835 241.290 61.660 241.075 61.660 ;
        RECT 241.290 61.815 245.285 61.835 ;
        POLYGON 245.285 61.860 245.385 61.860 245.285 61.815 ;
        POLYGON 255.915 61.860 256.015 61.860 256.015 61.815 ;
        RECT 256.015 61.815 260.415 61.860 ;
        RECT 241.290 61.725 245.095 61.815 ;
        POLYGON 245.095 61.815 245.285 61.815 245.095 61.725 ;
        POLYGON 256.015 61.815 256.145 61.815 256.145 61.760 ;
        RECT 256.145 61.760 260.415 61.815 ;
        POLYGON 256.145 61.760 256.200 61.760 256.200 61.735 ;
        RECT 256.200 61.735 260.415 61.760 ;
        POLYGON 256.200 61.735 256.215 61.735 256.215 61.725 ;
        RECT 256.215 61.725 260.415 61.735 ;
        RECT 241.290 61.660 244.915 61.725 ;
        RECT 231.580 61.470 236.725 61.660 ;
        POLYGON 236.725 61.660 236.875 61.660 236.725 61.470 ;
        POLYGON 241.075 61.660 241.075 61.605 241.010 61.605 ;
        RECT 241.075 61.645 244.915 61.660 ;
        POLYGON 244.915 61.725 245.095 61.725 244.915 61.645 ;
        POLYGON 256.215 61.725 256.375 61.725 256.375 61.645 ;
        RECT 256.375 61.645 260.415 61.725 ;
        RECT 241.075 61.635 244.900 61.645 ;
        POLYGON 244.900 61.645 244.915 61.645 244.900 61.635 ;
        POLYGON 256.375 61.645 256.400 61.645 256.400 61.635 ;
        RECT 256.400 61.635 260.415 61.645 ;
        RECT 241.075 61.605 244.550 61.635 ;
        POLYGON 241.010 61.605 241.010 61.470 240.865 61.470 ;
        RECT 241.010 61.470 244.550 61.605 ;
        RECT 231.580 61.450 236.710 61.470 ;
        POLYGON 236.710 61.470 236.725 61.470 236.710 61.450 ;
        POLYGON 240.865 61.470 240.865 61.450 240.845 61.450 ;
        RECT 240.865 61.460 244.550 61.470 ;
        POLYGON 244.550 61.635 244.900 61.635 244.550 61.460 ;
        POLYGON 256.400 61.635 256.535 61.635 256.535 61.570 ;
        RECT 256.535 61.570 260.415 61.635 ;
        POLYGON 256.540 61.570 256.570 61.570 256.570 61.555 ;
        RECT 256.570 61.555 260.415 61.570 ;
        POLYGON 260.415 62.005 260.970 61.555 260.415 61.555 ;
        POLYGON 265.820 62.005 265.900 62.005 265.900 61.915 ;
        RECT 265.900 61.975 273.695 62.005 ;
        POLYGON 273.695 62.005 273.720 61.975 273.695 61.975 ;
        RECT 265.900 61.915 273.720 61.975 ;
        POLYGON 265.900 61.915 265.920 61.915 265.920 61.890 ;
        RECT 265.920 61.890 273.720 61.915 ;
        POLYGON 265.920 61.890 265.950 61.890 265.950 61.855 ;
        RECT 265.950 61.855 273.720 61.890 ;
        POLYGON 265.950 61.855 266.075 61.855 266.075 61.710 ;
        RECT 266.075 61.780 273.720 61.855 ;
        POLYGON 273.720 61.975 273.840 61.780 273.720 61.780 ;
        RECT 287.515 61.970 303.120 62.210 ;
        POLYGON 287.515 61.970 287.535 61.970 287.535 61.795 ;
        RECT 287.535 61.780 303.120 61.970 ;
        RECT 266.075 61.710 273.840 61.780 ;
        POLYGON 266.075 61.710 266.095 61.710 266.095 61.690 ;
        RECT 266.095 61.690 273.840 61.710 ;
        POLYGON 266.095 61.690 266.210 61.690 266.210 61.555 ;
        RECT 266.210 61.555 273.840 61.690 ;
        POLYGON 256.570 61.555 256.715 61.555 256.715 61.475 ;
        RECT 256.715 61.490 260.970 61.555 ;
        POLYGON 260.970 61.555 261.050 61.490 260.970 61.490 ;
        POLYGON 266.210 61.555 266.230 61.555 266.230 61.535 ;
        RECT 266.230 61.535 273.840 61.555 ;
        POLYGON 266.230 61.535 266.245 61.535 266.245 61.515 ;
        RECT 266.245 61.515 273.840 61.535 ;
        POLYGON 266.245 61.515 266.255 61.515 266.255 61.505 ;
        RECT 266.255 61.505 273.840 61.515 ;
        POLYGON 266.255 61.505 266.265 61.505 266.265 61.490 ;
        RECT 266.265 61.490 273.840 61.505 ;
        RECT 256.715 61.475 261.050 61.490 ;
        POLYGON 261.050 61.490 261.070 61.475 261.050 61.475 ;
        POLYGON 266.265 61.490 266.275 61.490 266.275 61.475 ;
        RECT 266.275 61.475 273.840 61.490 ;
        POLYGON 256.720 61.475 256.745 61.475 256.745 61.460 ;
        RECT 256.745 61.460 261.070 61.475 ;
        RECT 240.865 61.450 244.535 61.460 ;
        POLYGON 244.535 61.460 244.550 61.460 244.535 61.450 ;
        POLYGON 256.745 61.460 256.765 61.460 256.765 61.450 ;
        RECT 256.765 61.450 261.070 61.460 ;
        POLYGON 261.070 61.475 261.095 61.450 261.070 61.450 ;
        POLYGON 266.275 61.475 266.295 61.475 266.295 61.450 ;
        RECT 266.295 61.450 273.840 61.475 ;
        POLYGON 273.840 61.780 274.045 61.450 273.840 61.450 ;
        POLYGON 287.535 61.780 287.575 61.780 287.575 61.450 ;
        RECT 206.340 61.405 223.235 61.445 ;
        RECT 179.105 61.310 193.750 61.405 ;
        POLYGON 179.105 61.310 179.120 61.310 179.120 61.285 ;
        RECT 179.120 61.285 193.750 61.310 ;
        RECT 166.335 61.270 171.435 61.285 ;
        RECT 117.570 61.250 145.525 61.270 ;
        POLYGON 145.525 61.270 145.545 61.270 145.525 61.250 ;
        POLYGON 149.155 61.270 149.155 61.250 149.120 61.250 ;
        RECT 149.155 61.250 162.120 61.270 ;
        RECT 117.570 61.215 145.485 61.250 ;
        POLYGON 145.485 61.250 145.525 61.250 145.485 61.215 ;
        POLYGON 149.120 61.250 149.120 61.215 149.065 61.215 ;
        RECT 149.120 61.215 162.120 61.250 ;
        RECT 117.570 60.880 145.230 61.215 ;
        POLYGON 145.230 61.215 145.485 61.215 145.230 60.960 ;
        POLYGON 149.065 61.215 149.065 61.200 149.040 61.200 ;
        RECT 149.065 61.200 162.120 61.215 ;
        POLYGON 149.030 61.200 149.030 61.075 148.830 61.075 ;
        RECT 149.030 61.175 162.120 61.200 ;
        RECT 149.030 61.170 154.915 61.175 ;
        POLYGON 154.915 61.175 155.495 61.175 154.915 61.170 ;
        POLYGON 155.495 61.175 155.855 61.175 155.855 61.170 ;
        RECT 155.855 61.170 162.120 61.175 ;
        RECT 149.030 61.160 154.410 61.170 ;
        POLYGON 154.410 61.170 154.655 61.170 154.410 61.160 ;
        POLYGON 156.335 61.170 156.365 61.170 156.365 61.165 ;
        RECT 156.365 61.165 162.120 61.170 ;
        POLYGON 156.375 61.165 156.530 61.165 156.530 61.160 ;
        RECT 156.530 61.160 162.120 61.165 ;
        RECT 149.030 61.155 154.290 61.160 ;
        POLYGON 154.290 61.160 154.400 61.160 154.290 61.155 ;
        POLYGON 156.570 61.160 156.645 61.160 156.645 61.155 ;
        RECT 156.645 61.155 162.120 61.160 ;
        RECT 149.030 61.145 153.955 61.155 ;
        POLYGON 153.955 61.155 154.280 61.155 153.955 61.145 ;
        POLYGON 156.660 61.155 156.925 61.155 156.925 61.145 ;
        RECT 156.925 61.145 162.120 61.155 ;
        RECT 149.030 61.140 153.905 61.145 ;
        POLYGON 153.905 61.145 153.955 61.145 153.905 61.140 ;
        POLYGON 157.035 61.145 157.090 61.145 157.090 61.140 ;
        RECT 157.090 61.140 162.120 61.145 ;
        RECT 149.030 61.125 153.735 61.140 ;
        POLYGON 153.735 61.140 153.900 61.140 153.735 61.125 ;
        POLYGON 157.105 61.140 157.130 61.140 157.130 61.135 ;
        RECT 157.130 61.135 162.120 61.140 ;
        POLYGON 157.140 61.135 157.180 61.135 157.180 61.130 ;
        RECT 157.180 61.130 162.120 61.135 ;
        POLYGON 157.185 61.130 157.260 61.130 157.260 61.125 ;
        RECT 157.260 61.125 162.120 61.130 ;
        RECT 149.030 61.120 153.645 61.125 ;
        POLYGON 153.645 61.125 153.725 61.125 153.645 61.120 ;
        POLYGON 157.260 61.125 157.340 61.125 157.340 61.120 ;
        RECT 157.340 61.120 162.120 61.125 ;
        RECT 149.030 61.095 153.400 61.120 ;
        POLYGON 153.400 61.120 153.645 61.120 153.400 61.095 ;
        POLYGON 157.340 61.120 157.435 61.120 157.435 61.110 ;
        RECT 157.435 61.110 162.120 61.120 ;
        POLYGON 157.440 61.110 157.580 61.110 157.580 61.095 ;
        RECT 157.580 61.095 162.120 61.110 ;
        RECT 149.030 61.090 153.360 61.095 ;
        POLYGON 153.360 61.095 153.395 61.095 153.360 61.090 ;
        POLYGON 157.580 61.095 157.630 61.095 157.630 61.090 ;
        RECT 157.630 61.090 162.120 61.095 ;
        RECT 149.030 61.075 153.180 61.090 ;
        POLYGON 148.830 61.075 148.830 61.060 148.800 61.060 ;
        RECT 148.830 61.060 153.180 61.075 ;
        POLYGON 153.180 61.090 153.360 61.090 153.180 61.060 ;
        RECT 157.640 61.085 162.120 61.090 ;
        POLYGON 157.640 61.085 157.690 61.085 157.690 61.080 ;
        RECT 157.690 61.080 162.120 61.085 ;
        POLYGON 162.120 61.270 162.460 61.080 162.120 61.080 ;
        POLYGON 166.335 61.270 166.390 61.270 166.390 61.220 ;
        RECT 166.390 61.220 171.435 61.270 ;
        POLYGON 166.390 61.220 166.515 61.220 166.515 61.100 ;
        RECT 166.515 61.100 171.435 61.220 ;
        POLYGON 166.515 61.100 166.535 61.100 166.535 61.080 ;
        RECT 166.535 61.080 171.435 61.100 ;
        POLYGON 157.695 61.080 157.830 61.080 157.830 61.060 ;
        RECT 157.830 61.060 162.460 61.080 ;
        POLYGON 148.800 61.060 148.800 60.980 148.680 60.980 ;
        RECT 148.800 61.050 153.090 61.060 ;
        POLYGON 153.090 61.060 153.175 61.060 153.090 61.050 ;
        POLYGON 157.830 61.060 157.900 61.060 157.900 61.050 ;
        RECT 157.900 61.050 162.460 61.060 ;
        RECT 148.800 61.045 153.060 61.050 ;
        POLYGON 153.060 61.050 153.090 61.050 153.060 61.045 ;
        POLYGON 157.900 61.050 157.920 61.050 157.920 61.045 ;
        RECT 157.920 61.045 162.460 61.050 ;
        RECT 148.800 61.015 152.910 61.045 ;
        POLYGON 152.910 61.045 153.055 61.045 152.910 61.015 ;
        POLYGON 157.920 61.045 157.940 61.045 157.940 61.040 ;
        RECT 157.940 61.040 162.460 61.045 ;
        POLYGON 157.945 61.040 158.075 61.040 158.075 61.015 ;
        RECT 158.075 61.015 162.460 61.040 ;
        RECT 148.800 61.000 152.830 61.015 ;
        POLYGON 152.830 61.015 152.905 61.015 152.830 61.000 ;
        POLYGON 158.075 61.015 158.160 61.015 158.160 61.000 ;
        RECT 158.160 61.000 162.460 61.015 ;
        RECT 148.800 60.980 152.750 61.000 ;
        POLYGON 152.750 61.000 152.830 61.000 152.750 60.980 ;
        POLYGON 158.160 61.000 158.170 61.000 158.170 60.995 ;
        RECT 158.170 60.995 162.460 61.000 ;
        POLYGON 158.170 60.995 158.210 60.995 158.210 60.990 ;
        RECT 158.210 60.990 162.460 60.995 ;
        POLYGON 158.210 60.990 158.240 60.990 158.240 60.980 ;
        RECT 158.240 60.980 162.460 60.990 ;
        POLYGON 148.680 60.980 148.680 60.960 148.650 60.960 ;
        RECT 148.680 60.960 152.655 60.980 ;
        POLYGON 145.230 60.960 145.250 60.880 145.230 60.880 ;
        RECT 117.570 60.810 145.250 60.880 ;
        POLYGON 148.650 60.960 148.650 60.875 148.520 60.875 ;
        RECT 148.650 60.955 152.655 60.960 ;
        POLYGON 152.655 60.980 152.750 60.980 152.655 60.955 ;
        POLYGON 158.240 60.980 158.345 60.980 158.345 60.955 ;
        RECT 158.345 60.955 162.460 60.980 ;
        RECT 148.650 60.940 152.575 60.955 ;
        POLYGON 152.575 60.955 152.655 60.955 152.575 60.940 ;
        POLYGON 158.345 60.955 158.410 60.955 158.410 60.940 ;
        RECT 158.410 60.940 162.460 60.955 ;
        RECT 148.650 60.905 152.470 60.940 ;
        POLYGON 152.470 60.940 152.575 60.940 152.470 60.905 ;
        POLYGON 158.410 60.940 158.525 60.940 158.525 60.905 ;
        RECT 158.525 60.905 162.460 60.940 ;
        POLYGON 162.460 61.080 162.740 60.905 162.460 60.905 ;
        POLYGON 166.535 61.080 166.665 61.080 166.665 60.960 ;
        RECT 166.665 60.960 171.435 61.080 ;
        POLYGON 166.665 60.960 166.725 60.960 166.725 60.905 ;
        RECT 166.725 60.905 171.435 60.960 ;
        RECT 148.650 60.890 152.420 60.905 ;
        POLYGON 152.420 60.905 152.465 60.905 152.420 60.890 ;
        POLYGON 158.525 60.905 158.575 60.905 158.575 60.890 ;
        RECT 158.575 60.890 162.740 60.905 ;
        RECT 148.650 60.875 152.325 60.890 ;
        POLYGON 148.520 60.875 148.520 60.870 148.510 60.870 ;
        RECT 148.520 60.870 152.325 60.875 ;
        POLYGON 145.250 60.870 145.265 60.810 145.250 60.810 ;
        RECT 117.570 60.710 145.265 60.810 ;
        POLYGON 148.510 60.870 148.510 60.790 148.390 60.790 ;
        RECT 148.510 60.865 152.325 60.870 ;
        POLYGON 152.325 60.890 152.415 60.890 152.325 60.865 ;
        POLYGON 158.575 60.890 158.660 60.890 158.660 60.865 ;
        RECT 158.660 60.865 162.740 60.890 ;
        RECT 148.510 60.825 152.200 60.865 ;
        POLYGON 152.200 60.865 152.325 60.865 152.200 60.825 ;
        POLYGON 158.660 60.865 158.765 60.865 158.765 60.830 ;
        RECT 158.765 60.830 162.740 60.865 ;
        POLYGON 158.770 60.830 158.780 60.830 158.780 60.825 ;
        RECT 158.780 60.825 162.740 60.830 ;
        RECT 148.510 60.805 152.150 60.825 ;
        POLYGON 152.150 60.825 152.200 60.825 152.150 60.805 ;
        POLYGON 158.785 60.825 158.840 60.825 158.840 60.805 ;
        RECT 158.840 60.815 162.740 60.825 ;
        POLYGON 162.740 60.905 162.880 60.815 162.740 60.815 ;
        POLYGON 166.725 60.905 166.825 60.905 166.825 60.815 ;
        RECT 166.825 60.815 171.435 60.905 ;
        RECT 158.840 60.805 162.880 60.815 ;
        RECT 148.510 60.790 152.070 60.805 ;
        POLYGON 145.265 60.790 145.285 60.710 145.265 60.710 ;
        POLYGON 148.390 60.790 148.390 60.710 148.280 60.710 ;
        RECT 148.390 60.780 152.070 60.790 ;
        POLYGON 152.070 60.805 152.150 60.805 152.070 60.780 ;
        POLYGON 158.840 60.805 158.915 60.805 158.915 60.780 ;
        RECT 158.915 60.790 162.880 60.805 ;
        POLYGON 162.880 60.815 162.920 60.790 162.880 60.790 ;
        POLYGON 166.825 60.815 166.850 60.815 166.850 60.790 ;
        RECT 166.850 60.790 171.435 60.815 ;
        RECT 158.915 60.780 162.920 60.790 ;
        RECT 148.390 60.730 151.945 60.780 ;
        POLYGON 151.945 60.780 152.070 60.780 151.945 60.730 ;
        POLYGON 158.915 60.780 159.020 60.780 159.020 60.740 ;
        RECT 159.020 60.740 162.920 60.780 ;
        POLYGON 159.025 60.740 159.050 60.740 159.050 60.730 ;
        RECT 159.050 60.730 162.920 60.740 ;
        RECT 148.390 60.715 151.910 60.730 ;
        POLYGON 151.910 60.730 151.935 60.730 151.910 60.715 ;
        POLYGON 159.050 60.730 159.085 60.730 159.085 60.715 ;
        RECT 159.085 60.715 162.920 60.730 ;
        RECT 148.390 60.710 151.805 60.715 ;
        RECT 117.570 60.640 145.285 60.710 ;
        POLYGON 148.280 60.710 148.280 60.705 148.275 60.705 ;
        RECT 148.280 60.705 151.805 60.710 ;
        POLYGON 148.275 60.705 148.275 60.695 148.260 60.695 ;
        RECT 148.275 60.695 151.805 60.705 ;
        POLYGON 145.285 60.695 145.300 60.640 145.285 60.640 ;
        POLYGON 148.260 60.695 148.260 60.640 148.180 60.640 ;
        RECT 148.260 60.680 151.805 60.695 ;
        POLYGON 151.805 60.715 151.910 60.715 151.805 60.680 ;
        POLYGON 159.085 60.715 159.180 60.715 159.180 60.680 ;
        RECT 159.180 60.680 162.920 60.715 ;
        RECT 148.260 60.640 151.700 60.680 ;
        RECT 117.570 60.525 145.300 60.640 ;
        RECT 117.500 60.520 145.300 60.525 ;
        POLYGON 145.300 60.640 145.325 60.520 145.300 60.520 ;
        POLYGON 148.180 60.640 148.180 60.520 148.010 60.520 ;
        RECT 148.180 60.630 151.700 60.640 ;
        POLYGON 151.700 60.680 151.805 60.680 151.700 60.630 ;
        POLYGON 159.180 60.680 159.200 60.680 159.200 60.670 ;
        RECT 159.200 60.670 162.920 60.680 ;
        POLYGON 159.200 60.670 159.275 60.670 159.275 60.640 ;
        RECT 159.275 60.640 162.920 60.670 ;
        POLYGON 159.275 60.640 159.295 60.640 159.295 60.630 ;
        RECT 159.295 60.630 162.920 60.640 ;
        RECT 148.180 60.620 151.675 60.630 ;
        POLYGON 151.675 60.630 151.700 60.630 151.675 60.620 ;
        POLYGON 159.295 60.630 159.320 60.630 159.320 60.620 ;
        RECT 159.320 60.620 162.920 60.630 ;
        RECT 148.180 60.530 151.465 60.620 ;
        POLYGON 151.465 60.620 151.675 60.620 151.465 60.530 ;
        POLYGON 159.320 60.620 159.445 60.620 159.445 60.565 ;
        RECT 159.445 60.565 162.920 60.620 ;
        POLYGON 159.445 60.565 159.515 60.565 159.515 60.535 ;
        RECT 159.515 60.555 162.920 60.565 ;
        POLYGON 162.920 60.790 163.265 60.555 162.920 60.555 ;
        POLYGON 166.850 60.790 166.930 60.790 166.930 60.710 ;
        RECT 166.930 60.720 171.435 60.790 ;
        POLYGON 171.435 61.285 171.875 60.720 171.435 60.720 ;
        POLYGON 179.120 61.285 179.200 61.285 179.200 61.165 ;
        RECT 179.200 61.165 193.750 61.285 ;
        POLYGON 179.200 61.165 179.410 61.165 179.410 60.825 ;
        RECT 179.410 60.825 193.750 61.165 ;
        POLYGON 179.410 60.825 179.465 60.825 179.465 60.725 ;
        RECT 179.465 60.720 193.750 60.825 ;
        RECT 166.930 60.710 171.875 60.720 ;
        POLYGON 166.930 60.710 167.020 60.710 167.020 60.615 ;
        RECT 167.020 60.615 171.875 60.710 ;
        POLYGON 167.020 60.615 167.080 60.615 167.080 60.555 ;
        RECT 167.080 60.590 171.875 60.615 ;
        POLYGON 171.875 60.720 171.980 60.590 171.875 60.590 ;
        POLYGON 179.465 60.720 179.540 60.720 179.540 60.590 ;
        RECT 179.540 60.590 193.750 60.720 ;
        RECT 167.080 60.555 171.980 60.590 ;
        RECT 159.515 60.540 163.265 60.555 ;
        POLYGON 163.265 60.555 163.285 60.540 163.265 60.540 ;
        POLYGON 167.080 60.555 167.095 60.555 167.095 60.540 ;
        RECT 167.095 60.540 171.980 60.555 ;
        RECT 159.515 60.535 163.285 60.540 ;
        POLYGON 159.515 60.535 159.525 60.535 159.525 60.530 ;
        RECT 159.525 60.530 163.285 60.535 ;
        RECT 148.180 60.525 151.460 60.530 ;
        RECT 148.180 60.520 151.445 60.525 ;
        POLYGON 151.445 60.525 151.460 60.525 151.445 60.520 ;
        POLYGON 159.525 60.530 159.545 60.530 159.545 60.520 ;
        RECT 159.545 60.520 163.285 60.530 ;
        POLYGON 117.500 60.495 117.500 60.455 117.495 60.455 ;
        RECT 117.500 60.470 145.325 60.520 ;
        POLYGON 148.010 60.520 148.010 60.510 147.995 60.510 ;
        RECT 148.010 60.510 151.235 60.520 ;
        POLYGON 145.325 60.510 145.335 60.470 145.325 60.470 ;
        RECT 117.500 60.455 145.335 60.470 ;
        RECT 50.380 60.015 111.200 60.450 ;
        POLYGON 111.200 60.450 111.225 60.450 111.200 60.015 ;
        POLYGON 117.495 60.445 117.495 60.395 117.490 60.395 ;
        RECT 117.495 60.420 145.335 60.455 ;
        POLYGON 147.995 60.510 147.995 60.450 147.920 60.450 ;
        RECT 147.995 60.450 151.235 60.510 ;
        POLYGON 145.335 60.450 145.345 60.420 145.335 60.420 ;
        RECT 117.495 60.395 145.345 60.420 ;
        POLYGON 147.920 60.450 147.920 60.415 147.875 60.415 ;
        RECT 147.920 60.430 151.235 60.450 ;
        POLYGON 151.235 60.520 151.445 60.520 151.235 60.430 ;
        POLYGON 159.545 60.520 159.695 60.520 159.695 60.455 ;
        RECT 159.695 60.495 163.285 60.520 ;
        POLYGON 163.285 60.540 163.350 60.495 163.285 60.495 ;
        POLYGON 167.095 60.540 167.110 60.540 167.110 60.530 ;
        RECT 167.110 60.530 171.980 60.540 ;
        POLYGON 167.110 60.530 167.140 60.530 167.140 60.495 ;
        RECT 167.140 60.495 171.980 60.530 ;
        RECT 159.695 60.455 163.350 60.495 ;
        POLYGON 159.700 60.455 159.750 60.455 159.750 60.430 ;
        RECT 159.750 60.430 163.350 60.455 ;
        RECT 147.920 60.425 151.225 60.430 ;
        POLYGON 151.225 60.430 151.235 60.430 151.225 60.425 ;
        POLYGON 159.750 60.430 159.760 60.430 159.760 60.425 ;
        RECT 159.760 60.425 163.350 60.430 ;
        RECT 147.920 60.420 151.220 60.425 ;
        POLYGON 151.220 60.425 151.225 60.425 151.220 60.420 ;
        POLYGON 159.760 60.425 159.770 60.425 159.770 60.420 ;
        RECT 159.770 60.420 163.350 60.425 ;
        RECT 147.920 60.415 150.995 60.420 ;
        POLYGON 147.875 60.415 147.875 60.405 147.860 60.405 ;
        RECT 147.875 60.405 150.995 60.415 ;
        POLYGON 117.490 60.385 117.490 60.035 117.465 60.035 ;
        RECT 117.490 60.350 145.345 60.395 ;
        POLYGON 145.345 60.405 145.360 60.350 145.345 60.350 ;
        POLYGON 147.860 60.405 147.860 60.350 147.790 60.350 ;
        RECT 147.860 60.350 150.995 60.405 ;
        RECT 117.490 60.220 145.360 60.350 ;
        POLYGON 145.360 60.350 145.390 60.220 145.360 60.220 ;
        RECT 117.490 60.180 145.390 60.220 ;
        POLYGON 147.790 60.350 147.790 60.210 147.605 60.210 ;
        RECT 147.790 60.315 150.995 60.350 ;
        POLYGON 150.995 60.420 151.220 60.420 150.995 60.315 ;
        POLYGON 159.770 60.420 159.930 60.420 159.930 60.345 ;
        RECT 159.930 60.345 163.350 60.420 ;
        POLYGON 159.930 60.345 159.990 60.345 159.990 60.315 ;
        RECT 159.990 60.315 163.350 60.345 ;
        RECT 147.790 60.305 150.980 60.315 ;
        POLYGON 150.980 60.315 150.995 60.315 150.980 60.305 ;
        POLYGON 159.990 60.315 160.010 60.315 160.010 60.305 ;
        RECT 160.010 60.305 163.350 60.315 ;
        RECT 147.790 60.250 150.860 60.305 ;
        POLYGON 150.860 60.305 150.980 60.305 150.860 60.250 ;
        POLYGON 160.010 60.305 160.130 60.305 160.130 60.250 ;
        RECT 160.130 60.250 163.350 60.305 ;
        POLYGON 163.350 60.495 163.685 60.250 163.350 60.250 ;
        POLYGON 167.140 60.495 167.180 60.495 167.180 60.455 ;
        RECT 167.180 60.470 171.980 60.495 ;
        POLYGON 171.980 60.590 172.060 60.470 171.980 60.470 ;
        POLYGON 179.540 60.590 179.605 60.590 179.605 60.470 ;
        RECT 179.605 60.470 193.750 60.590 ;
        RECT 167.180 60.455 172.060 60.470 ;
        POLYGON 167.180 60.455 167.375 60.455 167.375 60.255 ;
        RECT 167.375 60.250 172.060 60.455 ;
        RECT 147.790 60.210 150.570 60.250 ;
        POLYGON 145.390 60.210 145.400 60.180 145.390 60.180 ;
        RECT 117.490 60.135 145.400 60.180 ;
        POLYGON 147.605 60.210 147.605 60.160 147.550 60.160 ;
        RECT 147.605 60.160 150.570 60.210 ;
        POLYGON 145.400 60.160 145.410 60.135 145.400 60.135 ;
        POLYGON 147.550 60.160 147.550 60.135 147.515 60.135 ;
        RECT 147.550 60.135 150.570 60.160 ;
        RECT 117.490 60.035 145.410 60.135 ;
        POLYGON 147.515 60.135 147.515 60.130 147.510 60.130 ;
        RECT 147.515 60.130 150.570 60.135 ;
        RECT 50.380 60.000 111.175 60.015 ;
        RECT 5.000 58.000 27.000 60.000 ;
        POLYGON 50.380 60.000 50.710 60.000 50.710 58.490 ;
        RECT 50.710 58.490 111.175 60.000 ;
        POLYGON 50.710 58.490 50.815 58.490 50.815 58.110 ;
        RECT 50.815 58.110 111.175 58.490 ;
        POLYGON 50.815 58.110 50.845 58.110 50.845 58.000 ;
        RECT 50.845 58.000 111.175 58.110 ;
        RECT 5.000 50.000 25.000 58.000 ;
        POLYGON 50.845 58.000 51.940 58.000 51.940 54.005 ;
        RECT 51.940 56.390 111.175 58.000 ;
        POLYGON 111.175 60.015 111.200 60.015 111.175 57.055 ;
        POLYGON 117.465 60.015 117.465 59.750 117.445 59.750 ;
        RECT 117.465 60.010 145.410 60.035 ;
        POLYGON 145.410 60.130 145.440 60.010 145.410 60.010 ;
        RECT 117.465 59.925 145.440 60.010 ;
        POLYGON 147.510 60.130 147.510 59.995 147.350 59.995 ;
        RECT 147.510 60.110 150.570 60.130 ;
        POLYGON 150.570 60.250 150.860 60.250 150.570 60.110 ;
        POLYGON 160.130 60.250 160.185 60.250 160.185 60.225 ;
        RECT 160.185 60.220 163.685 60.250 ;
        POLYGON 160.185 60.220 160.390 60.220 160.390 60.125 ;
        RECT 160.390 60.125 163.685 60.220 ;
        POLYGON 160.390 60.125 160.415 60.125 160.415 60.110 ;
        RECT 160.415 60.110 163.685 60.125 ;
        RECT 147.510 60.095 150.540 60.110 ;
        POLYGON 150.540 60.110 150.570 60.110 150.540 60.095 ;
        POLYGON 160.415 60.110 160.445 60.110 160.445 60.095 ;
        RECT 160.445 60.095 163.685 60.110 ;
        RECT 147.510 60.070 150.495 60.095 ;
        POLYGON 150.495 60.095 150.540 60.095 150.495 60.070 ;
        POLYGON 160.445 60.095 160.495 60.095 160.495 60.070 ;
        RECT 160.495 60.070 163.685 60.095 ;
        RECT 147.510 60.065 150.485 60.070 ;
        POLYGON 150.485 60.070 150.495 60.070 150.485 60.065 ;
        POLYGON 160.495 60.070 160.500 60.070 160.500 60.065 ;
        RECT 160.500 60.065 163.685 60.070 ;
        RECT 147.510 59.995 150.135 60.065 ;
        POLYGON 145.440 59.995 145.460 59.925 145.440 59.925 ;
        RECT 117.465 59.905 145.460 59.925 ;
        POLYGON 147.350 59.995 147.350 59.910 147.250 59.910 ;
        RECT 147.350 59.910 150.135 59.995 ;
        POLYGON 145.460 59.910 145.465 59.905 145.460 59.905 ;
        RECT 117.465 59.860 145.465 59.905 ;
        POLYGON 147.250 59.910 147.250 59.895 147.230 59.895 ;
        RECT 147.250 59.895 150.135 59.910 ;
        POLYGON 145.465 59.895 145.475 59.860 145.465 59.860 ;
        POLYGON 147.230 59.895 147.230 59.860 147.190 59.860 ;
        RECT 147.230 59.880 150.135 59.895 ;
        POLYGON 150.135 60.065 150.480 60.065 150.135 59.880 ;
        POLYGON 160.500 60.065 160.660 60.065 160.660 59.985 ;
        RECT 160.660 60.050 163.685 60.065 ;
        POLYGON 163.685 60.250 163.940 60.050 163.685 60.050 ;
        POLYGON 167.375 60.250 167.415 60.250 167.415 60.210 ;
        RECT 167.415 60.210 172.060 60.250 ;
        POLYGON 167.415 60.210 167.555 60.210 167.555 60.050 ;
        RECT 167.555 60.165 172.060 60.210 ;
        POLYGON 172.060 60.470 172.270 60.165 172.060 60.165 ;
        POLYGON 179.605 60.470 179.775 60.470 179.775 60.165 ;
        RECT 179.775 60.165 193.750 60.470 ;
        RECT 167.555 60.050 172.270 60.165 ;
        RECT 160.660 60.005 163.940 60.050 ;
        POLYGON 163.940 60.050 164.000 60.005 163.940 60.005 ;
        POLYGON 167.555 60.050 167.595 60.050 167.595 60.005 ;
        RECT 167.595 60.005 172.270 60.050 ;
        RECT 160.660 59.985 164.000 60.005 ;
        POLYGON 160.665 59.985 160.750 59.985 160.750 59.940 ;
        RECT 160.750 59.955 164.000 59.985 ;
        POLYGON 164.000 60.005 164.060 59.955 164.000 59.955 ;
        POLYGON 167.595 60.005 167.620 60.005 167.620 59.980 ;
        RECT 167.620 59.980 172.270 60.005 ;
        POLYGON 167.620 59.980 167.635 59.980 167.635 59.960 ;
        RECT 167.635 59.955 172.270 59.980 ;
        RECT 160.750 59.950 164.060 59.955 ;
        POLYGON 164.060 59.955 164.065 59.950 164.060 59.950 ;
        POLYGON 167.635 59.955 167.640 59.955 167.640 59.950 ;
        RECT 167.640 59.950 172.270 59.955 ;
        RECT 160.750 59.940 164.065 59.950 ;
        POLYGON 155.370 59.940 155.370 59.935 154.915 59.935 ;
        RECT 155.370 59.935 155.420 59.940 ;
        POLYGON 155.420 59.940 155.495 59.935 155.420 59.935 ;
        POLYGON 160.750 59.940 160.760 59.940 160.760 59.935 ;
        RECT 160.760 59.935 164.065 59.940 ;
        POLYGON 154.850 59.935 154.850 59.925 154.655 59.925 ;
        RECT 154.850 59.925 155.495 59.935 ;
        POLYGON 154.645 59.925 154.645 59.910 154.410 59.910 ;
        RECT 154.645 59.915 155.495 59.925 ;
        POLYGON 155.495 59.935 155.975 59.915 155.495 59.915 ;
        POLYGON 160.760 59.935 160.800 59.935 160.800 59.915 ;
        RECT 160.800 59.915 164.065 59.935 ;
        RECT 154.645 59.910 155.995 59.915 ;
        POLYGON 155.995 59.915 156.065 59.910 155.995 59.910 ;
        POLYGON 160.800 59.915 160.810 59.915 160.810 59.910 ;
        RECT 160.810 59.910 164.065 59.915 ;
        POLYGON 154.400 59.910 154.400 59.905 154.280 59.905 ;
        RECT 154.400 59.905 156.065 59.910 ;
        POLYGON 154.280 59.905 154.280 59.880 154.050 59.880 ;
        RECT 154.280 59.885 156.065 59.905 ;
        POLYGON 156.065 59.910 156.330 59.885 156.065 59.885 ;
        POLYGON 160.810 59.910 160.835 59.910 160.835 59.895 ;
        RECT 160.835 59.895 164.065 59.910 ;
        POLYGON 160.835 59.895 160.860 59.895 160.860 59.885 ;
        RECT 160.860 59.885 164.065 59.895 ;
        RECT 154.280 59.880 156.335 59.885 ;
        POLYGON 156.335 59.885 156.375 59.880 156.335 59.880 ;
        POLYGON 160.860 59.885 160.865 59.885 160.865 59.880 ;
        RECT 160.865 59.880 164.065 59.885 ;
        RECT 147.230 59.860 150.090 59.880 ;
        RECT 117.465 59.775 145.475 59.860 ;
        POLYGON 145.475 59.860 145.495 59.775 145.475 59.775 ;
        RECT 117.465 59.750 145.495 59.775 ;
        POLYGON 147.190 59.860 147.190 59.770 147.090 59.770 ;
        RECT 147.190 59.855 150.090 59.860 ;
        POLYGON 150.090 59.880 150.135 59.880 150.090 59.855 ;
        POLYGON 154.050 59.880 154.050 59.870 153.955 59.870 ;
        RECT 154.050 59.870 156.375 59.880 ;
        POLYGON 153.950 59.870 153.950 59.865 153.905 59.865 ;
        RECT 153.950 59.865 156.375 59.870 ;
        POLYGON 156.375 59.880 156.550 59.865 156.375 59.865 ;
        POLYGON 160.865 59.880 160.895 59.880 160.895 59.865 ;
        RECT 160.895 59.865 164.065 59.880 ;
        POLYGON 153.900 59.865 153.900 59.855 153.820 59.855 ;
        RECT 153.900 59.860 156.555 59.865 ;
        POLYGON 156.555 59.865 156.570 59.860 156.555 59.860 ;
        POLYGON 160.895 59.865 160.905 59.865 160.905 59.860 ;
        RECT 160.905 59.860 164.065 59.865 ;
        RECT 153.900 59.855 156.570 59.860 ;
        RECT 147.190 59.775 149.940 59.855 ;
        POLYGON 149.940 59.855 150.090 59.855 149.940 59.775 ;
        POLYGON 153.820 59.855 153.820 59.845 153.735 59.845 ;
        RECT 153.820 59.850 156.570 59.855 ;
        POLYGON 156.570 59.860 156.660 59.850 156.570 59.850 ;
        POLYGON 160.905 59.860 160.920 59.860 160.920 59.850 ;
        RECT 160.920 59.850 164.065 59.860 ;
        RECT 153.820 59.845 156.660 59.850 ;
        POLYGON 153.725 59.845 153.725 59.830 153.650 59.830 ;
        RECT 153.725 59.830 156.660 59.845 ;
        POLYGON 153.645 59.830 153.645 59.790 153.400 59.790 ;
        RECT 153.645 59.815 156.660 59.830 ;
        POLYGON 156.660 59.850 156.925 59.815 156.660 59.815 ;
        POLYGON 160.920 59.850 160.985 59.850 160.985 59.815 ;
        RECT 160.985 59.815 164.065 59.850 ;
        RECT 153.645 59.800 156.930 59.815 ;
        POLYGON 156.930 59.815 157.035 59.800 156.930 59.800 ;
        POLYGON 160.985 59.815 161.010 59.815 161.010 59.800 ;
        RECT 161.010 59.800 164.065 59.815 ;
        RECT 153.645 59.790 157.035 59.800 ;
        POLYGON 157.035 59.800 157.095 59.790 157.035 59.790 ;
        POLYGON 161.010 59.800 161.030 59.800 161.030 59.790 ;
        RECT 161.030 59.790 164.065 59.800 ;
        POLYGON 153.395 59.790 153.395 59.785 153.360 59.785 ;
        RECT 153.395 59.785 157.105 59.790 ;
        POLYGON 157.105 59.790 157.140 59.785 157.105 59.785 ;
        POLYGON 161.030 59.790 161.040 59.790 161.040 59.785 ;
        RECT 161.040 59.785 164.065 59.790 ;
        POLYGON 153.360 59.785 153.360 59.775 153.300 59.775 ;
        RECT 153.360 59.775 157.140 59.785 ;
        POLYGON 157.140 59.785 157.185 59.775 157.140 59.775 ;
        POLYGON 161.040 59.785 161.055 59.785 161.055 59.775 ;
        RECT 161.055 59.775 164.065 59.785 ;
        RECT 147.190 59.770 149.885 59.775 ;
        POLYGON 117.445 59.725 117.445 59.000 117.390 59.000 ;
        RECT 117.445 59.715 145.495 59.750 ;
        POLYGON 145.495 59.770 145.510 59.715 145.495 59.715 ;
        RECT 117.445 59.650 145.510 59.715 ;
        POLYGON 147.090 59.770 147.090 59.705 147.020 59.705 ;
        RECT 147.090 59.750 149.885 59.770 ;
        POLYGON 149.885 59.775 149.940 59.775 149.885 59.750 ;
        POLYGON 153.300 59.775 153.300 59.755 153.180 59.755 ;
        RECT 153.300 59.755 157.190 59.775 ;
        POLYGON 153.175 59.755 153.175 59.750 153.155 59.750 ;
        RECT 153.175 59.750 157.190 59.755 ;
        RECT 147.090 59.705 149.780 59.750 ;
        POLYGON 145.510 59.705 145.525 59.650 145.510 59.650 ;
        POLYGON 147.020 59.705 147.020 59.650 146.960 59.650 ;
        RECT 147.020 59.685 149.780 59.705 ;
        POLYGON 149.780 59.750 149.885 59.750 149.780 59.685 ;
        POLYGON 153.155 59.750 153.155 59.735 153.090 59.735 ;
        RECT 153.155 59.735 157.190 59.750 ;
        POLYGON 153.090 59.735 153.090 59.730 153.055 59.730 ;
        RECT 153.090 59.730 157.190 59.735 ;
        POLYGON 153.055 59.730 153.055 59.695 152.905 59.695 ;
        RECT 153.055 59.725 157.190 59.730 ;
        POLYGON 157.190 59.775 157.440 59.725 157.190 59.725 ;
        POLYGON 161.055 59.775 161.130 59.775 161.130 59.735 ;
        RECT 161.130 59.735 164.065 59.775 ;
        POLYGON 161.130 59.735 161.145 59.735 161.145 59.725 ;
        RECT 161.145 59.725 164.065 59.735 ;
        RECT 153.055 59.695 157.440 59.725 ;
        POLYGON 152.905 59.695 152.905 59.685 152.855 59.685 ;
        RECT 152.905 59.690 157.440 59.695 ;
        POLYGON 157.440 59.725 157.625 59.690 157.440 59.690 ;
        POLYGON 161.145 59.725 161.195 59.725 161.195 59.700 ;
        RECT 161.195 59.700 164.065 59.725 ;
        POLYGON 161.195 59.700 161.210 59.700 161.210 59.690 ;
        RECT 161.210 59.690 164.065 59.700 ;
        RECT 152.905 59.685 157.640 59.690 ;
        RECT 147.020 59.650 149.650 59.685 ;
        RECT 117.445 59.610 145.525 59.650 ;
        POLYGON 145.525 59.650 145.535 59.610 145.525 59.610 ;
        RECT 117.445 59.590 145.535 59.610 ;
        POLYGON 146.960 59.650 146.960 59.605 146.910 59.605 ;
        RECT 146.960 59.605 149.650 59.650 ;
        POLYGON 149.650 59.685 149.780 59.685 149.650 59.605 ;
        POLYGON 152.855 59.685 152.855 59.680 152.830 59.680 ;
        RECT 152.855 59.680 157.640 59.685 ;
        POLYGON 157.640 59.690 157.690 59.680 157.640 59.680 ;
        POLYGON 161.210 59.690 161.225 59.690 161.225 59.680 ;
        RECT 161.225 59.680 164.065 59.690 ;
        POLYGON 152.830 59.680 152.830 59.665 152.750 59.665 ;
        RECT 152.830 59.665 157.695 59.680 ;
        POLYGON 161.225 59.680 161.230 59.680 161.230 59.675 ;
        RECT 161.230 59.675 164.065 59.680 ;
        POLYGON 152.750 59.665 152.750 59.640 152.655 59.640 ;
        RECT 152.750 59.640 157.695 59.665 ;
        POLYGON 152.655 59.640 152.655 59.620 152.575 59.620 ;
        RECT 152.655 59.630 157.695 59.640 ;
        POLYGON 157.695 59.675 157.895 59.630 157.695 59.630 ;
        POLYGON 161.230 59.675 161.265 59.675 161.265 59.655 ;
        RECT 161.265 59.655 164.065 59.675 ;
        POLYGON 161.265 59.655 161.305 59.655 161.305 59.630 ;
        RECT 161.305 59.635 164.065 59.655 ;
        POLYGON 164.065 59.950 164.435 59.635 164.065 59.635 ;
        POLYGON 167.640 59.950 167.840 59.950 167.840 59.730 ;
        RECT 167.840 59.730 172.270 59.950 ;
        POLYGON 167.840 59.730 167.865 59.730 167.865 59.705 ;
        RECT 167.865 59.705 172.270 59.730 ;
        POLYGON 167.865 59.705 167.915 59.705 167.915 59.640 ;
        RECT 167.915 59.665 172.270 59.705 ;
        POLYGON 172.270 60.165 172.615 59.665 172.270 59.665 ;
        POLYGON 179.775 60.165 180.050 60.165 180.050 59.665 ;
        RECT 180.050 60.015 193.750 60.165 ;
        POLYGON 193.750 61.405 194.390 60.015 193.750 60.015 ;
        RECT 180.050 59.995 194.390 60.015 ;
        POLYGON 206.335 61.390 206.335 60.005 206.245 60.005 ;
        RECT 206.335 61.335 223.235 61.405 ;
        POLYGON 223.235 61.445 223.270 61.445 223.235 61.335 ;
        POLYGON 231.400 61.450 231.400 61.335 231.340 61.335 ;
        RECT 231.400 61.335 236.575 61.450 ;
        RECT 206.335 60.710 223.035 61.335 ;
        POLYGON 223.035 61.335 223.235 61.335 223.035 60.710 ;
        POLYGON 231.340 61.335 231.340 61.215 231.280 61.215 ;
        RECT 231.340 61.275 236.575 61.335 ;
        POLYGON 236.575 61.450 236.710 61.450 236.575 61.275 ;
        POLYGON 240.845 61.450 240.845 61.280 240.660 61.280 ;
        RECT 240.845 61.395 244.440 61.450 ;
        POLYGON 244.440 61.450 244.535 61.450 244.440 61.395 ;
        POLYGON 256.765 61.450 256.870 61.450 256.870 61.395 ;
        RECT 256.870 61.395 261.095 61.450 ;
        RECT 240.845 61.300 244.260 61.395 ;
        POLYGON 244.260 61.395 244.440 61.395 244.260 61.300 ;
        POLYGON 256.870 61.395 256.930 61.395 256.930 61.365 ;
        RECT 256.930 61.365 261.095 61.395 ;
        POLYGON 256.930 61.365 257.045 61.365 257.045 61.300 ;
        RECT 257.045 61.300 261.095 61.365 ;
        RECT 240.845 61.280 244.195 61.300 ;
        POLYGON 240.660 61.280 240.660 61.275 240.655 61.275 ;
        RECT 240.660 61.275 244.195 61.280 ;
        RECT 231.340 61.215 236.485 61.275 ;
        POLYGON 231.280 61.215 231.280 60.910 231.140 60.910 ;
        RECT 231.280 61.150 236.485 61.215 ;
        POLYGON 236.485 61.275 236.575 61.275 236.485 61.150 ;
        POLYGON 240.655 61.275 240.655 61.150 240.520 61.150 ;
        RECT 240.655 61.260 244.195 61.275 ;
        POLYGON 244.195 61.300 244.260 61.300 244.195 61.260 ;
        POLYGON 257.045 61.300 257.115 61.300 257.115 61.260 ;
        RECT 257.115 61.260 261.095 61.300 ;
        RECT 240.655 61.150 243.960 61.260 ;
        RECT 231.280 61.010 236.390 61.150 ;
        POLYGON 236.390 61.150 236.485 61.150 236.390 61.010 ;
        POLYGON 240.520 61.150 240.520 61.135 240.505 61.135 ;
        RECT 240.520 61.135 243.960 61.150 ;
        POLYGON 240.505 61.135 240.505 61.010 240.370 61.010 ;
        RECT 240.505 61.125 243.960 61.135 ;
        POLYGON 243.960 61.260 244.195 61.260 243.960 61.125 ;
        POLYGON 257.115 61.260 257.165 61.260 257.165 61.235 ;
        RECT 257.165 61.235 261.095 61.260 ;
        POLYGON 257.165 61.235 257.275 61.235 257.275 61.170 ;
        RECT 257.275 61.170 261.095 61.235 ;
        POLYGON 257.275 61.170 257.280 61.170 257.280 61.165 ;
        RECT 257.280 61.165 261.095 61.170 ;
        POLYGON 250.365 61.165 250.365 61.160 249.785 61.160 ;
        RECT 250.365 61.160 250.620 61.165 ;
        POLYGON 250.620 61.165 251.105 61.160 250.620 61.160 ;
        POLYGON 257.280 61.165 257.290 61.165 257.290 61.160 ;
        RECT 257.290 61.160 261.095 61.165 ;
        POLYGON 249.760 61.160 249.760 61.155 249.665 61.155 ;
        RECT 249.760 61.155 251.265 61.160 ;
        POLYGON 251.265 61.160 251.345 61.155 251.265 61.155 ;
        POLYGON 257.290 61.160 257.300 61.160 257.300 61.155 ;
        RECT 257.300 61.155 261.095 61.160 ;
        POLYGON 249.610 61.155 249.610 61.145 249.370 61.145 ;
        RECT 249.610 61.150 251.480 61.155 ;
        POLYGON 251.480 61.155 251.505 61.150 251.480 61.150 ;
        POLYGON 257.300 61.155 257.305 61.155 257.305 61.150 ;
        RECT 257.305 61.150 261.095 61.155 ;
        RECT 249.610 61.145 251.530 61.150 ;
        POLYGON 251.530 61.150 251.655 61.145 251.530 61.145 ;
        POLYGON 257.305 61.150 257.315 61.150 257.315 61.145 ;
        RECT 257.315 61.145 261.095 61.150 ;
        POLYGON 249.355 61.145 249.355 61.130 248.965 61.130 ;
        RECT 249.355 61.140 251.680 61.145 ;
        POLYGON 251.680 61.145 251.855 61.140 251.680 61.140 ;
        POLYGON 257.315 61.145 257.325 61.145 257.325 61.140 ;
        RECT 257.325 61.140 261.095 61.145 ;
        RECT 249.355 61.130 251.855 61.140 ;
        POLYGON 251.855 61.140 252.040 61.130 251.855 61.130 ;
        POLYGON 257.325 61.140 257.345 61.140 257.345 61.130 ;
        RECT 257.345 61.130 261.095 61.140 ;
        POLYGON 248.965 61.130 248.965 61.125 248.910 61.125 ;
        RECT 248.965 61.125 252.090 61.130 ;
        POLYGON 252.090 61.130 252.155 61.125 252.090 61.125 ;
        POLYGON 257.345 61.130 257.350 61.130 257.350 61.125 ;
        RECT 257.350 61.125 261.095 61.130 ;
        RECT 240.505 61.120 243.955 61.125 ;
        POLYGON 243.955 61.125 243.960 61.125 243.955 61.120 ;
        POLYGON 248.905 61.125 248.905 61.120 248.810 61.120 ;
        RECT 248.905 61.120 252.155 61.125 ;
        RECT 240.505 61.050 243.840 61.120 ;
        POLYGON 243.840 61.120 243.955 61.120 243.840 61.050 ;
        POLYGON 248.805 61.120 248.805 61.110 248.660 61.110 ;
        RECT 248.805 61.110 252.155 61.120 ;
        POLYGON 252.155 61.125 252.335 61.110 252.155 61.110 ;
        POLYGON 257.350 61.125 257.375 61.125 257.375 61.110 ;
        RECT 257.375 61.110 261.095 61.125 ;
        POLYGON 248.660 61.110 248.660 61.080 248.370 61.080 ;
        RECT 248.660 61.100 252.350 61.110 ;
        POLYGON 252.350 61.110 252.435 61.100 252.350 61.100 ;
        POLYGON 257.375 61.110 257.395 61.110 257.395 61.100 ;
        RECT 257.395 61.100 261.095 61.110 ;
        RECT 248.660 61.095 252.435 61.100 ;
        POLYGON 252.435 61.100 252.500 61.095 252.435 61.095 ;
        POLYGON 257.395 61.100 257.400 61.100 257.400 61.095 ;
        RECT 257.400 61.095 261.095 61.100 ;
        RECT 248.660 61.080 252.505 61.095 ;
        POLYGON 252.505 61.095 252.635 61.080 252.505 61.080 ;
        POLYGON 257.400 61.095 257.425 61.095 257.425 61.080 ;
        RECT 257.425 61.080 261.095 61.095 ;
        POLYGON 248.370 61.080 248.370 61.070 248.315 61.070 ;
        RECT 248.370 61.070 252.635 61.080 ;
        POLYGON 252.635 61.080 252.705 61.070 252.635 61.070 ;
        POLYGON 257.425 61.080 257.445 61.080 257.445 61.070 ;
        RECT 257.445 61.070 261.095 61.080 ;
        POLYGON 248.315 61.070 248.315 61.050 248.170 61.050 ;
        RECT 248.315 61.050 252.705 61.070 ;
        RECT 240.505 61.010 243.660 61.050 ;
        RECT 231.280 60.910 236.295 61.010 ;
        POLYGON 231.140 60.910 231.140 60.710 231.050 60.710 ;
        RECT 231.140 60.875 236.295 60.910 ;
        POLYGON 236.295 61.010 236.390 61.010 236.295 60.875 ;
        POLYGON 240.370 61.010 240.370 60.980 240.335 60.980 ;
        RECT 240.370 60.980 243.660 61.010 ;
        POLYGON 240.335 60.980 240.335 60.895 240.255 60.895 ;
        RECT 240.335 60.940 243.660 60.980 ;
        POLYGON 243.660 61.050 243.840 61.050 243.660 60.940 ;
        POLYGON 248.170 61.050 248.170 61.040 248.100 61.040 ;
        RECT 248.170 61.040 252.705 61.050 ;
        POLYGON 252.705 61.070 252.905 61.040 252.705 61.040 ;
        POLYGON 257.445 61.070 257.495 61.070 257.495 61.040 ;
        RECT 257.495 61.040 261.095 61.070 ;
        POLYGON 248.100 61.040 248.100 61.030 248.055 61.030 ;
        RECT 248.100 61.035 252.905 61.040 ;
        POLYGON 252.905 61.040 252.915 61.035 252.905 61.035 ;
        POLYGON 257.495 61.040 257.500 61.040 257.500 61.035 ;
        RECT 257.500 61.035 261.095 61.040 ;
        RECT 248.100 61.030 252.915 61.035 ;
        POLYGON 248.055 61.030 248.055 61.020 247.995 61.020 ;
        RECT 248.055 61.025 252.915 61.030 ;
        POLYGON 252.915 61.035 252.970 61.025 252.915 61.025 ;
        POLYGON 257.500 61.035 257.520 61.035 257.520 61.025 ;
        RECT 257.520 61.025 261.095 61.035 ;
        RECT 248.055 61.020 252.970 61.025 ;
        POLYGON 247.995 61.020 247.995 60.990 247.840 60.990 ;
        RECT 247.995 60.990 252.970 61.020 ;
        POLYGON 252.970 61.025 253.165 60.990 252.970 60.990 ;
        POLYGON 257.520 61.025 257.575 61.025 257.575 60.990 ;
        RECT 257.575 60.990 261.095 61.025 ;
        POLYGON 247.840 60.990 247.840 60.940 247.650 60.940 ;
        RECT 247.840 60.985 253.165 60.990 ;
        POLYGON 253.165 60.990 253.190 60.985 253.165 60.985 ;
        POLYGON 257.575 60.990 257.585 60.990 257.585 60.985 ;
        RECT 257.585 60.985 261.095 60.990 ;
        RECT 247.840 60.975 253.195 60.985 ;
        POLYGON 253.195 60.985 253.230 60.975 253.195 60.975 ;
        POLYGON 257.585 60.985 257.605 60.985 257.605 60.975 ;
        RECT 257.605 60.975 261.095 60.985 ;
        RECT 247.840 60.950 253.235 60.975 ;
        POLYGON 253.235 60.975 253.325 60.950 253.235 60.950 ;
        POLYGON 257.605 60.975 257.615 60.975 257.615 60.970 ;
        RECT 257.615 60.970 261.095 60.975 ;
        POLYGON 257.615 60.970 257.645 60.970 257.645 60.950 ;
        RECT 257.645 60.950 261.095 60.970 ;
        RECT 247.840 60.940 253.325 60.950 ;
        RECT 240.335 60.925 243.645 60.940 ;
        POLYGON 243.645 60.940 243.660 60.940 243.645 60.925 ;
        POLYGON 247.650 60.940 247.650 60.925 247.590 60.925 ;
        RECT 247.650 60.930 253.325 60.940 ;
        POLYGON 253.325 60.950 253.415 60.930 253.325 60.930 ;
        POLYGON 257.645 60.950 257.675 60.950 257.675 60.930 ;
        RECT 257.675 60.930 261.095 60.950 ;
        RECT 247.650 60.925 253.415 60.930 ;
        RECT 240.335 60.895 243.495 60.925 ;
        POLYGON 240.255 60.895 240.255 60.875 240.235 60.875 ;
        RECT 240.255 60.875 243.495 60.895 ;
        RECT 231.140 60.710 236.145 60.875 ;
        RECT 206.335 60.485 222.965 60.710 ;
        POLYGON 222.965 60.710 223.035 60.710 222.965 60.490 ;
        POLYGON 231.050 60.710 231.050 60.610 231.005 60.610 ;
        RECT 231.050 60.660 236.145 60.710 ;
        POLYGON 236.145 60.875 236.295 60.875 236.145 60.660 ;
        POLYGON 240.235 60.875 240.235 60.660 240.030 60.660 ;
        RECT 240.235 60.830 243.495 60.875 ;
        POLYGON 243.495 60.925 243.645 60.925 243.495 60.830 ;
        POLYGON 247.590 60.925 247.590 60.895 247.485 60.895 ;
        RECT 247.590 60.905 253.415 60.925 ;
        POLYGON 253.415 60.930 253.505 60.905 253.415 60.905 ;
        POLYGON 257.675 60.930 257.710 60.930 257.710 60.905 ;
        RECT 257.710 60.905 261.095 60.930 ;
        RECT 247.590 60.895 253.505 60.905 ;
        POLYGON 247.485 60.895 247.485 60.855 247.340 60.855 ;
        RECT 247.485 60.855 253.505 60.895 ;
        POLYGON 253.505 60.905 253.670 60.855 253.505 60.855 ;
        POLYGON 257.710 60.905 257.785 60.905 257.785 60.855 ;
        RECT 257.785 60.855 261.095 60.905 ;
        POLYGON 247.335 60.855 247.335 60.830 247.265 60.830 ;
        RECT 247.335 60.830 253.670 60.855 ;
        POLYGON 253.670 60.855 253.735 60.830 253.670 60.830 ;
        POLYGON 257.785 60.855 257.825 60.855 257.825 60.830 ;
        RECT 257.825 60.850 261.095 60.855 ;
        POLYGON 261.095 61.450 261.760 60.850 261.095 60.850 ;
        POLYGON 266.295 61.450 266.365 61.450 266.365 61.365 ;
        RECT 266.365 61.365 274.045 61.450 ;
        POLYGON 266.365 61.365 266.470 61.365 266.470 61.225 ;
        RECT 266.470 61.225 274.045 61.365 ;
        POLYGON 266.470 61.225 266.490 61.225 266.490 61.205 ;
        RECT 266.490 61.205 274.045 61.225 ;
        POLYGON 266.490 61.205 266.570 61.205 266.570 61.100 ;
        RECT 266.570 61.100 274.045 61.205 ;
        POLYGON 266.570 61.100 266.580 61.100 266.580 61.085 ;
        RECT 266.580 61.085 274.045 61.100 ;
        POLYGON 266.580 61.085 266.645 61.085 266.645 61.005 ;
        RECT 266.645 61.080 274.045 61.085 ;
        POLYGON 274.045 61.450 274.275 61.080 274.045 61.080 ;
        RECT 287.575 61.405 303.120 61.780 ;
        POLYGON 287.575 61.405 287.610 61.405 287.610 61.085 ;
        RECT 287.610 61.080 303.120 61.405 ;
        RECT 266.645 61.005 274.275 61.080 ;
        POLYGON 266.645 61.005 266.650 61.005 266.650 60.995 ;
        RECT 266.650 60.995 274.275 61.005 ;
        POLYGON 266.650 60.995 266.695 60.995 266.695 60.935 ;
        RECT 266.695 60.935 274.275 60.995 ;
        POLYGON 266.695 60.935 266.700 60.935 266.700 60.930 ;
        RECT 266.700 60.930 274.275 60.935 ;
        POLYGON 266.700 60.930 266.725 60.930 266.725 60.895 ;
        RECT 266.725 60.895 274.275 60.930 ;
        POLYGON 266.725 60.895 266.740 60.895 266.740 60.880 ;
        RECT 266.740 60.880 274.275 60.895 ;
        POLYGON 266.740 60.880 266.760 60.880 266.760 60.850 ;
        RECT 266.760 60.850 274.275 60.880 ;
        RECT 257.825 60.830 261.760 60.850 ;
        RECT 240.235 60.750 243.375 60.830 ;
        POLYGON 243.375 60.830 243.495 60.830 243.375 60.750 ;
        POLYGON 247.265 60.830 247.265 60.810 247.210 60.810 ;
        RECT 247.265 60.810 253.735 60.830 ;
        POLYGON 247.200 60.810 247.200 60.785 247.130 60.785 ;
        RECT 247.200 60.785 253.735 60.810 ;
        POLYGON 247.130 60.785 247.130 60.770 247.085 60.770 ;
        RECT 247.130 60.770 253.735 60.785 ;
        POLYGON 253.735 60.830 253.925 60.770 253.735 60.770 ;
        POLYGON 257.825 60.830 257.915 60.830 257.915 60.770 ;
        RECT 257.915 60.770 261.760 60.830 ;
        POLYGON 247.085 60.770 247.085 60.750 247.035 60.750 ;
        RECT 247.085 60.750 253.925 60.770 ;
        RECT 240.235 60.660 243.190 60.750 ;
        RECT 231.050 60.610 236.055 60.660 ;
        POLYGON 231.005 60.610 231.005 60.490 230.955 60.490 ;
        RECT 231.005 60.530 236.055 60.610 ;
        POLYGON 236.055 60.660 236.145 60.660 236.055 60.530 ;
        POLYGON 240.030 60.660 240.030 60.535 239.910 60.535 ;
        RECT 240.030 60.620 243.190 60.660 ;
        POLYGON 243.190 60.750 243.375 60.750 243.190 60.620 ;
        POLYGON 247.035 60.750 247.035 60.665 246.820 60.665 ;
        RECT 247.035 60.725 253.925 60.750 ;
        POLYGON 253.925 60.770 254.045 60.725 253.925 60.725 ;
        POLYGON 257.915 60.770 257.935 60.770 257.935 60.760 ;
        RECT 257.935 60.760 261.760 60.770 ;
        POLYGON 257.935 60.760 257.985 60.760 257.985 60.725 ;
        RECT 257.985 60.725 261.760 60.760 ;
        RECT 247.035 60.705 254.045 60.725 ;
        POLYGON 254.045 60.725 254.090 60.705 254.045 60.705 ;
        POLYGON 257.985 60.725 258.010 60.725 258.010 60.710 ;
        RECT 258.010 60.710 261.760 60.725 ;
        POLYGON 258.010 60.710 258.015 60.710 258.015 60.705 ;
        RECT 258.015 60.705 261.760 60.710 ;
        RECT 247.035 60.685 254.090 60.705 ;
        POLYGON 254.090 60.705 254.140 60.685 254.090 60.685 ;
        POLYGON 258.015 60.705 258.050 60.705 258.050 60.685 ;
        RECT 258.050 60.685 261.760 60.705 ;
        RECT 247.035 60.670 254.145 60.685 ;
        POLYGON 254.145 60.685 254.185 60.670 254.145 60.670 ;
        POLYGON 258.050 60.685 258.070 60.685 258.070 60.670 ;
        RECT 258.070 60.670 261.760 60.685 ;
        RECT 247.035 60.665 254.185 60.670 ;
        POLYGON 246.820 60.665 246.820 60.660 246.805 60.660 ;
        RECT 246.820 60.660 254.185 60.665 ;
        POLYGON 246.805 60.660 246.805 60.620 246.715 60.620 ;
        RECT 246.805 60.620 254.185 60.660 ;
        RECT 240.030 60.560 243.100 60.620 ;
        POLYGON 243.100 60.620 243.190 60.620 243.100 60.560 ;
        POLYGON 246.715 60.620 246.715 60.560 246.575 60.560 ;
        RECT 246.715 60.560 254.185 60.620 ;
        RECT 240.030 60.535 242.885 60.560 ;
        RECT 231.005 60.515 236.045 60.530 ;
        POLYGON 236.045 60.530 236.055 60.530 236.045 60.515 ;
        POLYGON 239.910 60.530 239.910 60.515 239.895 60.515 ;
        RECT 239.910 60.515 242.885 60.535 ;
        RECT 231.005 60.490 236.005 60.515 ;
        RECT 206.335 60.005 222.835 60.485 ;
        POLYGON 222.835 60.485 222.965 60.485 222.835 60.010 ;
        POLYGON 230.955 60.490 230.955 60.010 230.750 60.010 ;
        RECT 230.955 60.450 236.005 60.490 ;
        POLYGON 236.005 60.515 236.045 60.515 236.005 60.450 ;
        POLYGON 239.895 60.515 239.895 60.450 239.830 60.450 ;
        RECT 239.895 60.450 242.885 60.515 ;
        RECT 230.955 60.420 235.985 60.450 ;
        POLYGON 235.985 60.450 236.005 60.450 235.985 60.420 ;
        POLYGON 239.830 60.450 239.830 60.420 239.805 60.420 ;
        RECT 239.830 60.420 242.885 60.450 ;
        RECT 230.955 60.400 235.975 60.420 ;
        POLYGON 235.975 60.420 235.985 60.420 235.975 60.400 ;
        POLYGON 239.805 60.420 239.805 60.400 239.785 60.400 ;
        RECT 239.805 60.400 242.885 60.420 ;
        POLYGON 242.885 60.560 243.100 60.560 242.885 60.400 ;
        POLYGON 246.575 60.560 246.575 60.530 246.505 60.530 ;
        RECT 246.575 60.530 254.185 60.560 ;
        POLYGON 246.505 60.530 246.505 60.495 246.420 60.495 ;
        RECT 246.505 60.510 254.185 60.530 ;
        POLYGON 254.185 60.670 254.550 60.510 254.185 60.510 ;
        POLYGON 258.070 60.670 258.135 60.670 258.135 60.625 ;
        RECT 258.135 60.655 261.760 60.670 ;
        POLYGON 261.760 60.850 261.950 60.655 261.760 60.655 ;
        POLYGON 266.760 60.850 266.830 60.850 266.830 60.765 ;
        RECT 266.830 60.765 274.275 60.850 ;
        POLYGON 266.830 60.765 266.915 60.765 266.915 60.655 ;
        RECT 266.915 60.680 274.275 60.765 ;
        POLYGON 274.275 61.080 274.500 60.680 274.275 60.680 ;
        POLYGON 287.610 61.080 287.655 61.080 287.655 60.680 ;
        RECT 287.655 60.680 303.120 61.080 ;
        RECT 266.915 60.655 274.500 60.680 ;
        RECT 258.135 60.625 261.950 60.655 ;
        POLYGON 258.135 60.625 258.245 60.625 258.245 60.545 ;
        RECT 258.245 60.545 261.950 60.625 ;
        POLYGON 258.245 60.545 258.295 60.545 258.295 60.510 ;
        RECT 258.295 60.510 261.950 60.545 ;
        RECT 246.505 60.495 254.550 60.510 ;
        POLYGON 246.420 60.495 246.420 60.475 246.380 60.475 ;
        RECT 246.420 60.475 254.550 60.495 ;
        POLYGON 246.375 60.475 246.375 60.420 246.245 60.420 ;
        RECT 246.375 60.420 254.550 60.475 ;
        POLYGON 254.550 60.510 254.755 60.420 254.550 60.420 ;
        POLYGON 258.295 60.510 258.405 60.510 258.405 60.435 ;
        RECT 258.405 60.490 261.950 60.510 ;
        POLYGON 261.950 60.655 262.115 60.490 261.950 60.490 ;
        POLYGON 266.915 60.655 266.975 60.655 266.975 60.580 ;
        RECT 266.975 60.580 274.500 60.655 ;
        POLYGON 266.975 60.580 267.015 60.580 267.015 60.515 ;
        RECT 267.015 60.515 274.500 60.580 ;
        POLYGON 267.015 60.515 267.030 60.515 267.030 60.490 ;
        RECT 267.030 60.490 274.500 60.515 ;
        RECT 258.405 60.435 262.115 60.490 ;
        POLYGON 258.410 60.435 258.425 60.435 258.425 60.420 ;
        RECT 258.425 60.420 262.115 60.435 ;
        POLYGON 246.245 60.420 246.245 60.405 246.220 60.405 ;
        RECT 246.245 60.415 254.755 60.420 ;
        POLYGON 254.755 60.420 254.770 60.415 254.755 60.415 ;
        POLYGON 258.425 60.420 258.430 60.420 258.430 60.415 ;
        RECT 258.430 60.415 262.115 60.420 ;
        RECT 246.245 60.405 254.770 60.415 ;
        POLYGON 246.220 60.405 246.220 60.400 246.210 60.400 ;
        RECT 246.220 60.400 254.770 60.405 ;
        RECT 230.955 60.065 235.765 60.400 ;
        POLYGON 235.765 60.400 235.975 60.400 235.765 60.065 ;
        POLYGON 239.785 60.400 239.785 60.375 239.760 60.375 ;
        RECT 239.785 60.375 242.840 60.400 ;
        POLYGON 239.760 60.375 239.760 60.300 239.690 60.300 ;
        RECT 239.760 60.365 242.840 60.375 ;
        POLYGON 242.840 60.400 242.885 60.400 242.840 60.365 ;
        POLYGON 246.210 60.400 246.210 60.365 246.135 60.365 ;
        RECT 246.210 60.365 254.770 60.400 ;
        RECT 239.760 60.355 242.825 60.365 ;
        POLYGON 242.825 60.365 242.840 60.365 242.825 60.355 ;
        POLYGON 246.135 60.365 246.135 60.355 246.115 60.355 ;
        RECT 246.135 60.360 254.770 60.365 ;
        POLYGON 254.770 60.415 254.885 60.360 254.770 60.360 ;
        POLYGON 258.430 60.415 258.505 60.415 258.505 60.360 ;
        RECT 258.505 60.360 262.115 60.415 ;
        RECT 246.135 60.355 254.885 60.360 ;
        RECT 239.760 60.300 242.585 60.355 ;
        POLYGON 239.690 60.300 239.690 60.280 239.670 60.280 ;
        RECT 239.690 60.280 242.585 60.300 ;
        POLYGON 239.670 60.280 239.670 60.210 239.615 60.210 ;
        RECT 239.670 60.210 242.585 60.280 ;
        POLYGON 239.615 60.210 239.615 60.065 239.490 60.065 ;
        RECT 239.615 60.165 242.585 60.210 ;
        POLYGON 242.585 60.355 242.825 60.355 242.585 60.165 ;
        POLYGON 246.115 60.355 246.115 60.320 246.040 60.320 ;
        RECT 246.115 60.325 254.885 60.355 ;
        POLYGON 254.885 60.360 254.955 60.325 254.885 60.325 ;
        POLYGON 258.505 60.360 258.545 60.360 258.545 60.330 ;
        RECT 258.545 60.330 262.115 60.360 ;
        POLYGON 258.545 60.330 258.550 60.330 258.550 60.325 ;
        RECT 258.550 60.325 262.115 60.330 ;
        RECT 246.115 60.320 254.955 60.325 ;
        POLYGON 246.040 60.320 246.040 60.270 245.945 60.270 ;
        RECT 246.040 60.270 254.955 60.320 ;
        POLYGON 245.940 60.270 245.940 60.165 245.720 60.165 ;
        RECT 245.940 60.170 254.955 60.270 ;
        POLYGON 254.955 60.325 255.280 60.170 254.955 60.170 ;
        POLYGON 258.550 60.325 258.760 60.325 258.760 60.170 ;
        RECT 258.760 60.190 262.115 60.325 ;
        POLYGON 262.115 60.490 262.405 60.190 262.115 60.190 ;
        POLYGON 267.030 60.490 267.235 60.490 267.235 60.190 ;
        RECT 267.235 60.190 274.500 60.490 ;
        RECT 258.760 60.170 262.405 60.190 ;
        RECT 245.940 60.165 255.280 60.170 ;
        RECT 239.615 60.100 242.505 60.165 ;
        POLYGON 242.505 60.165 242.585 60.165 242.505 60.100 ;
        POLYGON 245.720 60.165 245.720 60.140 245.665 60.140 ;
        RECT 245.720 60.140 255.280 60.165 ;
        POLYGON 245.665 60.140 245.665 60.135 245.660 60.135 ;
        RECT 245.665 60.135 255.280 60.140 ;
        POLYGON 255.280 60.170 255.350 60.135 255.280 60.135 ;
        POLYGON 258.760 60.170 258.790 60.170 258.790 60.150 ;
        RECT 258.790 60.150 262.405 60.170 ;
        POLYGON 258.790 60.150 258.805 60.150 258.805 60.135 ;
        RECT 258.805 60.135 262.405 60.150 ;
        POLYGON 245.660 60.135 245.660 60.100 245.580 60.100 ;
        RECT 245.660 60.100 255.355 60.135 ;
        POLYGON 255.355 60.135 255.420 60.100 255.355 60.100 ;
        POLYGON 258.805 60.135 258.830 60.135 258.830 60.115 ;
        RECT 258.830 60.115 262.405 60.135 ;
        POLYGON 258.830 60.115 258.845 60.115 258.845 60.100 ;
        RECT 258.845 60.100 262.405 60.115 ;
        RECT 239.615 60.065 242.440 60.100 ;
        RECT 230.955 60.010 235.725 60.065 ;
        POLYGON 194.390 60.005 194.395 59.995 194.390 59.995 ;
        RECT 180.050 59.720 194.395 59.995 ;
        POLYGON 194.395 59.995 194.510 59.720 194.395 59.720 ;
        RECT 180.050 59.665 194.510 59.720 ;
        RECT 167.915 59.635 172.615 59.665 ;
        RECT 161.305 59.630 164.435 59.635 ;
        RECT 152.655 59.620 157.900 59.630 ;
        POLYGON 152.575 59.620 152.575 59.605 152.525 59.605 ;
        RECT 152.575 59.615 157.900 59.620 ;
        POLYGON 157.900 59.630 157.945 59.615 157.900 59.615 ;
        POLYGON 161.305 59.630 161.330 59.630 161.330 59.615 ;
        RECT 161.330 59.615 164.435 59.630 ;
        RECT 152.575 59.605 157.950 59.615 ;
        POLYGON 145.535 59.605 145.540 59.590 145.535 59.590 ;
        POLYGON 146.910 59.605 146.910 59.590 146.895 59.590 ;
        RECT 146.910 59.590 149.435 59.605 ;
        RECT 117.445 59.570 145.540 59.590 ;
        POLYGON 145.540 59.590 145.545 59.570 145.540 59.570 ;
        RECT 117.445 59.545 145.545 59.570 ;
        POLYGON 146.895 59.590 146.895 59.565 146.865 59.565 ;
        RECT 146.895 59.565 149.435 59.590 ;
        POLYGON 145.545 59.565 145.550 59.545 145.545 59.545 ;
        POLYGON 146.865 59.565 146.865 59.545 146.845 59.545 ;
        RECT 146.865 59.545 149.435 59.565 ;
        RECT 117.445 59.380 145.550 59.545 ;
        POLYGON 145.550 59.545 145.590 59.380 145.550 59.380 ;
        RECT 117.445 59.235 145.590 59.380 ;
        POLYGON 146.845 59.545 146.845 59.375 146.670 59.375 ;
        RECT 146.845 59.475 149.435 59.545 ;
        POLYGON 149.435 59.605 149.650 59.605 149.435 59.475 ;
        POLYGON 152.525 59.605 152.525 59.590 152.470 59.590 ;
        RECT 152.525 59.590 157.950 59.605 ;
        POLYGON 152.465 59.590 152.465 59.575 152.415 59.575 ;
        RECT 152.465 59.575 157.950 59.590 ;
        POLYGON 152.415 59.575 152.415 59.550 152.325 59.550 ;
        RECT 152.415 59.565 157.950 59.575 ;
        POLYGON 157.950 59.615 158.155 59.565 157.950 59.565 ;
        POLYGON 161.330 59.615 161.415 59.615 161.415 59.565 ;
        RECT 161.415 59.565 164.435 59.615 ;
        RECT 152.415 59.560 158.160 59.565 ;
        POLYGON 158.160 59.565 158.170 59.560 158.160 59.560 ;
        POLYGON 161.415 59.565 161.425 59.565 161.425 59.560 ;
        RECT 161.425 59.560 164.435 59.565 ;
        POLYGON 164.435 59.635 164.520 59.560 164.435 59.560 ;
        POLYGON 167.915 59.635 167.950 59.635 167.950 59.595 ;
        RECT 167.950 59.615 172.615 59.635 ;
        POLYGON 172.615 59.665 172.650 59.615 172.615 59.615 ;
        POLYGON 180.050 59.665 180.075 59.665 180.075 59.620 ;
        RECT 180.075 59.615 194.510 59.665 ;
        RECT 167.950 59.595 172.650 59.615 ;
        POLYGON 167.950 59.595 167.975 59.595 167.975 59.560 ;
        RECT 167.975 59.585 172.650 59.595 ;
        POLYGON 172.650 59.615 172.665 59.585 172.650 59.585 ;
        POLYGON 180.075 59.615 180.085 59.615 180.085 59.605 ;
        RECT 180.085 59.605 194.510 59.615 ;
        POLYGON 180.085 59.605 180.090 59.605 180.090 59.590 ;
        RECT 180.090 59.585 194.510 59.605 ;
        RECT 167.975 59.560 172.665 59.585 ;
        RECT 152.415 59.550 158.170 59.560 ;
        POLYGON 158.170 59.560 158.210 59.550 158.170 59.550 ;
        POLYGON 161.425 59.560 161.440 59.560 161.440 59.550 ;
        RECT 161.440 59.550 164.520 59.560 ;
        POLYGON 152.325 59.550 152.325 59.515 152.200 59.515 ;
        RECT 152.325 59.545 158.210 59.550 ;
        POLYGON 158.210 59.550 158.240 59.545 158.210 59.545 ;
        POLYGON 161.440 59.550 161.450 59.550 161.450 59.545 ;
        RECT 161.450 59.545 164.520 59.550 ;
        RECT 152.325 59.515 158.240 59.545 ;
        POLYGON 152.200 59.515 152.200 59.500 152.150 59.500 ;
        RECT 152.200 59.500 158.240 59.515 ;
        POLYGON 152.150 59.500 152.150 59.475 152.085 59.475 ;
        RECT 152.150 59.490 158.240 59.500 ;
        POLYGON 158.240 59.545 158.410 59.490 158.240 59.490 ;
        POLYGON 161.450 59.545 161.545 59.545 161.545 59.490 ;
        RECT 161.545 59.490 164.520 59.545 ;
        RECT 152.150 59.475 158.410 59.490 ;
        RECT 146.845 59.470 149.425 59.475 ;
        POLYGON 149.425 59.475 149.430 59.475 149.425 59.470 ;
        POLYGON 152.085 59.475 152.085 59.470 152.070 59.470 ;
        RECT 152.085 59.470 158.410 59.475 ;
        RECT 146.845 59.375 149.245 59.470 ;
        POLYGON 145.590 59.375 145.625 59.235 145.590 59.235 ;
        RECT 117.445 59.090 145.625 59.235 ;
        POLYGON 146.670 59.375 146.670 59.220 146.515 59.220 ;
        RECT 146.670 59.360 149.245 59.375 ;
        POLYGON 149.245 59.470 149.425 59.470 149.245 59.360 ;
        POLYGON 152.070 59.470 152.070 59.430 151.945 59.430 ;
        RECT 152.070 59.430 158.410 59.470 ;
        POLYGON 151.945 59.430 151.945 59.425 151.935 59.425 ;
        RECT 151.945 59.425 158.410 59.430 ;
        POLYGON 151.935 59.425 151.935 59.420 151.910 59.420 ;
        RECT 151.935 59.420 158.410 59.425 ;
        POLYGON 151.910 59.420 151.910 59.380 151.805 59.380 ;
        RECT 151.910 59.415 158.410 59.420 ;
        POLYGON 158.410 59.490 158.660 59.415 158.410 59.415 ;
        POLYGON 161.545 59.490 161.555 59.490 161.555 59.485 ;
        RECT 161.555 59.485 164.520 59.490 ;
        POLYGON 161.555 59.485 161.565 59.485 161.565 59.475 ;
        RECT 161.565 59.475 164.520 59.485 ;
        POLYGON 161.565 59.475 161.585 59.475 161.585 59.465 ;
        RECT 161.585 59.465 164.520 59.475 ;
        POLYGON 161.585 59.465 161.660 59.465 161.660 59.415 ;
        RECT 161.660 59.415 164.520 59.465 ;
        RECT 151.910 59.405 158.660 59.415 ;
        POLYGON 158.660 59.415 158.690 59.405 158.660 59.405 ;
        POLYGON 161.660 59.415 161.675 59.415 161.675 59.405 ;
        RECT 161.675 59.405 164.520 59.415 ;
        RECT 151.910 59.380 158.690 59.405 ;
        POLYGON 158.690 59.405 158.770 59.380 158.690 59.380 ;
        POLYGON 161.675 59.405 161.710 59.405 161.710 59.380 ;
        RECT 161.710 59.380 164.520 59.405 ;
        POLYGON 151.805 59.380 151.805 59.360 151.755 59.360 ;
        RECT 151.805 59.375 158.770 59.380 ;
        POLYGON 158.770 59.380 158.785 59.375 158.770 59.375 ;
        POLYGON 161.710 59.380 161.720 59.380 161.720 59.375 ;
        RECT 161.720 59.375 164.520 59.380 ;
        RECT 151.805 59.360 158.785 59.375 ;
        RECT 146.670 59.345 149.220 59.360 ;
        POLYGON 149.220 59.360 149.245 59.360 149.220 59.345 ;
        POLYGON 151.755 59.360 151.755 59.345 151.715 59.345 ;
        RECT 151.755 59.345 158.785 59.360 ;
        RECT 146.670 59.255 149.090 59.345 ;
        POLYGON 149.090 59.345 149.220 59.345 149.090 59.255 ;
        POLYGON 151.715 59.345 151.715 59.340 151.700 59.340 ;
        RECT 151.715 59.340 158.785 59.345 ;
        POLYGON 151.700 59.340 151.700 59.330 151.675 59.330 ;
        RECT 151.700 59.330 158.785 59.340 ;
        POLYGON 158.785 59.375 158.915 59.330 158.785 59.330 ;
        POLYGON 161.720 59.375 161.790 59.375 161.790 59.330 ;
        RECT 161.790 59.330 164.520 59.375 ;
        POLYGON 151.675 59.330 151.675 59.255 151.500 59.255 ;
        RECT 151.675 59.290 158.915 59.330 ;
        POLYGON 158.915 59.330 159.025 59.290 158.915 59.290 ;
        POLYGON 161.790 59.330 161.850 59.330 161.850 59.290 ;
        RECT 161.850 59.305 164.520 59.330 ;
        POLYGON 164.520 59.560 164.795 59.305 164.520 59.305 ;
        POLYGON 167.975 59.560 168.030 59.560 168.030 59.495 ;
        RECT 168.030 59.495 172.665 59.560 ;
        POLYGON 168.030 59.495 168.050 59.495 168.050 59.470 ;
        RECT 168.050 59.470 172.665 59.495 ;
        POLYGON 168.050 59.470 168.180 59.470 168.180 59.305 ;
        RECT 168.180 59.390 172.665 59.470 ;
        POLYGON 172.665 59.585 172.790 59.390 172.665 59.390 ;
        POLYGON 180.090 59.585 180.185 59.585 180.185 59.395 ;
        RECT 180.185 59.390 194.510 59.585 ;
        RECT 168.180 59.305 172.790 59.390 ;
        RECT 161.850 59.290 164.795 59.305 ;
        RECT 151.675 59.255 159.025 59.290 ;
        RECT 146.670 59.220 148.940 59.255 ;
        POLYGON 145.625 59.220 145.660 59.090 145.625 59.090 ;
        RECT 117.445 59.000 145.660 59.090 ;
        POLYGON 146.515 59.220 146.515 59.080 146.380 59.080 ;
        RECT 146.515 59.155 148.940 59.220 ;
        POLYGON 148.940 59.255 149.090 59.255 148.940 59.155 ;
        POLYGON 151.500 59.255 151.500 59.240 151.465 59.240 ;
        RECT 151.500 59.240 159.025 59.255 ;
        POLYGON 151.460 59.240 151.460 59.235 151.445 59.235 ;
        RECT 151.460 59.235 159.025 59.240 ;
        POLYGON 151.445 59.235 151.445 59.155 151.275 59.155 ;
        RECT 151.445 59.230 159.025 59.235 ;
        POLYGON 159.025 59.290 159.180 59.230 159.025 59.230 ;
        POLYGON 161.850 59.290 161.885 59.290 161.885 59.270 ;
        RECT 161.885 59.270 164.795 59.290 ;
        POLYGON 164.795 59.305 164.830 59.270 164.795 59.270 ;
        POLYGON 168.180 59.305 168.205 59.305 168.205 59.275 ;
        RECT 168.205 59.275 172.790 59.305 ;
        POLYGON 168.205 59.275 168.210 59.275 168.210 59.270 ;
        RECT 168.210 59.270 172.790 59.275 ;
        POLYGON 161.890 59.270 161.925 59.270 161.925 59.245 ;
        RECT 161.925 59.245 164.830 59.270 ;
        POLYGON 161.925 59.245 161.945 59.245 161.945 59.230 ;
        RECT 161.945 59.230 164.830 59.245 ;
        RECT 151.445 59.225 159.180 59.230 ;
        POLYGON 159.180 59.230 159.200 59.225 159.180 59.225 ;
        POLYGON 161.945 59.230 161.950 59.230 161.950 59.225 ;
        RECT 161.950 59.225 164.830 59.230 ;
        RECT 151.445 59.195 159.200 59.225 ;
        POLYGON 159.200 59.225 159.275 59.195 159.200 59.195 ;
        POLYGON 161.950 59.225 161.995 59.225 161.995 59.195 ;
        RECT 161.995 59.195 164.830 59.225 ;
        RECT 151.445 59.155 159.275 59.195 ;
        RECT 146.515 59.150 148.935 59.155 ;
        POLYGON 148.935 59.155 148.940 59.155 148.935 59.150 ;
        POLYGON 151.275 59.155 151.275 59.150 151.265 59.150 ;
        RECT 151.275 59.150 159.275 59.155 ;
        RECT 146.515 59.080 148.800 59.150 ;
        POLYGON 117.390 58.975 117.390 58.280 117.340 58.280 ;
        RECT 117.390 58.970 145.660 59.000 ;
        POLYGON 145.660 59.080 145.690 58.970 145.660 58.970 ;
        RECT 117.390 58.945 145.690 58.970 ;
        POLYGON 146.380 59.080 146.380 58.965 146.270 58.965 ;
        RECT 146.380 59.055 148.800 59.080 ;
        POLYGON 148.800 59.150 148.930 59.150 148.800 59.055 ;
        POLYGON 151.265 59.150 151.265 59.135 151.235 59.135 ;
        RECT 151.265 59.135 159.275 59.150 ;
        POLYGON 151.230 59.135 151.230 59.125 151.220 59.125 ;
        RECT 151.230 59.125 159.275 59.135 ;
        POLYGON 151.220 59.125 151.220 59.055 151.085 59.055 ;
        RECT 151.220 59.120 159.275 59.125 ;
        POLYGON 159.275 59.195 159.445 59.120 159.275 59.120 ;
        POLYGON 161.995 59.195 162.025 59.195 162.025 59.175 ;
        RECT 162.025 59.175 164.830 59.195 ;
        POLYGON 162.025 59.175 162.065 59.175 162.065 59.150 ;
        RECT 162.065 59.150 164.830 59.175 ;
        POLYGON 162.065 59.150 162.105 59.150 162.105 59.120 ;
        RECT 162.105 59.120 164.830 59.150 ;
        RECT 151.220 59.090 159.445 59.120 ;
        POLYGON 159.445 59.120 159.515 59.090 159.445 59.090 ;
        POLYGON 162.105 59.120 162.150 59.120 162.150 59.090 ;
        RECT 162.150 59.090 164.830 59.120 ;
        RECT 151.220 59.055 159.515 59.090 ;
        RECT 146.380 59.025 148.760 59.055 ;
        POLYGON 148.760 59.055 148.800 59.055 148.760 59.025 ;
        POLYGON 151.085 59.055 151.085 59.025 151.025 59.025 ;
        RECT 151.085 59.025 159.515 59.055 ;
        RECT 146.380 58.965 148.645 59.025 ;
        POLYGON 145.690 58.965 145.695 58.945 145.690 58.945 ;
        RECT 117.390 58.865 145.695 58.945 ;
        POLYGON 146.270 58.965 146.270 58.945 146.250 58.945 ;
        RECT 146.270 58.945 148.645 58.965 ;
        RECT 146.250 58.940 148.645 58.945 ;
        POLYGON 148.645 59.025 148.760 59.025 148.645 58.940 ;
        POLYGON 151.025 59.025 151.025 59.010 150.995 59.010 ;
        RECT 151.025 59.010 159.515 59.025 ;
        POLYGON 150.995 59.010 150.995 59.000 150.980 59.000 ;
        RECT 150.995 59.005 159.515 59.010 ;
        POLYGON 159.515 59.090 159.695 59.005 159.515 59.005 ;
        POLYGON 162.150 59.090 162.210 59.090 162.210 59.050 ;
        RECT 162.210 59.060 164.830 59.090 ;
        POLYGON 164.830 59.270 165.045 59.060 164.830 59.060 ;
        POLYGON 168.210 59.270 168.240 59.270 168.240 59.240 ;
        RECT 168.240 59.240 172.790 59.270 ;
        POLYGON 168.240 59.240 168.325 59.240 168.325 59.130 ;
        RECT 168.325 59.195 172.790 59.240 ;
        POLYGON 172.790 59.390 172.905 59.195 172.790 59.195 ;
        POLYGON 180.185 59.390 180.280 59.390 180.280 59.200 ;
        RECT 180.280 59.195 194.510 59.390 ;
        RECT 168.325 59.130 172.905 59.195 ;
        POLYGON 168.325 59.130 168.365 59.130 168.365 59.075 ;
        RECT 168.365 59.075 172.905 59.130 ;
        POLYGON 168.365 59.075 168.375 59.075 168.375 59.060 ;
        RECT 168.375 59.060 172.905 59.075 ;
        RECT 162.210 59.050 165.045 59.060 ;
        POLYGON 162.210 59.050 162.275 59.050 162.275 59.005 ;
        RECT 162.275 59.020 165.045 59.050 ;
        POLYGON 165.045 59.060 165.090 59.020 165.045 59.020 ;
        POLYGON 168.375 59.060 168.405 59.060 168.405 59.020 ;
        RECT 168.405 59.020 172.905 59.060 ;
        RECT 162.275 59.005 165.090 59.020 ;
        RECT 150.995 59.000 159.700 59.005 ;
        POLYGON 150.980 59.000 150.980 58.940 150.860 58.940 ;
        RECT 150.980 58.940 159.700 59.000 ;
        POLYGON 145.695 58.940 145.715 58.865 145.695 58.865 ;
        POLYGON 146.250 58.940 146.250 58.865 146.180 58.865 ;
        RECT 146.250 58.865 148.455 58.940 ;
        RECT 117.390 58.845 145.715 58.865 ;
        POLYGON 146.180 58.865 146.180 58.850 146.170 58.850 ;
        RECT 146.180 58.850 148.455 58.865 ;
        POLYGON 145.715 58.850 145.720 58.845 145.715 58.845 ;
        POLYGON 146.170 58.850 146.170 58.845 146.165 58.845 ;
        RECT 146.170 58.845 148.455 58.850 ;
        RECT 117.390 58.800 145.720 58.845 ;
        POLYGON 145.720 58.845 145.730 58.800 145.720 58.800 ;
        RECT 117.390 58.740 145.730 58.800 ;
        POLYGON 146.165 58.845 146.165 58.790 146.115 58.790 ;
        RECT 146.165 58.795 148.455 58.845 ;
        POLYGON 148.455 58.940 148.645 58.940 148.455 58.795 ;
        POLYGON 150.860 58.940 150.860 58.795 150.620 58.795 ;
        RECT 150.860 58.890 159.700 58.940 ;
        POLYGON 159.700 59.005 159.930 58.890 159.700 58.890 ;
        POLYGON 162.275 59.005 162.430 59.005 162.430 58.890 ;
        RECT 162.430 58.965 165.090 59.005 ;
        POLYGON 165.090 59.020 165.140 58.965 165.090 58.965 ;
        POLYGON 168.405 59.020 168.440 59.020 168.440 58.970 ;
        RECT 168.440 58.965 172.905 59.020 ;
        RECT 162.430 58.890 165.140 58.965 ;
        RECT 150.860 58.885 154.975 58.890 ;
        POLYGON 154.975 58.890 155.350 58.890 154.975 58.885 ;
        POLYGON 155.540 58.890 155.660 58.890 155.660 58.885 ;
        RECT 155.660 58.885 159.930 58.890 ;
        RECT 150.860 58.880 154.925 58.885 ;
        POLYGON 154.925 58.885 154.975 58.885 154.925 58.880 ;
        POLYGON 155.660 58.885 155.780 58.885 155.780 58.880 ;
        RECT 155.780 58.880 159.930 58.885 ;
        RECT 150.860 58.875 154.850 58.880 ;
        POLYGON 154.850 58.880 154.915 58.880 154.850 58.875 ;
        POLYGON 155.780 58.880 155.905 58.880 155.905 58.875 ;
        RECT 155.905 58.875 159.930 58.880 ;
        RECT 150.860 58.860 154.630 58.875 ;
        POLYGON 154.630 58.875 154.850 58.875 154.630 58.860 ;
        POLYGON 155.920 58.875 155.945 58.875 155.945 58.870 ;
        RECT 155.945 58.870 159.930 58.875 ;
        POLYGON 155.995 58.870 156.105 58.870 156.105 58.865 ;
        RECT 156.105 58.865 159.930 58.870 ;
        POLYGON 156.105 58.865 156.145 58.865 156.145 58.860 ;
        RECT 156.145 58.860 159.930 58.865 ;
        RECT 150.860 58.845 154.425 58.860 ;
        POLYGON 154.425 58.860 154.625 58.860 154.425 58.845 ;
        POLYGON 156.145 58.860 156.265 58.860 156.265 58.845 ;
        RECT 156.265 58.845 159.930 58.860 ;
        RECT 150.860 58.825 154.280 58.845 ;
        POLYGON 154.280 58.845 154.410 58.845 154.280 58.825 ;
        POLYGON 156.265 58.845 156.385 58.845 156.385 58.830 ;
        RECT 156.385 58.830 159.930 58.845 ;
        POLYGON 156.410 58.830 156.445 58.830 156.445 58.825 ;
        RECT 156.445 58.825 159.930 58.830 ;
        RECT 150.860 58.815 154.185 58.825 ;
        POLYGON 154.185 58.825 154.280 58.825 154.185 58.815 ;
        POLYGON 156.445 58.825 156.525 58.825 156.525 58.815 ;
        RECT 156.525 58.815 159.930 58.825 ;
        RECT 150.860 58.795 153.935 58.815 ;
        RECT 146.165 58.790 148.435 58.795 ;
        POLYGON 145.730 58.790 145.745 58.740 145.730 58.740 ;
        RECT 117.390 58.680 145.745 58.740 ;
        POLYGON 146.115 58.790 146.115 58.730 146.060 58.730 ;
        RECT 146.115 58.780 148.435 58.790 ;
        POLYGON 148.435 58.795 148.455 58.795 148.435 58.780 ;
        POLYGON 150.620 58.795 150.620 58.780 150.595 58.780 ;
        RECT 150.620 58.780 153.935 58.795 ;
        POLYGON 153.935 58.815 154.180 58.815 153.935 58.780 ;
        POLYGON 156.525 58.815 156.565 58.815 156.565 58.810 ;
        RECT 156.565 58.810 159.930 58.815 ;
        POLYGON 156.570 58.810 156.670 58.810 156.670 58.800 ;
        RECT 156.670 58.800 159.930 58.810 ;
        POLYGON 156.670 58.800 156.790 58.800 156.790 58.780 ;
        RECT 156.790 58.785 159.930 58.800 ;
        POLYGON 159.930 58.890 160.130 58.785 159.930 58.785 ;
        POLYGON 162.430 58.890 162.440 58.890 162.440 58.885 ;
        RECT 162.440 58.885 165.140 58.890 ;
        POLYGON 162.440 58.885 162.460 58.885 162.460 58.870 ;
        RECT 162.460 58.870 165.140 58.885 ;
        POLYGON 162.460 58.870 162.525 58.870 162.525 58.820 ;
        RECT 162.525 58.820 165.140 58.870 ;
        POLYGON 162.525 58.820 162.570 58.820 162.570 58.785 ;
        RECT 162.570 58.785 165.140 58.820 ;
        RECT 156.790 58.780 160.130 58.785 ;
        RECT 146.115 58.745 148.390 58.780 ;
        POLYGON 148.390 58.780 148.435 58.780 148.390 58.745 ;
        POLYGON 150.595 58.780 150.595 58.765 150.570 58.765 ;
        RECT 150.595 58.770 153.850 58.780 ;
        POLYGON 153.850 58.780 153.930 58.780 153.850 58.770 ;
        POLYGON 156.790 58.780 156.825 58.780 156.825 58.775 ;
        RECT 156.825 58.775 160.130 58.780 ;
        POLYGON 156.830 58.775 156.855 58.775 156.855 58.770 ;
        RECT 156.855 58.770 160.130 58.775 ;
        RECT 150.595 58.765 153.725 58.770 ;
        POLYGON 150.565 58.765 150.565 58.750 150.540 58.750 ;
        RECT 150.565 58.750 153.725 58.765 ;
        POLYGON 150.540 58.750 150.540 58.745 150.530 58.745 ;
        RECT 150.540 58.745 153.725 58.750 ;
        POLYGON 153.725 58.770 153.850 58.770 153.725 58.745 ;
        POLYGON 156.855 58.770 156.905 58.770 156.905 58.760 ;
        RECT 156.905 58.760 160.130 58.770 ;
        POLYGON 156.905 58.760 156.950 58.760 156.950 58.755 ;
        RECT 156.950 58.755 160.130 58.760 ;
        POLYGON 156.950 58.755 157.000 58.755 157.000 58.745 ;
        RECT 157.000 58.750 160.130 58.755 ;
        POLYGON 160.130 58.785 160.185 58.750 160.130 58.750 ;
        POLYGON 162.570 58.785 162.610 58.785 162.610 58.760 ;
        RECT 162.610 58.760 165.140 58.785 ;
        POLYGON 162.610 58.760 162.620 58.760 162.620 58.750 ;
        RECT 162.620 58.750 165.140 58.760 ;
        RECT 157.000 58.745 160.185 58.750 ;
        RECT 146.115 58.730 148.360 58.745 ;
        POLYGON 145.745 58.730 145.760 58.680 145.745 58.680 ;
        POLYGON 146.060 58.730 146.060 58.680 146.015 58.680 ;
        RECT 146.060 58.725 148.360 58.730 ;
        POLYGON 148.360 58.745 148.390 58.745 148.360 58.725 ;
        POLYGON 150.530 58.745 150.530 58.725 150.495 58.725 ;
        RECT 150.530 58.725 153.435 58.745 ;
        RECT 146.060 58.680 148.130 58.725 ;
        RECT 117.390 58.655 145.760 58.680 ;
        POLYGON 145.760 58.680 145.765 58.655 145.760 58.655 ;
        POLYGON 146.015 58.680 146.015 58.655 145.995 58.655 ;
        RECT 146.015 58.655 148.130 58.680 ;
        RECT 117.390 58.575 145.765 58.655 ;
        POLYGON 145.765 58.655 145.785 58.575 145.765 58.575 ;
        POLYGON 145.995 58.655 145.995 58.615 145.960 58.615 ;
        RECT 145.995 58.615 148.130 58.655 ;
        RECT 117.390 58.470 145.785 58.575 ;
        POLYGON 145.960 58.615 145.960 58.570 145.925 58.570 ;
        RECT 145.960 58.570 148.130 58.615 ;
        POLYGON 145.785 58.570 145.810 58.470 145.785 58.470 ;
        POLYGON 145.925 58.570 145.925 58.490 145.855 58.490 ;
        RECT 145.925 58.530 148.130 58.570 ;
        POLYGON 148.130 58.725 148.360 58.725 148.130 58.530 ;
        POLYGON 150.495 58.725 150.495 58.715 150.480 58.715 ;
        RECT 150.495 58.715 153.435 58.725 ;
        POLYGON 150.480 58.715 150.480 58.530 150.195 58.530 ;
        RECT 150.480 58.685 153.435 58.715 ;
        POLYGON 153.435 58.745 153.720 58.745 153.435 58.685 ;
        POLYGON 157.000 58.745 157.135 58.745 157.135 58.720 ;
        RECT 157.135 58.720 160.185 58.745 ;
        POLYGON 157.140 58.720 157.235 58.720 157.235 58.700 ;
        RECT 157.235 58.700 160.185 58.720 ;
        POLYGON 157.235 58.700 157.265 58.700 157.265 58.690 ;
        RECT 157.265 58.690 160.185 58.700 ;
        POLYGON 157.265 58.690 157.285 58.690 157.285 58.685 ;
        RECT 157.285 58.685 160.185 58.690 ;
        RECT 150.480 58.665 153.325 58.685 ;
        POLYGON 153.325 58.685 153.435 58.685 153.325 58.665 ;
        POLYGON 157.285 58.685 157.370 58.685 157.370 58.665 ;
        RECT 157.370 58.665 160.185 58.685 ;
        RECT 150.480 58.630 153.180 58.665 ;
        POLYGON 153.180 58.665 153.320 58.665 153.180 58.630 ;
        POLYGON 157.370 58.665 157.395 58.665 157.395 58.660 ;
        RECT 157.395 58.660 160.185 58.665 ;
        POLYGON 157.395 58.660 157.515 58.660 157.515 58.635 ;
        RECT 157.515 58.635 160.185 58.660 ;
        POLYGON 160.185 58.750 160.390 58.635 160.185 58.635 ;
        POLYGON 162.620 58.750 162.765 58.750 162.765 58.635 ;
        RECT 162.765 58.635 165.140 58.750 ;
        POLYGON 157.515 58.635 157.530 58.635 157.530 58.630 ;
        RECT 157.530 58.630 160.390 58.635 ;
        RECT 150.480 58.565 152.950 58.630 ;
        POLYGON 152.950 58.630 153.180 58.630 152.950 58.565 ;
        POLYGON 157.530 58.630 157.695 58.630 157.695 58.585 ;
        RECT 157.695 58.620 160.390 58.630 ;
        POLYGON 160.390 58.635 160.415 58.620 160.390 58.620 ;
        POLYGON 162.765 58.635 162.780 58.635 162.780 58.620 ;
        RECT 162.780 58.620 165.140 58.635 ;
        RECT 157.695 58.585 160.415 58.620 ;
        POLYGON 157.700 58.585 157.770 58.585 157.770 58.565 ;
        RECT 157.770 58.570 160.415 58.585 ;
        POLYGON 160.415 58.620 160.495 58.570 160.415 58.570 ;
        POLYGON 162.780 58.620 162.790 58.620 162.790 58.615 ;
        RECT 162.790 58.615 165.140 58.620 ;
        POLYGON 165.140 58.965 165.475 58.615 165.140 58.615 ;
        POLYGON 168.440 58.965 168.510 58.965 168.510 58.875 ;
        RECT 168.510 58.875 172.905 58.965 ;
        POLYGON 168.510 58.875 168.555 58.875 168.555 58.815 ;
        RECT 168.555 58.815 172.905 58.875 ;
        POLYGON 168.555 58.815 168.640 58.815 168.640 58.695 ;
        RECT 168.640 58.695 172.905 58.815 ;
        POLYGON 168.640 58.695 168.700 58.695 168.700 58.615 ;
        POLYGON 162.790 58.615 162.825 58.615 162.825 58.585 ;
        RECT 162.825 58.585 165.475 58.615 ;
        RECT 168.700 58.610 172.905 58.695 ;
        POLYGON 162.825 58.585 162.845 58.585 162.845 58.570 ;
        RECT 162.845 58.570 165.475 58.585 ;
        RECT 157.770 58.565 160.495 58.570 ;
        RECT 150.480 58.555 152.900 58.565 ;
        POLYGON 152.900 58.565 152.950 58.565 152.900 58.555 ;
        POLYGON 157.770 58.565 157.790 58.565 157.790 58.560 ;
        RECT 157.790 58.560 160.495 58.565 ;
        POLYGON 157.790 58.560 157.805 58.560 157.805 58.555 ;
        RECT 157.805 58.555 160.495 58.560 ;
        RECT 150.480 58.530 152.655 58.555 ;
        RECT 145.925 58.495 148.085 58.530 ;
        POLYGON 148.085 58.530 148.130 58.530 148.085 58.495 ;
        POLYGON 150.195 58.530 150.195 58.495 150.145 58.495 ;
        RECT 150.195 58.495 152.655 58.530 ;
        RECT 145.925 58.490 147.995 58.495 ;
        RECT 117.390 58.440 145.810 58.470 ;
        POLYGON 145.855 58.490 145.855 58.455 145.825 58.455 ;
        RECT 145.855 58.455 147.995 58.490 ;
        POLYGON 145.825 58.455 145.825 58.450 145.820 58.450 ;
        RECT 145.825 58.450 147.995 58.455 ;
        POLYGON 145.810 58.450 145.815 58.440 145.810 58.440 ;
        POLYGON 145.820 58.450 145.820 58.440 145.815 58.440 ;
        RECT 145.820 58.440 147.995 58.450 ;
        RECT 117.390 58.415 147.995 58.440 ;
        POLYGON 147.995 58.495 148.085 58.495 147.995 58.415 ;
        POLYGON 150.145 58.495 150.145 58.490 150.135 58.490 ;
        RECT 150.145 58.490 152.655 58.495 ;
        POLYGON 150.135 58.490 150.135 58.460 150.090 58.460 ;
        RECT 150.135 58.485 152.655 58.490 ;
        POLYGON 152.655 58.555 152.900 58.555 152.655 58.485 ;
        POLYGON 157.805 58.555 158.050 58.555 158.050 58.485 ;
        RECT 158.050 58.485 160.495 58.555 ;
        RECT 150.135 58.460 152.485 58.485 ;
        POLYGON 150.090 58.460 150.090 58.415 150.030 58.415 ;
        RECT 150.090 58.425 152.485 58.460 ;
        POLYGON 152.485 58.485 152.655 58.485 152.485 58.425 ;
        POLYGON 158.050 58.485 158.070 58.485 158.070 58.480 ;
        RECT 158.070 58.480 160.495 58.485 ;
        POLYGON 158.070 58.480 158.125 58.480 158.125 58.460 ;
        RECT 158.125 58.470 160.495 58.480 ;
        POLYGON 160.495 58.570 160.660 58.470 160.495 58.470 ;
        POLYGON 162.845 58.570 162.880 58.570 162.880 58.545 ;
        RECT 162.880 58.545 165.475 58.570 ;
        POLYGON 162.880 58.545 162.935 58.545 162.935 58.500 ;
        RECT 162.935 58.500 165.475 58.545 ;
        POLYGON 162.935 58.500 162.970 58.500 162.970 58.470 ;
        RECT 162.970 58.470 165.475 58.500 ;
        RECT 158.125 58.460 160.665 58.470 ;
        POLYGON 158.130 58.460 158.240 58.460 158.240 58.425 ;
        RECT 150.090 58.420 152.460 58.425 ;
        POLYGON 152.460 58.425 152.485 58.425 152.460 58.420 ;
        RECT 158.240 58.420 160.665 58.460 ;
        RECT 150.090 58.415 152.225 58.420 ;
        RECT 117.390 58.280 147.830 58.415 ;
        RECT 117.340 58.270 147.830 58.280 ;
        POLYGON 147.830 58.415 147.995 58.415 147.830 58.270 ;
        POLYGON 150.030 58.415 150.030 58.350 149.940 58.350 ;
        RECT 150.030 58.350 152.225 58.415 ;
        POLYGON 149.940 58.350 149.940 58.315 149.885 58.315 ;
        RECT 149.940 58.340 152.225 58.350 ;
        POLYGON 152.225 58.420 152.460 58.420 152.225 58.340 ;
        POLYGON 158.240 58.420 158.345 58.420 158.345 58.390 ;
        RECT 158.345 58.390 160.665 58.420 ;
        POLYGON 158.345 58.390 158.355 58.390 158.355 58.385 ;
        RECT 158.355 58.385 160.665 58.390 ;
        POLYGON 158.355 58.385 158.470 58.385 158.470 58.340 ;
        RECT 158.470 58.375 160.665 58.385 ;
        POLYGON 160.665 58.470 160.810 58.375 160.665 58.375 ;
        POLYGON 162.970 58.470 163.080 58.470 163.080 58.375 ;
        RECT 163.080 58.375 165.475 58.470 ;
        RECT 158.470 58.345 160.810 58.375 ;
        POLYGON 160.810 58.375 160.860 58.345 160.810 58.345 ;
        POLYGON 163.080 58.375 163.120 58.375 163.120 58.345 ;
        RECT 163.120 58.345 165.475 58.375 ;
        RECT 158.470 58.340 160.860 58.345 ;
        RECT 149.940 58.315 152.155 58.340 ;
        POLYGON 149.885 58.315 149.885 58.270 149.820 58.270 ;
        RECT 149.885 58.310 152.155 58.315 ;
        POLYGON 152.155 58.340 152.225 58.340 152.155 58.310 ;
        POLYGON 158.470 58.340 158.550 58.340 158.550 58.310 ;
        RECT 158.550 58.310 160.860 58.340 ;
        RECT 149.885 58.280 152.075 58.310 ;
        POLYGON 152.075 58.310 152.150 58.310 152.075 58.280 ;
        POLYGON 158.550 58.310 158.615 58.310 158.615 58.285 ;
        RECT 158.615 58.285 160.860 58.310 ;
        POLYGON 158.615 58.285 158.625 58.285 158.625 58.280 ;
        RECT 158.625 58.280 160.860 58.285 ;
        RECT 149.885 58.270 151.985 58.280 ;
        POLYGON 117.340 58.270 117.340 57.990 117.320 57.990 ;
        RECT 117.340 58.265 147.820 58.270 ;
        POLYGON 147.820 58.270 147.830 58.270 147.820 58.265 ;
        POLYGON 149.820 58.270 149.820 58.265 149.815 58.265 ;
        RECT 149.820 58.265 151.985 58.270 ;
        RECT 117.340 58.060 147.605 58.265 ;
        POLYGON 147.605 58.265 147.820 58.265 147.605 58.060 ;
        POLYGON 149.815 58.265 149.815 58.240 149.780 58.240 ;
        RECT 149.815 58.245 151.985 58.265 ;
        POLYGON 151.985 58.280 152.075 58.280 151.985 58.245 ;
        POLYGON 158.625 58.280 158.715 58.280 158.715 58.245 ;
        RECT 158.715 58.245 160.860 58.280 ;
        RECT 149.815 58.240 151.910 58.245 ;
        POLYGON 149.780 58.240 149.780 58.140 149.650 58.140 ;
        RECT 149.780 58.215 151.910 58.240 ;
        POLYGON 151.910 58.245 151.985 58.245 151.910 58.215 ;
        POLYGON 158.715 58.245 158.770 58.245 158.770 58.225 ;
        RECT 158.770 58.225 160.860 58.245 ;
        POLYGON 158.770 58.225 158.790 58.225 158.790 58.215 ;
        RECT 158.790 58.215 160.860 58.225 ;
        RECT 149.780 58.140 151.705 58.215 ;
        POLYGON 149.650 58.140 149.650 58.060 149.550 58.060 ;
        RECT 149.650 58.130 151.705 58.140 ;
        POLYGON 151.705 58.215 151.910 58.215 151.705 58.130 ;
        POLYGON 158.790 58.215 158.825 58.215 158.825 58.200 ;
        RECT 158.825 58.200 160.860 58.215 ;
        POLYGON 158.825 58.200 158.885 58.200 158.885 58.175 ;
        RECT 158.885 58.175 160.860 58.200 ;
        POLYGON 158.885 58.175 158.965 58.175 158.965 58.140 ;
        RECT 158.965 58.155 160.860 58.175 ;
        POLYGON 160.860 58.345 161.130 58.155 160.860 58.155 ;
        POLYGON 163.120 58.345 163.125 58.345 163.125 58.340 ;
        RECT 163.125 58.340 165.475 58.345 ;
        POLYGON 163.125 58.340 163.245 58.340 163.245 58.235 ;
        RECT 163.245 58.250 165.475 58.340 ;
        POLYGON 165.475 58.610 165.790 58.250 165.475 58.250 ;
        POLYGON 168.700 58.610 168.755 58.610 168.755 58.545 ;
        RECT 168.755 58.595 172.905 58.610 ;
        POLYGON 172.905 59.195 173.275 58.595 172.905 58.595 ;
        POLYGON 180.280 59.195 180.420 59.195 180.420 58.915 ;
        RECT 180.420 58.915 194.510 59.195 ;
        POLYGON 180.420 58.915 180.570 58.915 180.570 58.595 ;
        RECT 180.570 58.595 194.510 58.915 ;
        RECT 168.755 58.540 173.275 58.595 ;
        POLYGON 168.755 58.540 168.795 58.540 168.795 58.480 ;
        RECT 168.795 58.480 173.275 58.540 ;
        POLYGON 168.795 58.480 168.840 58.480 168.840 58.410 ;
        RECT 168.840 58.410 173.275 58.480 ;
        POLYGON 168.840 58.410 168.850 58.410 168.850 58.400 ;
        RECT 168.850 58.400 173.275 58.410 ;
        POLYGON 168.850 58.400 168.890 58.400 168.890 58.340 ;
        RECT 168.890 58.375 173.275 58.400 ;
        POLYGON 173.275 58.595 173.390 58.375 173.275 58.375 ;
        POLYGON 180.570 58.595 180.675 58.595 180.675 58.375 ;
        RECT 180.675 58.590 194.510 58.595 ;
        POLYGON 194.510 59.720 194.980 58.590 194.510 58.590 ;
        POLYGON 206.245 59.720 206.245 58.610 206.235 58.610 ;
        RECT 206.245 59.715 222.755 60.005 ;
        POLYGON 222.755 60.005 222.835 60.005 222.755 59.725 ;
        POLYGON 230.750 60.005 230.750 59.995 230.745 59.995 ;
        RECT 230.750 60.000 235.725 60.010 ;
        POLYGON 235.725 60.065 235.765 60.065 235.725 60.005 ;
        POLYGON 239.490 60.065 239.490 60.005 239.440 60.005 ;
        RECT 239.490 60.050 242.440 60.065 ;
        POLYGON 242.440 60.100 242.505 60.100 242.440 60.050 ;
        POLYGON 245.580 60.100 245.580 60.085 245.560 60.085 ;
        RECT 245.580 60.085 255.420 60.100 ;
        POLYGON 245.555 60.085 245.555 60.050 245.490 60.050 ;
        RECT 245.555 60.050 255.420 60.085 ;
        RECT 239.490 60.005 242.385 60.050 ;
        POLYGON 242.385 60.050 242.440 60.050 242.385 60.005 ;
        POLYGON 245.490 60.050 245.490 60.005 245.405 60.005 ;
        RECT 245.490 60.005 255.420 60.050 ;
        RECT 230.750 59.995 235.595 60.000 ;
        POLYGON 230.745 59.995 230.745 59.725 230.640 59.725 ;
        RECT 230.745 59.795 235.595 59.995 ;
        POLYGON 235.595 60.000 235.725 60.000 235.595 59.795 ;
        POLYGON 239.440 60.005 239.440 59.795 239.260 59.795 ;
        RECT 239.440 59.965 242.340 60.005 ;
        POLYGON 242.340 60.005 242.385 60.005 242.340 59.965 ;
        POLYGON 245.405 60.005 245.405 59.995 245.385 59.995 ;
        RECT 245.405 59.995 255.420 60.005 ;
        POLYGON 245.385 59.995 245.385 59.965 245.330 59.965 ;
        RECT 245.385 59.965 255.420 59.995 ;
        RECT 239.440 59.835 242.190 59.965 ;
        POLYGON 242.190 59.965 242.340 59.965 242.190 59.835 ;
        POLYGON 245.330 59.965 245.330 59.940 245.285 59.940 ;
        RECT 245.330 59.940 255.420 59.965 ;
        POLYGON 245.285 59.940 245.285 59.840 245.095 59.840 ;
        RECT 245.285 59.935 255.420 59.940 ;
        POLYGON 255.420 60.100 255.750 59.935 255.420 59.935 ;
        POLYGON 258.845 60.100 258.905 60.100 258.905 60.050 ;
        RECT 258.905 60.050 262.405 60.100 ;
        POLYGON 258.905 60.050 258.960 60.050 258.960 60.005 ;
        RECT 258.960 60.005 262.405 60.050 ;
        POLYGON 262.405 60.190 262.565 60.005 262.405 60.005 ;
        POLYGON 267.235 60.190 267.365 60.190 267.365 60.005 ;
        RECT 267.365 60.170 274.500 60.190 ;
        POLYGON 274.500 60.680 274.785 60.170 274.500 60.170 ;
        POLYGON 287.655 60.680 287.710 60.680 287.710 60.185 ;
        RECT 287.710 60.170 303.120 60.680 ;
        RECT 267.365 60.005 274.785 60.170 ;
        POLYGON 274.785 60.170 274.870 60.005 274.785 60.005 ;
        POLYGON 287.710 60.170 287.730 60.170 287.730 60.005 ;
        POLYGON 258.960 60.005 259.045 60.005 259.045 59.935 ;
        RECT 259.045 59.935 262.565 60.005 ;
        RECT 245.285 59.930 255.750 59.935 ;
        RECT 245.285 59.925 249.890 59.930 ;
        POLYGON 249.890 59.930 250.430 59.930 249.890 59.925 ;
        POLYGON 250.430 59.930 250.550 59.930 250.550 59.925 ;
        RECT 250.550 59.925 255.750 59.930 ;
        RECT 245.285 59.915 249.695 59.925 ;
        POLYGON 249.695 59.925 249.860 59.925 249.695 59.915 ;
        POLYGON 250.550 59.925 250.790 59.925 250.790 59.915 ;
        RECT 250.790 59.920 255.750 59.925 ;
        POLYGON 255.750 59.935 255.775 59.920 255.750 59.920 ;
        POLYGON 259.045 59.935 259.065 59.935 259.065 59.920 ;
        RECT 259.065 59.920 262.565 59.935 ;
        RECT 250.790 59.915 255.775 59.920 ;
        RECT 245.285 59.900 249.380 59.915 ;
        POLYGON 249.380 59.915 249.655 59.915 249.380 59.900 ;
        POLYGON 250.790 59.915 250.910 59.915 250.910 59.910 ;
        RECT 250.910 59.910 255.775 59.915 ;
        POLYGON 250.915 59.910 251.005 59.910 251.005 59.905 ;
        RECT 251.005 59.905 255.775 59.910 ;
        POLYGON 251.005 59.905 251.060 59.905 251.060 59.900 ;
        RECT 251.060 59.900 255.775 59.905 ;
        POLYGON 255.775 59.920 255.815 59.900 255.775 59.900 ;
        POLYGON 259.065 59.920 259.090 59.920 259.090 59.900 ;
        RECT 259.090 59.900 262.565 59.920 ;
        RECT 245.285 59.895 249.290 59.900 ;
        POLYGON 249.290 59.900 249.380 59.900 249.290 59.895 ;
        POLYGON 251.060 59.900 251.115 59.900 251.115 59.895 ;
        RECT 251.115 59.895 255.815 59.900 ;
        RECT 245.285 59.860 248.965 59.895 ;
        POLYGON 248.965 59.895 249.290 59.895 248.965 59.860 ;
        POLYGON 251.115 59.895 251.335 59.895 251.335 59.875 ;
        RECT 251.335 59.875 255.815 59.895 ;
        POLYGON 251.345 59.875 251.415 59.875 251.415 59.865 ;
        RECT 251.415 59.865 255.815 59.875 ;
        POLYGON 251.425 59.865 251.475 59.865 251.475 59.860 ;
        RECT 251.475 59.860 255.815 59.865 ;
        RECT 245.285 59.855 248.940 59.860 ;
        POLYGON 248.940 59.860 248.960 59.860 248.940 59.855 ;
        POLYGON 251.475 59.860 251.525 59.860 251.525 59.855 ;
        RECT 251.525 59.855 255.815 59.860 ;
        RECT 245.285 59.850 248.875 59.855 ;
        POLYGON 248.875 59.855 248.940 59.855 248.875 59.850 ;
        POLYGON 251.525 59.855 251.580 59.855 251.580 59.850 ;
        RECT 251.580 59.850 255.815 59.855 ;
        RECT 245.285 59.840 248.735 59.850 ;
        POLYGON 245.090 59.840 245.090 59.835 245.080 59.835 ;
        RECT 245.090 59.835 248.735 59.840 ;
        POLYGON 248.735 59.850 248.875 59.850 248.735 59.835 ;
        POLYGON 251.605 59.850 251.710 59.850 251.710 59.835 ;
        RECT 251.710 59.835 255.815 59.850 ;
        RECT 239.440 59.810 242.160 59.835 ;
        POLYGON 242.160 59.835 242.190 59.835 242.160 59.810 ;
        POLYGON 245.080 59.835 245.080 59.810 245.035 59.810 ;
        RECT 245.080 59.820 248.660 59.835 ;
        POLYGON 248.660 59.835 248.735 59.835 248.660 59.820 ;
        POLYGON 251.710 59.835 251.820 59.835 251.820 59.820 ;
        RECT 251.820 59.820 255.815 59.835 ;
        RECT 245.080 59.810 248.380 59.820 ;
        RECT 239.440 59.795 242.105 59.810 ;
        RECT 230.745 59.725 235.555 59.795 ;
        POLYGON 235.555 59.795 235.595 59.795 235.555 59.725 ;
        POLYGON 239.260 59.795 239.260 59.725 239.200 59.725 ;
        RECT 239.260 59.760 242.105 59.795 ;
        POLYGON 242.105 59.810 242.160 59.810 242.105 59.760 ;
        POLYGON 245.035 59.810 245.035 59.760 244.945 59.760 ;
        RECT 245.035 59.775 248.380 59.810 ;
        POLYGON 248.380 59.820 248.660 59.820 248.380 59.775 ;
        POLYGON 251.820 59.820 251.860 59.820 251.860 59.815 ;
        RECT 251.860 59.815 255.815 59.820 ;
        POLYGON 251.860 59.815 251.915 59.815 251.915 59.805 ;
        RECT 251.915 59.805 255.815 59.815 ;
        POLYGON 251.925 59.805 252.040 59.805 252.040 59.790 ;
        RECT 252.040 59.790 255.815 59.805 ;
        POLYGON 252.040 59.790 252.090 59.790 252.090 59.780 ;
        RECT 252.090 59.780 255.815 59.790 ;
        POLYGON 252.095 59.780 252.145 59.780 252.145 59.775 ;
        RECT 252.145 59.775 255.815 59.780 ;
        RECT 245.035 59.765 248.315 59.775 ;
        POLYGON 248.315 59.775 248.370 59.775 248.315 59.765 ;
        POLYGON 252.145 59.775 252.195 59.775 252.195 59.765 ;
        RECT 252.195 59.765 255.815 59.775 ;
        RECT 245.035 59.760 248.190 59.765 ;
        RECT 239.260 59.725 242.065 59.760 ;
        POLYGON 242.065 59.760 242.105 59.760 242.065 59.725 ;
        POLYGON 244.945 59.760 244.945 59.745 244.915 59.745 ;
        RECT 244.945 59.745 248.190 59.760 ;
        POLYGON 248.190 59.765 248.295 59.765 248.190 59.745 ;
        POLYGON 252.195 59.765 252.295 59.765 252.295 59.745 ;
        RECT 252.295 59.745 255.815 59.765 ;
        POLYGON 244.915 59.745 244.915 59.740 244.900 59.740 ;
        RECT 244.915 59.740 248.010 59.745 ;
        POLYGON 244.900 59.740 244.900 59.725 244.875 59.725 ;
        RECT 244.900 59.725 248.010 59.740 ;
        RECT 206.245 58.990 222.585 59.715 ;
        POLYGON 222.585 59.715 222.755 59.715 222.585 59.000 ;
        POLYGON 230.640 59.720 230.640 59.370 230.505 59.370 ;
        RECT 230.640 59.370 235.190 59.725 ;
        POLYGON 230.505 59.370 230.505 59.000 230.375 59.000 ;
        RECT 230.505 59.065 235.190 59.370 ;
        POLYGON 235.190 59.725 235.555 59.725 235.190 59.065 ;
        POLYGON 239.200 59.725 239.200 59.635 239.125 59.635 ;
        RECT 239.200 59.635 241.880 59.725 ;
        POLYGON 239.125 59.635 239.125 59.425 238.965 59.425 ;
        RECT 239.125 59.560 241.880 59.635 ;
        POLYGON 241.880 59.725 242.065 59.725 241.880 59.560 ;
        POLYGON 244.875 59.725 244.875 59.650 244.750 59.650 ;
        RECT 244.875 59.705 248.010 59.725 ;
        POLYGON 248.010 59.745 248.190 59.745 248.010 59.705 ;
        POLYGON 252.295 59.745 252.320 59.745 252.320 59.740 ;
        RECT 252.320 59.740 255.815 59.745 ;
        POLYGON 252.325 59.740 252.345 59.740 252.345 59.735 ;
        RECT 252.345 59.735 255.815 59.740 ;
        POLYGON 252.350 59.735 252.390 59.735 252.390 59.725 ;
        RECT 252.390 59.725 255.815 59.735 ;
        POLYGON 255.815 59.900 256.135 59.725 255.815 59.725 ;
        POLYGON 259.090 59.900 259.105 59.900 259.105 59.890 ;
        RECT 259.105 59.890 262.565 59.900 ;
        POLYGON 259.105 59.890 259.130 59.890 259.130 59.875 ;
        RECT 259.130 59.875 262.565 59.890 ;
        POLYGON 259.130 59.875 259.150 59.875 259.150 59.855 ;
        RECT 259.150 59.855 262.565 59.875 ;
        POLYGON 259.150 59.855 259.300 59.855 259.300 59.725 ;
        RECT 259.300 59.775 262.565 59.855 ;
        POLYGON 262.565 60.005 262.770 59.775 262.565 59.775 ;
        POLYGON 267.365 60.005 267.520 60.005 267.520 59.780 ;
        RECT 267.520 59.850 274.870 60.005 ;
        POLYGON 274.870 60.005 274.950 59.850 274.870 59.850 ;
        RECT 287.730 59.995 303.120 60.170 ;
        POLYGON 287.730 59.995 287.745 59.995 287.745 59.860 ;
        RECT 287.745 59.850 303.120 59.995 ;
        RECT 267.520 59.775 274.950 59.850 ;
        RECT 259.300 59.725 262.770 59.775 ;
        POLYGON 262.770 59.775 262.810 59.725 262.770 59.725 ;
        POLYGON 267.520 59.775 267.555 59.775 267.555 59.725 ;
        RECT 267.555 59.730 274.950 59.775 ;
        POLYGON 274.950 59.850 275.010 59.730 274.950 59.730 ;
        RECT 267.555 59.725 275.010 59.730 ;
        POLYGON 287.745 59.850 287.760 59.850 287.760 59.725 ;
        POLYGON 252.390 59.725 252.415 59.725 252.415 59.720 ;
        RECT 252.415 59.720 256.135 59.725 ;
        POLYGON 256.135 59.725 256.145 59.720 256.135 59.720 ;
        POLYGON 259.300 59.725 259.305 59.725 259.305 59.720 ;
        RECT 259.305 59.720 262.810 59.725 ;
        POLYGON 252.415 59.720 252.505 59.720 252.505 59.705 ;
        RECT 252.505 59.705 256.145 59.720 ;
        RECT 244.875 59.685 247.895 59.705 ;
        POLYGON 247.895 59.705 248.010 59.705 247.895 59.685 ;
        POLYGON 252.505 59.705 252.540 59.705 252.540 59.700 ;
        RECT 252.540 59.700 256.145 59.705 ;
        POLYGON 252.545 59.700 252.605 59.700 252.605 59.685 ;
        RECT 252.605 59.690 256.145 59.700 ;
        POLYGON 256.145 59.720 256.200 59.690 256.145 59.690 ;
        POLYGON 259.305 59.720 259.340 59.720 259.340 59.690 ;
        RECT 259.340 59.690 262.810 59.720 ;
        RECT 252.605 59.685 256.200 59.690 ;
        RECT 244.875 59.670 247.840 59.685 ;
        POLYGON 247.840 59.685 247.895 59.685 247.840 59.670 ;
        POLYGON 252.605 59.685 252.630 59.685 252.630 59.680 ;
        RECT 252.630 59.680 256.200 59.685 ;
        POLYGON 252.635 59.680 252.680 59.680 252.680 59.670 ;
        RECT 252.680 59.670 256.200 59.680 ;
        RECT 244.875 59.650 247.665 59.670 ;
        POLYGON 244.750 59.650 244.750 59.560 244.605 59.560 ;
        RECT 244.750 59.635 247.665 59.650 ;
        POLYGON 247.665 59.670 247.840 59.670 247.665 59.635 ;
        POLYGON 252.680 59.670 252.705 59.670 252.705 59.665 ;
        RECT 252.705 59.665 256.200 59.670 ;
        POLYGON 252.705 59.665 252.760 59.665 252.760 59.655 ;
        RECT 252.760 59.655 256.200 59.665 ;
        POLYGON 256.200 59.690 256.255 59.655 256.200 59.655 ;
        POLYGON 259.340 59.690 259.365 59.690 259.365 59.670 ;
        RECT 259.365 59.670 262.810 59.690 ;
        POLYGON 259.370 59.670 259.385 59.670 259.385 59.655 ;
        RECT 259.385 59.655 262.810 59.670 ;
        POLYGON 252.760 59.655 252.835 59.655 252.835 59.635 ;
        RECT 252.835 59.635 256.255 59.655 ;
        RECT 244.750 59.610 247.590 59.635 ;
        POLYGON 247.590 59.635 247.665 59.635 247.590 59.610 ;
        POLYGON 252.835 59.635 252.895 59.635 252.895 59.620 ;
        RECT 252.895 59.620 256.255 59.635 ;
        POLYGON 252.905 59.620 252.940 59.620 252.940 59.610 ;
        RECT 252.940 59.610 256.255 59.620 ;
        RECT 244.750 59.580 247.490 59.610 ;
        POLYGON 247.490 59.610 247.590 59.610 247.490 59.580 ;
        POLYGON 252.940 59.610 252.975 59.610 252.975 59.600 ;
        RECT 252.975 59.600 256.255 59.610 ;
        POLYGON 252.980 59.600 253.060 59.600 253.060 59.580 ;
        RECT 253.060 59.580 256.255 59.600 ;
        RECT 244.750 59.565 247.425 59.580 ;
        POLYGON 247.425 59.580 247.485 59.580 247.425 59.565 ;
        POLYGON 253.060 59.580 253.120 59.580 253.120 59.565 ;
        RECT 253.120 59.565 256.255 59.580 ;
        RECT 244.750 59.560 247.340 59.565 ;
        RECT 239.125 59.425 241.710 59.560 ;
        POLYGON 238.965 59.425 238.965 59.080 238.710 59.080 ;
        RECT 238.965 59.395 241.710 59.425 ;
        POLYGON 241.710 59.560 241.880 59.560 241.710 59.395 ;
        POLYGON 244.605 59.560 244.605 59.525 244.550 59.525 ;
        RECT 244.605 59.540 247.340 59.560 ;
        POLYGON 247.340 59.565 247.425 59.565 247.340 59.540 ;
        POLYGON 253.120 59.565 253.165 59.565 253.165 59.555 ;
        RECT 253.165 59.555 256.255 59.565 ;
        POLYGON 253.165 59.555 253.225 59.555 253.225 59.540 ;
        RECT 253.225 59.540 256.255 59.555 ;
        RECT 244.605 59.525 247.245 59.540 ;
        POLYGON 244.550 59.525 244.550 59.460 244.440 59.460 ;
        RECT 244.550 59.515 247.245 59.525 ;
        POLYGON 247.245 59.540 247.335 59.540 247.245 59.515 ;
        POLYGON 253.225 59.540 253.250 59.540 253.250 59.535 ;
        RECT 253.250 59.535 256.255 59.540 ;
        POLYGON 253.250 59.535 253.310 59.535 253.310 59.515 ;
        RECT 253.310 59.515 256.255 59.535 ;
        RECT 244.550 59.500 247.195 59.515 ;
        POLYGON 247.195 59.515 247.245 59.515 247.195 59.500 ;
        POLYGON 253.310 59.515 253.355 59.515 253.355 59.500 ;
        RECT 253.355 59.500 256.255 59.515 ;
        RECT 244.550 59.490 247.165 59.500 ;
        POLYGON 247.165 59.500 247.195 59.500 247.165 59.490 ;
        POLYGON 253.355 59.500 253.395 59.500 253.395 59.490 ;
        RECT 253.395 59.490 256.255 59.500 ;
        POLYGON 256.255 59.655 256.535 59.490 256.255 59.490 ;
        POLYGON 259.385 59.655 259.475 59.655 259.475 59.575 ;
        RECT 259.475 59.575 262.810 59.655 ;
        POLYGON 259.475 59.575 259.495 59.575 259.495 59.555 ;
        RECT 259.495 59.570 262.810 59.575 ;
        POLYGON 262.810 59.725 262.950 59.570 262.810 59.570 ;
        POLYGON 267.555 59.725 267.575 59.725 267.575 59.700 ;
        RECT 267.575 59.700 275.010 59.725 ;
        POLYGON 267.575 59.700 267.645 59.700 267.645 59.605 ;
        RECT 267.645 59.605 275.010 59.700 ;
        POLYGON 267.645 59.605 267.665 59.605 267.665 59.570 ;
        RECT 267.665 59.570 275.010 59.605 ;
        RECT 259.495 59.555 262.950 59.570 ;
        POLYGON 259.495 59.555 259.565 59.555 259.565 59.490 ;
        RECT 259.565 59.490 262.950 59.555 ;
        POLYGON 262.950 59.570 263.020 59.490 262.950 59.490 ;
        POLYGON 267.665 59.570 267.710 59.570 267.710 59.495 ;
        RECT 267.710 59.565 275.010 59.570 ;
        POLYGON 275.010 59.725 275.095 59.565 275.010 59.565 ;
        RECT 287.760 59.720 303.120 59.850 ;
        POLYGON 287.760 59.720 287.775 59.720 287.775 59.580 ;
        RECT 287.775 59.565 303.120 59.720 ;
        RECT 267.710 59.490 275.095 59.565 ;
        RECT 244.550 59.465 247.085 59.490 ;
        POLYGON 247.085 59.490 247.165 59.490 247.085 59.465 ;
        POLYGON 253.395 59.490 253.415 59.490 253.415 59.485 ;
        RECT 253.415 59.485 256.535 59.490 ;
        POLYGON 256.535 59.490 256.540 59.485 256.535 59.485 ;
        POLYGON 259.565 59.490 259.570 59.490 259.570 59.485 ;
        RECT 259.570 59.485 263.020 59.490 ;
        POLYGON 253.415 59.485 253.420 59.485 253.420 59.480 ;
        RECT 253.420 59.480 256.540 59.485 ;
        POLYGON 253.420 59.480 253.470 59.480 253.470 59.465 ;
        RECT 253.470 59.465 256.540 59.480 ;
        POLYGON 256.540 59.485 256.570 59.465 256.540 59.465 ;
        POLYGON 259.570 59.485 259.595 59.485 259.595 59.465 ;
        RECT 259.595 59.465 263.020 59.485 ;
        RECT 244.550 59.460 247.010 59.465 ;
        POLYGON 244.435 59.460 244.435 59.395 244.330 59.395 ;
        RECT 244.435 59.435 247.010 59.460 ;
        POLYGON 247.010 59.465 247.085 59.465 247.010 59.435 ;
        POLYGON 253.470 59.465 253.580 59.465 253.580 59.435 ;
        RECT 253.580 59.435 256.570 59.465 ;
        RECT 244.435 59.425 246.970 59.435 ;
        POLYGON 246.970 59.435 247.010 59.435 246.970 59.425 ;
        POLYGON 253.580 59.435 253.605 59.435 253.605 59.425 ;
        RECT 253.605 59.425 256.570 59.435 ;
        RECT 244.435 59.410 246.920 59.425 ;
        POLYGON 246.920 59.425 246.970 59.425 246.920 59.410 ;
        POLYGON 253.605 59.425 253.650 59.425 253.650 59.410 ;
        RECT 253.650 59.410 256.570 59.425 ;
        RECT 244.435 59.395 246.820 59.410 ;
        RECT 238.965 59.350 241.670 59.395 ;
        POLYGON 241.670 59.395 241.710 59.395 241.670 59.350 ;
        POLYGON 244.330 59.395 244.330 59.350 244.260 59.350 ;
        RECT 244.330 59.370 246.820 59.395 ;
        POLYGON 246.820 59.410 246.920 59.410 246.820 59.370 ;
        POLYGON 253.650 59.410 253.665 59.410 253.665 59.405 ;
        RECT 253.665 59.405 256.570 59.410 ;
        POLYGON 253.670 59.405 253.775 59.405 253.775 59.375 ;
        RECT 253.775 59.375 256.570 59.405 ;
        POLYGON 256.570 59.465 256.720 59.375 256.570 59.375 ;
        POLYGON 259.595 59.465 259.620 59.465 259.620 59.445 ;
        RECT 259.620 59.445 263.020 59.465 ;
        POLYGON 259.620 59.445 259.655 59.445 259.655 59.405 ;
        RECT 259.655 59.405 263.020 59.445 ;
        POLYGON 259.655 59.405 259.685 59.405 259.685 59.375 ;
        RECT 259.685 59.375 263.020 59.405 ;
        POLYGON 253.775 59.375 253.785 59.375 253.785 59.370 ;
        RECT 253.785 59.370 256.720 59.375 ;
        RECT 244.330 59.355 246.775 59.370 ;
        POLYGON 246.775 59.370 246.820 59.370 246.775 59.355 ;
        POLYGON 253.785 59.370 253.795 59.370 253.795 59.365 ;
        RECT 253.795 59.365 256.720 59.370 ;
        POLYGON 253.800 59.365 253.825 59.365 253.825 59.355 ;
        RECT 253.825 59.355 256.720 59.365 ;
        RECT 244.330 59.350 246.750 59.355 ;
        RECT 238.965 59.270 241.585 59.350 ;
        POLYGON 241.585 59.350 241.670 59.350 241.585 59.270 ;
        POLYGON 244.260 59.350 244.260 59.305 244.195 59.305 ;
        RECT 244.260 59.345 246.750 59.350 ;
        POLYGON 246.750 59.355 246.775 59.355 246.750 59.345 ;
        POLYGON 253.825 59.355 253.850 59.355 253.850 59.345 ;
        RECT 253.850 59.345 256.720 59.355 ;
        RECT 244.260 59.320 246.685 59.345 ;
        POLYGON 246.685 59.345 246.750 59.345 246.685 59.320 ;
        POLYGON 253.850 59.345 253.895 59.345 253.895 59.330 ;
        RECT 253.895 59.330 256.720 59.345 ;
        POLYGON 253.895 59.330 253.920 59.330 253.920 59.320 ;
        RECT 253.920 59.320 256.720 59.330 ;
        RECT 244.260 59.305 246.545 59.320 ;
        POLYGON 244.195 59.305 244.195 59.270 244.140 59.270 ;
        RECT 244.195 59.270 246.545 59.305 ;
        RECT 238.965 59.160 241.480 59.270 ;
        POLYGON 241.480 59.270 241.585 59.270 241.480 59.160 ;
        POLYGON 244.140 59.270 244.140 59.160 243.975 59.160 ;
        RECT 244.140 59.260 246.545 59.270 ;
        POLYGON 246.545 59.320 246.685 59.320 246.545 59.260 ;
        POLYGON 253.925 59.320 254.010 59.320 254.010 59.290 ;
        RECT 254.010 59.290 256.720 59.320 ;
        POLYGON 254.015 59.290 254.030 59.290 254.030 59.280 ;
        RECT 254.030 59.280 256.720 59.290 ;
        POLYGON 254.030 59.280 254.080 59.280 254.080 59.260 ;
        RECT 254.080 59.260 256.720 59.280 ;
        RECT 244.140 59.255 246.540 59.260 ;
        POLYGON 246.540 59.260 246.545 59.260 246.540 59.255 ;
        POLYGON 254.080 59.260 254.090 59.260 254.090 59.255 ;
        RECT 254.090 59.255 256.720 59.260 ;
        RECT 244.140 59.225 246.460 59.255 ;
        POLYGON 246.460 59.255 246.535 59.255 246.460 59.225 ;
        POLYGON 254.090 59.255 254.170 59.255 254.170 59.225 ;
        RECT 254.170 59.245 256.720 59.255 ;
        POLYGON 256.720 59.375 256.920 59.245 256.720 59.245 ;
        POLYGON 259.685 59.375 259.815 59.375 259.815 59.260 ;
        RECT 259.815 59.325 263.020 59.375 ;
        POLYGON 263.020 59.490 263.145 59.325 263.020 59.325 ;
        POLYGON 267.710 59.490 267.780 59.490 267.780 59.380 ;
        RECT 267.780 59.380 275.095 59.490 ;
        POLYGON 267.780 59.380 267.810 59.380 267.810 59.330 ;
        RECT 267.810 59.325 275.095 59.380 ;
        RECT 259.815 59.260 263.145 59.325 ;
        POLYGON 259.815 59.260 259.830 59.260 259.830 59.245 ;
        RECT 259.830 59.245 263.145 59.260 ;
        RECT 254.170 59.235 256.920 59.245 ;
        POLYGON 256.920 59.245 256.930 59.235 256.920 59.235 ;
        POLYGON 259.830 59.245 259.840 59.245 259.840 59.235 ;
        RECT 259.840 59.235 263.145 59.245 ;
        RECT 254.170 59.225 256.930 59.235 ;
        RECT 244.140 59.160 246.310 59.225 ;
        RECT 238.965 59.150 241.465 59.160 ;
        POLYGON 241.465 59.160 241.480 59.160 241.465 59.150 ;
        POLYGON 243.975 59.160 243.975 59.150 243.960 59.150 ;
        RECT 243.975 59.155 246.310 59.160 ;
        POLYGON 246.310 59.225 246.460 59.225 246.310 59.155 ;
        POLYGON 254.170 59.225 254.185 59.225 254.185 59.220 ;
        RECT 254.185 59.220 256.930 59.225 ;
        POLYGON 254.185 59.220 254.220 59.220 254.220 59.210 ;
        RECT 254.220 59.210 256.930 59.220 ;
        POLYGON 254.220 59.210 254.230 59.210 254.230 59.205 ;
        RECT 254.230 59.205 256.930 59.210 ;
        POLYGON 254.230 59.205 254.280 59.205 254.280 59.185 ;
        RECT 254.280 59.185 256.930 59.205 ;
        POLYGON 254.280 59.185 254.345 59.185 254.345 59.155 ;
        RECT 254.345 59.155 256.930 59.185 ;
        RECT 243.975 59.150 246.250 59.155 ;
        RECT 238.965 59.080 241.295 59.150 ;
        POLYGON 238.705 59.080 238.705 59.065 238.695 59.065 ;
        RECT 238.705 59.065 241.295 59.080 ;
        RECT 230.505 59.005 235.160 59.065 ;
        POLYGON 235.160 59.065 235.190 59.065 235.160 59.005 ;
        POLYGON 238.695 59.065 238.695 59.005 238.650 59.005 ;
        RECT 238.695 59.005 241.295 59.065 ;
        RECT 230.505 59.000 235.135 59.005 ;
        RECT 206.245 58.610 222.515 58.990 ;
        POLYGON 222.515 58.990 222.585 58.990 222.515 58.610 ;
        POLYGON 230.375 58.995 230.375 58.735 230.285 58.735 ;
        RECT 230.375 58.965 235.135 59.000 ;
        POLYGON 235.135 59.005 235.160 59.005 235.135 58.965 ;
        POLYGON 238.650 59.005 238.650 58.965 238.620 58.965 ;
        RECT 238.650 58.970 241.295 59.005 ;
        POLYGON 241.295 59.150 241.465 59.150 241.295 58.970 ;
        POLYGON 243.960 59.150 243.960 59.145 243.955 59.145 ;
        RECT 243.960 59.145 246.250 59.150 ;
        POLYGON 243.955 59.145 243.955 59.065 243.840 59.065 ;
        RECT 243.955 59.125 246.250 59.145 ;
        POLYGON 246.250 59.155 246.310 59.155 246.250 59.125 ;
        POLYGON 254.345 59.155 254.415 59.155 254.415 59.125 ;
        RECT 254.415 59.125 256.930 59.155 ;
        RECT 243.955 59.120 246.240 59.125 ;
        POLYGON 246.240 59.125 246.245 59.125 246.240 59.120 ;
        POLYGON 254.415 59.125 254.425 59.125 254.425 59.120 ;
        RECT 254.425 59.120 256.930 59.125 ;
        RECT 243.955 59.065 245.945 59.120 ;
        POLYGON 243.840 59.065 243.840 58.970 243.710 58.970 ;
        RECT 243.840 58.970 245.945 59.065 ;
        RECT 238.650 58.965 241.270 58.970 ;
        RECT 230.375 58.735 234.965 58.965 ;
        POLYGON 230.285 58.735 230.285 58.610 230.245 58.610 ;
        RECT 230.285 58.610 234.965 58.735 ;
        POLYGON 234.965 58.965 235.135 58.965 234.965 58.615 ;
        POLYGON 238.620 58.965 238.620 58.945 238.605 58.945 ;
        RECT 238.620 58.945 241.270 58.965 ;
        POLYGON 241.270 58.970 241.295 58.970 241.270 58.945 ;
        POLYGON 243.710 58.970 243.710 58.945 243.675 58.945 ;
        RECT 243.710 58.965 245.945 58.970 ;
        POLYGON 245.945 59.120 246.235 59.120 245.945 58.965 ;
        POLYGON 254.425 59.120 254.520 59.120 254.520 59.080 ;
        RECT 254.520 59.080 256.930 59.120 ;
        POLYGON 254.520 59.080 254.545 59.080 254.545 59.070 ;
        RECT 254.545 59.075 256.930 59.080 ;
        POLYGON 256.930 59.235 257.165 59.075 256.930 59.075 ;
        POLYGON 259.840 59.235 260.000 59.235 260.000 59.075 ;
        RECT 260.000 59.205 263.145 59.235 ;
        POLYGON 263.145 59.325 263.240 59.205 263.145 59.205 ;
        POLYGON 267.810 59.325 267.885 59.325 267.885 59.205 ;
        RECT 267.885 59.240 275.095 59.325 ;
        POLYGON 275.095 59.565 275.260 59.240 275.095 59.240 ;
        POLYGON 287.775 59.565 287.810 59.565 287.810 59.255 ;
        RECT 287.810 59.240 303.120 59.565 ;
        RECT 267.885 59.205 275.260 59.240 ;
        RECT 260.000 59.075 263.240 59.205 ;
        RECT 254.545 59.070 257.165 59.075 ;
        POLYGON 254.550 59.070 254.755 59.070 254.755 58.970 ;
        RECT 254.755 59.000 257.165 59.070 ;
        POLYGON 257.165 59.075 257.275 59.000 257.165 59.000 ;
        POLYGON 260.000 59.075 260.080 59.075 260.080 59.000 ;
        RECT 260.080 59.000 263.240 59.075 ;
        RECT 254.755 58.980 257.275 59.000 ;
        POLYGON 257.275 59.000 257.300 58.980 257.275 58.980 ;
        POLYGON 260.080 59.000 260.100 59.000 260.100 58.980 ;
        RECT 260.100 58.980 263.240 59.000 ;
        RECT 254.755 58.970 257.300 58.980 ;
        POLYGON 254.760 58.970 254.765 58.970 254.765 58.965 ;
        RECT 254.765 58.965 257.300 58.970 ;
        RECT 243.710 58.945 245.875 58.965 ;
        POLYGON 238.605 58.945 238.605 58.615 238.385 58.615 ;
        RECT 238.605 58.745 241.090 58.945 ;
        POLYGON 241.090 58.945 241.270 58.945 241.090 58.745 ;
        POLYGON 243.675 58.945 243.675 58.935 243.660 58.935 ;
        RECT 243.675 58.935 245.875 58.945 ;
        POLYGON 243.660 58.935 243.660 58.920 243.645 58.920 ;
        RECT 243.660 58.930 245.875 58.935 ;
        POLYGON 245.875 58.965 245.945 58.965 245.875 58.930 ;
        POLYGON 254.765 58.965 254.830 58.965 254.830 58.930 ;
        RECT 254.830 58.950 257.300 58.965 ;
        POLYGON 257.300 58.980 257.345 58.950 257.300 58.950 ;
        POLYGON 260.100 58.980 260.130 58.980 260.130 58.950 ;
        RECT 260.130 58.950 263.240 58.980 ;
        RECT 254.830 58.930 257.345 58.950 ;
        RECT 243.660 58.920 245.815 58.930 ;
        POLYGON 243.645 58.920 243.645 58.805 243.495 58.805 ;
        RECT 243.645 58.895 245.815 58.920 ;
        POLYGON 245.815 58.930 245.875 58.930 245.815 58.895 ;
        POLYGON 254.830 58.930 254.860 58.930 254.860 58.915 ;
        RECT 254.860 58.915 257.345 58.930 ;
        POLYGON 254.865 58.915 254.900 58.915 254.900 58.895 ;
        RECT 254.900 58.895 257.345 58.915 ;
        RECT 243.645 58.805 245.660 58.895 ;
        POLYGON 245.660 58.895 245.815 58.895 245.660 58.805 ;
        POLYGON 250.405 58.895 250.405 58.890 249.890 58.890 ;
        RECT 250.405 58.890 250.435 58.895 ;
        POLYGON 249.860 58.890 249.860 58.875 249.695 58.875 ;
        RECT 249.860 58.875 250.435 58.890 ;
        POLYGON 250.435 58.895 250.915 58.875 250.435 58.875 ;
        POLYGON 254.900 58.895 254.940 58.895 254.940 58.875 ;
        RECT 254.940 58.875 257.345 58.895 ;
        POLYGON 249.655 58.875 249.655 58.855 249.380 58.855 ;
        RECT 249.655 58.870 250.915 58.875 ;
        POLYGON 250.915 58.875 251.005 58.870 250.915 58.870 ;
        POLYGON 254.940 58.875 254.950 58.875 254.950 58.870 ;
        RECT 254.950 58.870 257.345 58.875 ;
        RECT 249.655 58.865 251.005 58.870 ;
        POLYGON 251.005 58.870 251.060 58.865 251.005 58.865 ;
        POLYGON 254.950 58.870 254.960 58.870 254.960 58.865 ;
        RECT 254.960 58.865 257.345 58.870 ;
        RECT 249.655 58.855 251.065 58.865 ;
        POLYGON 249.380 58.855 249.380 58.845 249.290 58.845 ;
        RECT 249.380 58.845 251.065 58.855 ;
        POLYGON 249.290 58.845 249.290 58.805 248.965 58.805 ;
        RECT 249.290 58.840 251.065 58.845 ;
        POLYGON 251.065 58.865 251.345 58.840 251.065 58.840 ;
        POLYGON 254.960 58.865 255.005 58.865 255.005 58.840 ;
        RECT 255.005 58.840 257.345 58.865 ;
        RECT 249.290 58.830 251.350 58.840 ;
        POLYGON 251.350 58.840 251.425 58.830 251.350 58.830 ;
        POLYGON 255.005 58.840 255.025 58.840 255.025 58.830 ;
        RECT 255.025 58.830 257.345 58.840 ;
        RECT 249.290 58.810 251.425 58.830 ;
        POLYGON 251.425 58.830 251.580 58.810 251.425 58.810 ;
        POLYGON 255.025 58.830 255.065 58.830 255.065 58.810 ;
        RECT 255.065 58.810 257.345 58.830 ;
        RECT 249.290 58.805 251.580 58.810 ;
        POLYGON 251.580 58.810 251.605 58.805 251.580 58.805 ;
        POLYGON 255.065 58.810 255.075 58.810 255.075 58.805 ;
        RECT 255.075 58.805 257.345 58.810 ;
        POLYGON 243.495 58.805 243.495 58.745 243.415 58.745 ;
        RECT 243.495 58.760 245.585 58.805 ;
        POLYGON 245.585 58.805 245.660 58.805 245.585 58.760 ;
        POLYGON 248.935 58.805 248.935 58.795 248.875 58.795 ;
        RECT 248.935 58.795 251.615 58.805 ;
        POLYGON 248.875 58.795 248.875 58.770 248.735 58.770 ;
        RECT 248.875 58.770 251.615 58.795 ;
        POLYGON 251.615 58.805 251.860 58.770 251.615 58.770 ;
        POLYGON 255.075 58.805 255.145 58.805 255.145 58.770 ;
        RECT 255.145 58.770 257.345 58.805 ;
        POLYGON 248.735 58.770 248.735 58.760 248.660 58.760 ;
        RECT 248.735 58.760 251.860 58.770 ;
        POLYGON 251.860 58.770 251.925 58.760 251.860 58.760 ;
        POLYGON 255.145 58.770 255.165 58.770 255.165 58.760 ;
        RECT 255.165 58.765 257.345 58.770 ;
        POLYGON 257.345 58.950 257.595 58.765 257.345 58.765 ;
        POLYGON 260.130 58.950 260.150 58.950 260.150 58.930 ;
        RECT 260.150 58.930 263.240 58.950 ;
        POLYGON 260.150 58.930 260.290 58.930 260.290 58.785 ;
        RECT 260.290 58.875 263.240 58.930 ;
        POLYGON 263.240 59.205 263.495 58.875 263.240 58.875 ;
        POLYGON 267.885 59.205 268.090 59.205 268.090 58.875 ;
        RECT 268.090 58.875 275.260 59.205 ;
        RECT 260.290 58.785 263.495 58.875 ;
        POLYGON 260.290 58.785 260.305 58.785 260.305 58.765 ;
        RECT 260.305 58.765 263.495 58.785 ;
        RECT 255.165 58.760 257.595 58.765 ;
        RECT 243.495 58.745 245.510 58.760 ;
        RECT 238.605 58.660 241.015 58.745 ;
        POLYGON 241.015 58.745 241.090 58.745 241.015 58.660 ;
        POLYGON 243.415 58.745 243.415 58.715 243.375 58.715 ;
        RECT 243.415 58.715 245.510 58.745 ;
        POLYGON 245.510 58.760 245.580 58.760 245.510 58.715 ;
        POLYGON 248.655 58.760 248.655 58.715 248.410 58.715 ;
        RECT 248.655 58.740 251.925 58.760 ;
        POLYGON 251.925 58.760 252.040 58.740 251.925 58.740 ;
        POLYGON 255.165 58.760 255.195 58.760 255.195 58.740 ;
        RECT 255.195 58.750 257.595 58.760 ;
        POLYGON 257.595 58.765 257.615 58.750 257.595 58.750 ;
        POLYGON 260.305 58.765 260.320 58.765 260.320 58.750 ;
        RECT 260.320 58.750 263.495 58.765 ;
        RECT 255.195 58.740 257.615 58.750 ;
        RECT 248.655 58.725 252.040 58.740 ;
        POLYGON 252.040 58.740 252.095 58.725 252.040 58.725 ;
        POLYGON 255.195 58.740 255.220 58.740 255.220 58.725 ;
        RECT 255.220 58.725 257.615 58.740 ;
        RECT 248.655 58.720 252.100 58.725 ;
        POLYGON 252.100 58.725 252.145 58.720 252.100 58.720 ;
        POLYGON 255.220 58.725 255.230 58.725 255.230 58.720 ;
        RECT 255.230 58.720 257.615 58.725 ;
        RECT 248.655 58.715 252.145 58.720 ;
        POLYGON 243.375 58.715 243.375 58.660 243.310 58.660 ;
        RECT 243.375 58.660 245.380 58.715 ;
        RECT 238.605 58.655 241.010 58.660 ;
        POLYGON 241.010 58.660 241.015 58.660 241.010 58.655 ;
        POLYGON 243.310 58.660 243.310 58.655 243.305 58.655 ;
        RECT 243.310 58.655 245.380 58.660 ;
        RECT 238.605 58.615 240.970 58.655 ;
        RECT 238.385 58.610 240.970 58.615 ;
        POLYGON 240.970 58.655 241.010 58.655 240.970 58.610 ;
        POLYGON 243.305 58.655 243.305 58.610 243.250 58.610 ;
        RECT 243.305 58.630 245.380 58.655 ;
        POLYGON 245.380 58.715 245.510 58.715 245.380 58.630 ;
        POLYGON 248.410 58.715 248.410 58.710 248.380 58.710 ;
        RECT 248.410 58.710 252.145 58.715 ;
        POLYGON 248.370 58.710 248.370 58.695 248.315 58.695 ;
        RECT 248.370 58.695 252.145 58.710 ;
        POLYGON 248.315 58.695 248.315 58.690 248.295 58.690 ;
        RECT 248.315 58.690 252.145 58.695 ;
        POLYGON 248.295 58.690 248.295 58.670 248.190 58.670 ;
        RECT 248.295 58.680 252.145 58.690 ;
        POLYGON 252.145 58.720 252.325 58.680 252.145 58.680 ;
        POLYGON 255.230 58.720 255.300 58.720 255.300 58.680 ;
        RECT 255.300 58.700 257.615 58.720 ;
        POLYGON 257.615 58.750 257.675 58.700 257.615 58.700 ;
        POLYGON 260.320 58.750 260.370 58.750 260.370 58.700 ;
        RECT 260.370 58.745 263.495 58.750 ;
        POLYGON 263.495 58.875 263.600 58.745 263.495 58.745 ;
        POLYGON 268.090 58.875 268.170 58.875 268.170 58.745 ;
        RECT 268.170 58.745 275.260 58.875 ;
        RECT 260.370 58.700 263.600 58.745 ;
        RECT 255.300 58.680 257.675 58.700 ;
        RECT 248.295 58.675 252.325 58.680 ;
        POLYGON 252.325 58.680 252.350 58.675 252.325 58.675 ;
        POLYGON 255.300 58.680 255.305 58.680 255.305 58.675 ;
        RECT 255.305 58.675 257.675 58.680 ;
        RECT 248.295 58.670 252.350 58.675 ;
        POLYGON 248.190 58.670 248.190 58.645 248.100 58.645 ;
        RECT 248.190 58.665 252.350 58.670 ;
        POLYGON 252.350 58.675 252.415 58.665 252.350 58.665 ;
        POLYGON 255.305 58.675 255.325 58.675 255.325 58.665 ;
        RECT 255.325 58.665 257.675 58.675 ;
        RECT 248.190 58.645 252.415 58.665 ;
        POLYGON 248.100 58.645 248.100 58.630 248.035 58.630 ;
        RECT 248.100 58.630 252.415 58.645 ;
        POLYGON 252.415 58.665 252.545 58.630 252.415 58.630 ;
        POLYGON 255.325 58.665 255.385 58.665 255.385 58.630 ;
        RECT 255.385 58.630 257.675 58.665 ;
        RECT 243.305 58.610 245.350 58.630 ;
        POLYGON 245.350 58.630 245.380 58.630 245.350 58.610 ;
        POLYGON 248.035 58.630 248.035 58.625 248.010 58.625 ;
        RECT 248.035 58.625 252.545 58.630 ;
        POLYGON 248.010 58.625 248.010 58.610 247.940 58.610 ;
        RECT 248.010 58.610 252.545 58.625 ;
        POLYGON 252.545 58.630 252.635 58.610 252.545 58.610 ;
        POLYGON 255.385 58.630 255.420 58.630 255.420 58.610 ;
        RECT 255.420 58.610 257.675 58.630 ;
        POLYGON 257.675 58.700 257.785 58.610 257.675 58.610 ;
        POLYGON 260.370 58.700 260.385 58.700 260.385 58.685 ;
        RECT 260.385 58.685 263.600 58.700 ;
        POLYGON 260.385 58.685 260.420 58.685 260.420 58.645 ;
        RECT 260.420 58.645 263.600 58.685 ;
        POLYGON 260.420 58.645 260.455 58.645 260.455 58.610 ;
        RECT 260.455 58.610 263.600 58.645 ;
        POLYGON 263.600 58.745 263.690 58.610 263.600 58.610 ;
        POLYGON 268.170 58.745 268.250 58.745 268.250 58.615 ;
        RECT 268.250 58.610 275.260 58.745 ;
        POLYGON 275.260 59.240 275.550 58.610 275.260 58.610 ;
        POLYGON 287.810 59.240 287.880 59.240 287.880 58.610 ;
        RECT 206.235 58.605 222.515 58.610 ;
        RECT 180.675 58.580 194.980 58.590 ;
        POLYGON 194.980 58.590 194.985 58.580 194.980 58.580 ;
        RECT 180.675 58.375 194.985 58.580 ;
        RECT 168.890 58.340 173.390 58.375 ;
        POLYGON 168.890 58.340 168.930 58.340 168.930 58.275 ;
        RECT 168.930 58.275 173.390 58.340 ;
        POLYGON 168.930 58.275 168.945 58.275 168.945 58.250 ;
        RECT 168.945 58.250 173.390 58.275 ;
        RECT 163.245 58.235 165.790 58.250 ;
        POLYGON 163.245 58.235 163.325 58.235 163.325 58.155 ;
        RECT 163.325 58.185 165.790 58.235 ;
        POLYGON 165.790 58.250 165.845 58.185 165.790 58.185 ;
        POLYGON 168.945 58.250 168.965 58.250 168.965 58.225 ;
        RECT 168.965 58.225 173.390 58.250 ;
        POLYGON 168.965 58.225 168.990 58.225 168.990 58.185 ;
        RECT 168.990 58.185 173.390 58.225 ;
        RECT 163.325 58.155 165.845 58.185 ;
        RECT 158.965 58.140 161.130 58.155 ;
        POLYGON 158.965 58.140 158.985 58.140 158.985 58.130 ;
        RECT 158.985 58.130 161.130 58.140 ;
        RECT 149.650 58.115 151.675 58.130 ;
        POLYGON 151.675 58.130 151.705 58.130 151.675 58.120 ;
        POLYGON 158.985 58.130 159.010 58.130 159.010 58.120 ;
        RECT 159.010 58.120 161.130 58.130 ;
        POLYGON 159.010 58.120 159.025 58.120 159.025 58.115 ;
        RECT 159.025 58.115 161.130 58.120 ;
        RECT 149.650 58.060 151.515 58.115 ;
        RECT 117.340 57.990 147.320 58.060 ;
        POLYGON 117.320 57.990 117.320 57.510 117.310 57.510 ;
        RECT 117.320 57.775 147.320 57.990 ;
        POLYGON 147.320 58.060 147.605 58.060 147.320 57.775 ;
        POLYGON 149.550 58.060 149.550 57.970 149.435 57.970 ;
        RECT 149.550 58.040 151.515 58.060 ;
        POLYGON 151.515 58.115 151.670 58.115 151.515 58.040 ;
        POLYGON 155.065 58.115 155.065 58.110 154.975 58.110 ;
        RECT 155.065 58.110 155.350 58.115 ;
        POLYGON 155.350 58.115 155.360 58.110 155.350 58.110 ;
        POLYGON 159.025 58.115 159.035 58.115 159.035 58.110 ;
        RECT 159.035 58.110 161.130 58.115 ;
        POLYGON 161.130 58.155 161.195 58.110 161.130 58.110 ;
        POLYGON 163.325 58.155 163.375 58.155 163.375 58.110 ;
        RECT 163.375 58.110 165.845 58.155 ;
        POLYGON 154.915 58.110 154.915 58.105 154.850 58.105 ;
        RECT 154.915 58.105 155.540 58.110 ;
        POLYGON 154.845 58.105 154.845 58.100 154.625 58.100 ;
        RECT 154.845 58.100 155.540 58.105 ;
        POLYGON 154.625 58.100 154.625 58.080 154.425 58.080 ;
        RECT 154.625 58.080 155.540 58.100 ;
        POLYGON 155.540 58.110 155.920 58.080 155.540 58.080 ;
        POLYGON 159.035 58.110 159.100 58.110 159.100 58.080 ;
        RECT 159.100 58.100 161.195 58.110 ;
        POLYGON 161.195 58.110 161.210 58.100 161.195 58.100 ;
        POLYGON 163.375 58.110 163.385 58.110 163.385 58.100 ;
        RECT 163.385 58.100 165.845 58.110 ;
        RECT 159.100 58.080 161.210 58.100 ;
        POLYGON 154.410 58.080 154.410 58.065 154.280 58.065 ;
        RECT 154.410 58.075 155.945 58.080 ;
        POLYGON 155.945 58.080 155.995 58.075 155.945 58.075 ;
        POLYGON 159.100 58.080 159.110 58.080 159.110 58.075 ;
        RECT 159.110 58.075 161.210 58.080 ;
        RECT 154.410 58.065 155.995 58.075 ;
        POLYGON 154.280 58.065 154.280 58.055 154.185 58.055 ;
        RECT 154.280 58.060 155.995 58.065 ;
        POLYGON 155.995 58.075 156.100 58.060 155.995 58.060 ;
        POLYGON 159.110 58.075 159.140 58.075 159.140 58.060 ;
        RECT 159.140 58.060 161.210 58.075 ;
        POLYGON 161.210 58.100 161.265 58.060 161.210 58.060 ;
        POLYGON 163.385 58.100 163.395 58.100 163.395 58.095 ;
        RECT 163.395 58.095 165.845 58.100 ;
        POLYGON 163.395 58.095 163.440 58.095 163.440 58.060 ;
        RECT 163.440 58.060 165.845 58.095 ;
        RECT 154.280 58.055 156.105 58.060 ;
        POLYGON 154.180 58.055 154.180 58.040 154.085 58.040 ;
        RECT 154.180 58.040 156.105 58.055 ;
        RECT 149.550 58.010 151.445 58.040 ;
        POLYGON 151.445 58.040 151.510 58.040 151.445 58.010 ;
        POLYGON 154.085 58.040 154.085 58.015 153.930 58.015 ;
        RECT 154.085 58.025 156.105 58.040 ;
        POLYGON 156.105 58.060 156.390 58.025 156.105 58.025 ;
        POLYGON 159.140 58.060 159.155 58.060 159.155 58.055 ;
        RECT 159.155 58.055 161.265 58.060 ;
        POLYGON 159.155 58.055 159.215 58.055 159.215 58.025 ;
        RECT 159.215 58.025 161.265 58.055 ;
        RECT 154.085 58.020 156.390 58.025 ;
        POLYGON 156.390 58.025 156.410 58.020 156.390 58.020 ;
        POLYGON 159.215 58.025 159.225 58.025 159.225 58.020 ;
        RECT 159.225 58.020 161.265 58.025 ;
        RECT 154.085 58.015 156.415 58.020 ;
        POLYGON 153.925 58.015 153.925 58.010 153.890 58.010 ;
        RECT 153.925 58.010 156.415 58.015 ;
        RECT 149.550 57.970 151.285 58.010 ;
        POLYGON 149.430 57.970 149.430 57.965 149.425 57.965 ;
        RECT 149.430 57.965 151.285 57.970 ;
        POLYGON 149.425 57.965 149.425 57.815 149.245 57.815 ;
        RECT 149.425 57.935 151.285 57.965 ;
        POLYGON 151.285 58.010 151.445 58.010 151.285 57.935 ;
        POLYGON 153.890 58.010 153.890 58.005 153.850 58.005 ;
        RECT 153.890 58.005 156.415 58.010 ;
        POLYGON 153.850 58.005 153.850 57.990 153.750 57.990 ;
        RECT 153.850 57.990 156.415 58.005 ;
        POLYGON 156.415 58.020 156.570 57.990 156.415 57.990 ;
        POLYGON 159.225 58.020 159.270 58.020 159.270 58.000 ;
        RECT 159.270 58.000 161.265 58.020 ;
        POLYGON 159.275 58.000 159.290 58.000 159.290 57.990 ;
        RECT 159.290 57.990 161.265 58.000 ;
        POLYGON 153.750 57.990 153.750 57.985 153.725 57.985 ;
        RECT 153.750 57.985 156.570 57.990 ;
        POLYGON 153.720 57.985 153.720 57.935 153.485 57.935 ;
        RECT 153.720 57.970 156.570 57.985 ;
        POLYGON 156.570 57.990 156.670 57.970 156.570 57.970 ;
        POLYGON 159.290 57.990 159.330 57.990 159.330 57.970 ;
        RECT 159.330 57.970 161.265 57.990 ;
        RECT 153.720 57.940 156.670 57.970 ;
        POLYGON 156.670 57.970 156.830 57.940 156.670 57.940 ;
        POLYGON 159.330 57.970 159.375 57.970 159.375 57.950 ;
        RECT 159.375 57.950 161.265 57.970 ;
        POLYGON 159.375 57.950 159.395 57.950 159.395 57.940 ;
        RECT 159.395 57.940 161.265 57.950 ;
        RECT 153.720 57.935 156.830 57.940 ;
        RECT 149.425 57.890 151.195 57.935 ;
        POLYGON 151.195 57.935 151.285 57.935 151.195 57.890 ;
        POLYGON 153.485 57.935 153.485 57.925 153.435 57.925 ;
        RECT 153.485 57.925 156.830 57.935 ;
        POLYGON 156.830 57.940 156.905 57.925 156.830 57.925 ;
        POLYGON 159.395 57.940 159.420 57.940 159.420 57.930 ;
        RECT 159.420 57.930 161.265 57.940 ;
        POLYGON 159.420 57.930 159.425 57.930 159.425 57.925 ;
        RECT 159.425 57.925 161.265 57.930 ;
        POLYGON 153.435 57.925 153.435 57.900 153.325 57.900 ;
        RECT 153.435 57.915 156.905 57.925 ;
        POLYGON 156.905 57.925 156.950 57.915 156.905 57.915 ;
        POLYGON 159.425 57.925 159.445 57.925 159.445 57.915 ;
        RECT 159.445 57.915 161.265 57.925 ;
        RECT 153.435 57.900 156.950 57.915 ;
        POLYGON 153.320 57.900 153.320 57.895 153.300 57.895 ;
        RECT 153.320 57.895 156.950 57.900 ;
        POLYGON 153.300 57.895 153.300 57.890 153.285 57.890 ;
        RECT 153.300 57.890 156.950 57.895 ;
        RECT 149.425 57.815 151.050 57.890 ;
        POLYGON 149.245 57.815 149.245 57.775 149.195 57.775 ;
        RECT 149.245 57.810 151.050 57.815 ;
        POLYGON 151.050 57.890 151.195 57.890 151.050 57.810 ;
        POLYGON 153.285 57.890 153.285 57.860 153.180 57.860 ;
        RECT 153.285 57.865 156.950 57.890 ;
        POLYGON 156.950 57.915 157.140 57.865 156.950 57.865 ;
        POLYGON 159.445 57.915 159.515 57.915 159.515 57.875 ;
        RECT 159.515 57.875 161.265 57.915 ;
        POLYGON 159.515 57.875 159.530 57.875 159.530 57.865 ;
        RECT 159.530 57.865 161.265 57.875 ;
        RECT 153.285 57.860 157.140 57.865 ;
        POLYGON 153.180 57.860 153.180 57.810 152.990 57.810 ;
        RECT 153.180 57.845 157.140 57.860 ;
        POLYGON 157.140 57.865 157.235 57.845 157.140 57.845 ;
        POLYGON 159.530 57.865 159.570 57.865 159.570 57.845 ;
        RECT 159.570 57.845 161.265 57.865 ;
        RECT 153.180 57.835 157.235 57.845 ;
        POLYGON 157.235 57.845 157.265 57.835 157.235 57.835 ;
        POLYGON 159.570 57.845 159.590 57.845 159.590 57.835 ;
        RECT 159.590 57.840 161.265 57.845 ;
        POLYGON 161.265 58.060 161.555 57.840 161.265 57.840 ;
        POLYGON 163.440 58.060 163.545 58.060 163.545 57.960 ;
        RECT 163.545 57.960 165.845 58.060 ;
        POLYGON 163.545 57.960 163.665 57.960 163.665 57.845 ;
        RECT 163.665 57.935 165.845 57.960 ;
        POLYGON 165.845 58.185 166.050 57.935 165.845 57.935 ;
        POLYGON 168.990 58.185 168.995 58.185 168.995 58.180 ;
        RECT 168.995 58.180 173.390 58.185 ;
        POLYGON 168.995 58.180 169.020 58.180 169.020 58.140 ;
        RECT 169.020 58.160 173.390 58.180 ;
        POLYGON 173.390 58.375 173.505 58.160 173.390 58.160 ;
        POLYGON 180.675 58.375 180.685 58.375 180.685 58.355 ;
        RECT 180.685 58.355 194.985 58.375 ;
        POLYGON 180.685 58.355 180.765 58.355 180.765 58.160 ;
        RECT 180.765 58.190 194.985 58.355 ;
        POLYGON 194.985 58.580 195.130 58.190 194.985 58.190 ;
        RECT 206.235 58.270 222.455 58.605 ;
        POLYGON 222.455 58.605 222.515 58.605 222.455 58.275 ;
        POLYGON 230.245 58.605 230.245 58.275 230.140 58.275 ;
        RECT 230.245 58.315 234.820 58.610 ;
        POLYGON 234.820 58.610 234.965 58.610 234.820 58.315 ;
        POLYGON 238.385 58.610 238.385 58.590 238.370 58.590 ;
        RECT 238.385 58.590 240.915 58.610 ;
        POLYGON 238.370 58.590 238.370 58.515 238.320 58.515 ;
        RECT 238.370 58.545 240.915 58.590 ;
        POLYGON 240.915 58.610 240.970 58.610 240.915 58.545 ;
        POLYGON 243.250 58.610 243.250 58.560 243.190 58.560 ;
        RECT 243.250 58.560 245.265 58.610 ;
        POLYGON 243.190 58.560 243.190 58.545 243.170 58.545 ;
        RECT 243.190 58.555 245.265 58.560 ;
        POLYGON 245.265 58.610 245.350 58.610 245.265 58.555 ;
        POLYGON 247.940 58.610 247.940 58.600 247.895 58.600 ;
        RECT 247.940 58.600 252.635 58.610 ;
        POLYGON 247.895 58.600 247.895 58.585 247.840 58.585 ;
        RECT 247.895 58.590 252.635 58.600 ;
        POLYGON 252.635 58.610 252.700 58.590 252.635 58.590 ;
        POLYGON 255.420 58.610 255.455 58.610 255.455 58.590 ;
        RECT 255.455 58.590 257.785 58.610 ;
        RECT 247.895 58.585 252.705 58.590 ;
        POLYGON 247.840 58.585 247.840 58.555 247.740 58.555 ;
        RECT 247.840 58.575 252.705 58.585 ;
        POLYGON 252.705 58.590 252.760 58.575 252.705 58.575 ;
        POLYGON 255.460 58.590 255.485 58.590 255.485 58.575 ;
        RECT 255.485 58.575 257.785 58.590 ;
        RECT 247.840 58.555 252.760 58.575 ;
        RECT 243.190 58.545 245.150 58.555 ;
        RECT 238.370 58.515 240.830 58.545 ;
        POLYGON 238.320 58.515 238.320 58.315 238.185 58.315 ;
        RECT 238.320 58.445 240.830 58.515 ;
        POLYGON 240.830 58.545 240.915 58.545 240.830 58.445 ;
        POLYGON 243.170 58.545 243.170 58.535 243.160 58.535 ;
        RECT 243.170 58.535 245.150 58.545 ;
        POLYGON 243.160 58.535 243.160 58.490 243.100 58.490 ;
        RECT 243.160 58.490 245.150 58.535 ;
        POLYGON 243.100 58.490 243.100 58.445 243.050 58.445 ;
        RECT 243.100 58.485 245.150 58.490 ;
        POLYGON 245.150 58.555 245.260 58.555 245.150 58.485 ;
        POLYGON 247.740 58.555 247.740 58.535 247.665 58.535 ;
        RECT 247.740 58.540 252.760 58.555 ;
        POLYGON 252.760 58.575 252.895 58.540 252.760 58.540 ;
        POLYGON 255.485 58.575 255.505 58.575 255.505 58.565 ;
        RECT 255.505 58.565 257.785 58.575 ;
        POLYGON 255.505 58.565 255.540 58.565 255.540 58.540 ;
        RECT 255.540 58.540 257.785 58.565 ;
        RECT 247.740 58.535 252.895 58.540 ;
        POLYGON 252.895 58.540 252.905 58.535 252.895 58.535 ;
        POLYGON 255.540 58.540 255.550 58.540 255.550 58.535 ;
        RECT 255.550 58.535 257.785 58.540 ;
        POLYGON 247.665 58.535 247.665 58.510 247.590 58.510 ;
        RECT 247.665 58.515 252.905 58.535 ;
        POLYGON 252.905 58.535 252.980 58.515 252.905 58.515 ;
        POLYGON 255.550 58.535 255.580 58.535 255.580 58.515 ;
        RECT 255.580 58.515 257.785 58.535 ;
        RECT 247.665 58.510 252.980 58.515 ;
        POLYGON 247.590 58.510 247.590 58.485 247.505 58.485 ;
        RECT 247.590 58.485 252.980 58.510 ;
        RECT 243.100 58.455 245.110 58.485 ;
        POLYGON 245.110 58.485 245.150 58.485 245.110 58.455 ;
        POLYGON 247.505 58.485 247.505 58.465 247.425 58.465 ;
        RECT 247.505 58.465 252.980 58.485 ;
        POLYGON 247.425 58.465 247.425 58.455 247.395 58.455 ;
        RECT 247.425 58.455 252.980 58.465 ;
        POLYGON 252.980 58.515 253.165 58.455 252.980 58.455 ;
        POLYGON 255.580 58.515 255.670 58.515 255.670 58.455 ;
        RECT 255.670 58.495 257.785 58.515 ;
        POLYGON 257.785 58.610 257.935 58.495 257.785 58.495 ;
        POLYGON 260.455 58.610 260.490 58.610 260.490 58.575 ;
        RECT 260.490 58.575 263.690 58.610 ;
        POLYGON 260.490 58.575 260.560 58.575 260.560 58.495 ;
        RECT 260.560 58.495 263.690 58.575 ;
        RECT 255.670 58.455 257.935 58.495 ;
        RECT 243.100 58.445 244.900 58.455 ;
        RECT 238.320 58.350 240.755 58.445 ;
        POLYGON 240.755 58.445 240.830 58.445 240.755 58.350 ;
        POLYGON 243.050 58.445 243.050 58.350 242.945 58.350 ;
        RECT 243.050 58.350 244.900 58.445 ;
        RECT 238.320 58.335 240.745 58.350 ;
        POLYGON 240.745 58.350 240.755 58.350 240.745 58.335 ;
        POLYGON 242.945 58.350 242.945 58.335 242.930 58.335 ;
        RECT 242.945 58.335 244.900 58.350 ;
        RECT 238.320 58.315 240.630 58.335 ;
        RECT 230.245 58.275 234.760 58.315 ;
        RECT 180.765 58.160 195.130 58.190 ;
        RECT 169.020 58.140 173.505 58.160 ;
        POLYGON 169.020 58.140 169.080 58.140 169.080 58.050 ;
        RECT 169.080 58.050 173.505 58.140 ;
        POLYGON 169.080 58.050 169.085 58.050 169.085 58.045 ;
        RECT 169.085 58.045 173.505 58.050 ;
        POLYGON 169.085 58.045 169.150 58.045 169.150 57.940 ;
        RECT 169.150 57.935 173.505 58.045 ;
        RECT 163.665 57.875 166.050 57.935 ;
        POLYGON 166.050 57.935 166.095 57.875 166.050 57.875 ;
        POLYGON 169.150 57.935 169.160 57.935 169.160 57.925 ;
        RECT 169.160 57.925 173.505 57.935 ;
        POLYGON 169.160 57.925 169.190 57.925 169.190 57.875 ;
        RECT 169.190 57.875 173.505 57.925 ;
        RECT 163.665 57.845 166.095 57.875 ;
        POLYGON 163.665 57.845 163.670 57.845 163.670 57.840 ;
        RECT 163.670 57.840 166.095 57.845 ;
        RECT 159.590 57.835 161.555 57.840 ;
        POLYGON 161.555 57.840 161.565 57.835 161.555 57.835 ;
        POLYGON 163.670 57.840 163.675 57.840 163.675 57.835 ;
        RECT 163.675 57.835 166.095 57.840 ;
        RECT 153.180 57.810 157.265 57.835 ;
        RECT 149.245 57.775 150.950 57.810 ;
        RECT 117.320 57.730 147.285 57.775 ;
        POLYGON 147.285 57.775 147.320 57.775 147.285 57.730 ;
        POLYGON 149.195 57.775 149.195 57.730 149.145 57.730 ;
        RECT 149.195 57.760 150.950 57.775 ;
        POLYGON 150.950 57.810 151.050 57.810 150.950 57.760 ;
        POLYGON 152.990 57.810 152.990 57.800 152.950 57.800 ;
        RECT 152.990 57.800 157.265 57.810 ;
        POLYGON 152.945 57.800 152.945 57.785 152.900 57.785 ;
        RECT 152.945 57.795 157.265 57.800 ;
        POLYGON 157.265 57.835 157.395 57.795 157.265 57.795 ;
        POLYGON 159.590 57.835 159.670 57.835 159.670 57.795 ;
        RECT 159.670 57.820 161.565 57.835 ;
        POLYGON 161.565 57.835 161.585 57.820 161.565 57.820 ;
        POLYGON 163.675 57.835 163.690 57.835 163.690 57.820 ;
        RECT 163.690 57.820 166.095 57.835 ;
        RECT 159.670 57.795 161.585 57.820 ;
        RECT 152.945 57.785 157.395 57.795 ;
        POLYGON 152.895 57.785 152.895 57.760 152.820 57.760 ;
        RECT 152.895 57.760 157.395 57.785 ;
        POLYGON 157.395 57.795 157.510 57.760 157.395 57.760 ;
        POLYGON 159.670 57.795 159.680 57.795 159.680 57.790 ;
        RECT 159.680 57.790 161.585 57.795 ;
        POLYGON 159.680 57.790 159.730 57.790 159.730 57.760 ;
        RECT 159.730 57.760 161.585 57.790 ;
        RECT 149.195 57.735 150.910 57.760 ;
        POLYGON 150.910 57.760 150.950 57.760 150.910 57.735 ;
        POLYGON 152.820 57.760 152.820 57.735 152.745 57.735 ;
        RECT 152.820 57.735 157.515 57.760 ;
        RECT 149.195 57.730 150.860 57.735 ;
        RECT 117.320 57.675 147.230 57.730 ;
        POLYGON 147.230 57.730 147.285 57.730 147.230 57.675 ;
        POLYGON 149.145 57.730 149.145 57.685 149.090 57.685 ;
        RECT 149.145 57.710 150.860 57.730 ;
        POLYGON 150.860 57.735 150.910 57.735 150.860 57.710 ;
        POLYGON 152.745 57.735 152.745 57.710 152.670 57.710 ;
        RECT 152.745 57.710 157.515 57.735 ;
        RECT 149.145 57.685 150.705 57.710 ;
        POLYGON 149.090 57.685 149.090 57.675 149.080 57.675 ;
        RECT 149.090 57.675 150.705 57.685 ;
        RECT 117.320 57.565 147.130 57.675 ;
        POLYGON 147.130 57.675 147.230 57.675 147.130 57.565 ;
        POLYGON 149.080 57.675 149.080 57.565 148.955 57.565 ;
        RECT 149.080 57.620 150.705 57.675 ;
        POLYGON 150.705 57.710 150.860 57.710 150.705 57.620 ;
        POLYGON 152.670 57.710 152.670 57.705 152.655 57.705 ;
        RECT 152.670 57.705 157.515 57.710 ;
        POLYGON 157.515 57.760 157.695 57.705 157.515 57.705 ;
        POLYGON 159.730 57.760 159.750 57.760 159.750 57.750 ;
        RECT 159.750 57.750 161.585 57.760 ;
        POLYGON 159.750 57.750 159.825 57.750 159.825 57.705 ;
        RECT 159.825 57.745 161.585 57.750 ;
        POLYGON 161.585 57.820 161.675 57.745 161.585 57.745 ;
        POLYGON 163.690 57.820 163.765 57.820 163.765 57.745 ;
        RECT 163.765 57.755 166.095 57.820 ;
        POLYGON 166.095 57.875 166.190 57.755 166.095 57.755 ;
        POLYGON 169.190 57.875 169.260 57.875 169.260 57.755 ;
        RECT 169.260 57.755 173.505 57.875 ;
        RECT 163.765 57.745 166.190 57.755 ;
        RECT 159.825 57.705 161.675 57.745 ;
        POLYGON 152.655 57.705 152.655 57.645 152.485 57.645 ;
        RECT 152.655 57.670 157.700 57.705 ;
        POLYGON 157.700 57.705 157.790 57.670 157.700 57.670 ;
        POLYGON 159.825 57.705 159.885 57.705 159.885 57.670 ;
        RECT 159.885 57.670 161.675 57.705 ;
        RECT 152.655 57.645 157.790 57.670 ;
        POLYGON 152.485 57.645 152.485 57.640 152.460 57.640 ;
        RECT 152.485 57.640 157.790 57.645 ;
        POLYGON 157.790 57.670 157.875 57.640 157.790 57.640 ;
        POLYGON 159.885 57.670 159.940 57.670 159.940 57.640 ;
        RECT 159.940 57.640 161.675 57.670 ;
        POLYGON 152.460 57.640 152.460 57.620 152.410 57.620 ;
        RECT 152.460 57.620 157.880 57.640 ;
        RECT 149.080 57.565 150.595 57.620 ;
        RECT 117.320 57.520 147.090 57.565 ;
        POLYGON 147.090 57.565 147.130 57.565 147.090 57.520 ;
        POLYGON 148.955 57.565 148.955 57.550 148.940 57.550 ;
        RECT 148.955 57.550 150.595 57.565 ;
        POLYGON 150.595 57.620 150.705 57.620 150.595 57.550 ;
        POLYGON 152.410 57.620 152.410 57.550 152.235 57.550 ;
        RECT 152.410 57.570 157.880 57.620 ;
        POLYGON 157.880 57.640 158.065 57.570 157.880 57.570 ;
        POLYGON 159.940 57.640 160.055 57.640 160.055 57.570 ;
        RECT 160.055 57.570 161.675 57.640 ;
        POLYGON 161.675 57.745 161.890 57.570 161.675 57.570 ;
        POLYGON 163.765 57.745 163.830 57.745 163.830 57.680 ;
        RECT 163.830 57.680 166.190 57.745 ;
        POLYGON 163.830 57.680 163.915 57.680 163.915 57.585 ;
        RECT 163.915 57.595 166.190 57.680 ;
        POLYGON 166.190 57.755 166.310 57.595 166.190 57.595 ;
        POLYGON 169.260 57.755 169.355 57.755 169.355 57.600 ;
        RECT 169.355 57.595 173.505 57.755 ;
        RECT 163.915 57.585 166.310 57.595 ;
        POLYGON 163.915 57.585 163.930 57.585 163.930 57.570 ;
        RECT 163.930 57.570 166.310 57.585 ;
        RECT 152.410 57.550 158.070 57.570 ;
        POLYGON 158.070 57.570 158.130 57.550 158.070 57.550 ;
        POLYGON 160.055 57.570 160.085 57.570 160.085 57.550 ;
        RECT 160.085 57.550 161.890 57.570 ;
        POLYGON 148.940 57.550 148.940 57.545 148.930 57.545 ;
        RECT 148.940 57.545 150.545 57.550 ;
        POLYGON 148.930 57.545 148.930 57.520 148.905 57.520 ;
        RECT 148.930 57.520 150.545 57.545 ;
        POLYGON 150.545 57.550 150.595 57.550 150.545 57.520 ;
        POLYGON 152.235 57.550 152.235 57.545 152.225 57.545 ;
        RECT 152.235 57.545 158.130 57.550 ;
        POLYGON 152.225 57.545 152.225 57.520 152.165 57.520 ;
        RECT 152.225 57.520 158.130 57.545 ;
        RECT 117.320 57.510 147.035 57.520 ;
        RECT 117.310 57.460 147.035 57.510 ;
        POLYGON 147.035 57.520 147.090 57.520 147.035 57.460 ;
        POLYGON 148.905 57.520 148.905 57.460 148.840 57.460 ;
        RECT 148.905 57.490 150.500 57.520 ;
        POLYGON 150.500 57.520 150.545 57.520 150.500 57.490 ;
        POLYGON 152.165 57.520 152.165 57.515 152.150 57.515 ;
        RECT 152.165 57.515 158.130 57.520 ;
        POLYGON 152.150 57.515 152.150 57.490 152.090 57.490 ;
        RECT 152.150 57.500 158.130 57.515 ;
        POLYGON 158.130 57.550 158.240 57.500 158.130 57.500 ;
        POLYGON 160.085 57.550 160.130 57.550 160.130 57.525 ;
        RECT 160.130 57.535 161.890 57.550 ;
        POLYGON 161.890 57.570 161.925 57.535 161.890 57.535 ;
        POLYGON 163.930 57.570 163.965 57.570 163.965 57.535 ;
        RECT 163.965 57.535 166.310 57.570 ;
        RECT 160.130 57.525 161.925 57.535 ;
        POLYGON 160.130 57.525 160.160 57.525 160.160 57.505 ;
        RECT 160.160 57.505 161.925 57.525 ;
        POLYGON 160.165 57.505 160.170 57.505 160.170 57.500 ;
        RECT 160.170 57.500 161.925 57.505 ;
        RECT 152.150 57.490 158.240 57.500 ;
        RECT 148.905 57.470 150.465 57.490 ;
        POLYGON 150.465 57.490 150.495 57.490 150.465 57.470 ;
        POLYGON 152.090 57.490 152.090 57.485 152.075 57.485 ;
        RECT 152.090 57.485 158.240 57.490 ;
        POLYGON 152.075 57.485 152.075 57.470 152.040 57.470 ;
        RECT 152.075 57.470 158.240 57.485 ;
        RECT 148.905 57.460 150.230 57.470 ;
        POLYGON 111.175 57.055 111.200 56.390 111.175 56.390 ;
        POLYGON 117.310 57.455 117.310 56.390 117.290 56.390 ;
        RECT 117.310 57.260 146.865 57.460 ;
        POLYGON 146.865 57.460 147.035 57.460 146.865 57.260 ;
        POLYGON 148.840 57.460 148.840 57.390 148.760 57.390 ;
        RECT 148.840 57.390 150.230 57.460 ;
        POLYGON 148.760 57.390 148.760 57.280 148.645 57.280 ;
        RECT 148.760 57.315 150.230 57.390 ;
        POLYGON 150.230 57.470 150.465 57.470 150.230 57.315 ;
        POLYGON 152.040 57.470 152.040 57.445 151.985 57.445 ;
        RECT 152.040 57.455 158.240 57.470 ;
        POLYGON 158.240 57.500 158.340 57.455 158.240 57.455 ;
        POLYGON 160.170 57.500 160.185 57.500 160.185 57.490 ;
        RECT 160.185 57.490 161.925 57.500 ;
        POLYGON 160.185 57.490 160.195 57.490 160.195 57.485 ;
        RECT 160.195 57.485 161.925 57.490 ;
        POLYGON 160.195 57.485 160.235 57.485 160.235 57.455 ;
        RECT 160.235 57.455 161.925 57.485 ;
        RECT 152.040 57.450 158.345 57.455 ;
        POLYGON 158.345 57.455 158.355 57.450 158.345 57.450 ;
        POLYGON 160.235 57.455 160.245 57.455 160.245 57.450 ;
        RECT 160.245 57.450 161.925 57.455 ;
        RECT 152.040 57.445 158.355 57.450 ;
        POLYGON 151.985 57.445 151.985 57.410 151.910 57.410 ;
        RECT 151.985 57.430 158.355 57.445 ;
        RECT 151.985 57.425 155.075 57.430 ;
        POLYGON 155.075 57.430 155.170 57.430 155.075 57.425 ;
        POLYGON 155.505 57.430 155.540 57.430 155.540 57.425 ;
        RECT 155.540 57.425 158.355 57.430 ;
        RECT 151.985 57.420 155.010 57.425 ;
        POLYGON 155.010 57.425 155.065 57.425 155.010 57.420 ;
        POLYGON 155.565 57.425 155.695 57.425 155.695 57.420 ;
        RECT 155.695 57.420 158.355 57.425 ;
        RECT 151.985 57.410 154.785 57.420 ;
        POLYGON 154.785 57.420 154.905 57.420 154.785 57.410 ;
        POLYGON 155.695 57.420 155.810 57.420 155.810 57.410 ;
        RECT 155.810 57.410 158.355 57.420 ;
        POLYGON 151.910 57.410 151.910 57.315 151.705 57.315 ;
        RECT 151.910 57.405 154.775 57.410 ;
        POLYGON 154.775 57.410 154.785 57.410 154.775 57.405 ;
        POLYGON 155.850 57.410 155.890 57.410 155.890 57.405 ;
        RECT 155.890 57.405 158.355 57.410 ;
        RECT 151.910 57.395 154.640 57.405 ;
        POLYGON 154.640 57.405 154.770 57.405 154.640 57.395 ;
        POLYGON 155.890 57.405 155.935 57.405 155.935 57.400 ;
        RECT 155.935 57.400 158.355 57.405 ;
        POLYGON 155.955 57.400 155.995 57.400 155.995 57.395 ;
        RECT 155.995 57.395 158.355 57.400 ;
        RECT 151.910 57.385 154.565 57.395 ;
        POLYGON 154.565 57.395 154.625 57.395 154.565 57.385 ;
        POLYGON 155.995 57.395 156.085 57.395 156.085 57.385 ;
        RECT 156.085 57.385 158.355 57.395 ;
        RECT 151.910 57.380 154.515 57.385 ;
        POLYGON 154.515 57.385 154.565 57.385 154.515 57.380 ;
        POLYGON 156.085 57.385 156.115 57.385 156.115 57.380 ;
        RECT 156.115 57.380 158.355 57.385 ;
        RECT 151.910 57.365 154.375 57.380 ;
        POLYGON 154.375 57.380 154.515 57.380 154.375 57.365 ;
        POLYGON 156.115 57.380 156.150 57.380 156.150 57.375 ;
        RECT 156.150 57.375 158.355 57.380 ;
        POLYGON 156.155 57.375 156.220 57.375 156.220 57.370 ;
        RECT 156.220 57.370 158.355 57.375 ;
        POLYGON 156.220 57.370 156.245 57.370 156.245 57.365 ;
        RECT 156.245 57.365 158.355 57.370 ;
        POLYGON 158.355 57.450 158.550 57.365 158.355 57.365 ;
        POLYGON 160.245 57.450 160.370 57.450 160.370 57.365 ;
        RECT 160.370 57.445 161.925 57.450 ;
        POLYGON 161.925 57.535 162.025 57.445 161.925 57.445 ;
        POLYGON 163.965 57.535 164.010 57.535 164.010 57.490 ;
        RECT 164.010 57.490 166.310 57.535 ;
        POLYGON 166.310 57.595 166.390 57.490 166.310 57.490 ;
        POLYGON 169.355 57.595 169.375 57.595 169.375 57.570 ;
        RECT 169.375 57.570 173.505 57.595 ;
        POLYGON 169.375 57.570 169.420 57.570 169.420 57.495 ;
        RECT 169.420 57.525 173.505 57.570 ;
        POLYGON 173.505 58.160 173.850 57.525 173.505 57.525 ;
        POLYGON 180.765 58.160 180.925 58.160 180.925 57.780 ;
        RECT 180.925 57.935 195.130 58.160 ;
        POLYGON 195.130 58.190 195.225 57.935 195.130 57.935 ;
        RECT 180.925 57.780 195.225 57.935 ;
        POLYGON 206.235 58.190 206.235 58.100 206.230 58.100 ;
        RECT 206.235 58.100 222.435 58.270 ;
        POLYGON 222.435 58.270 222.455 58.270 222.435 58.110 ;
        POLYGON 230.140 58.265 230.140 58.190 230.115 58.190 ;
        RECT 230.140 58.190 234.760 58.275 ;
        POLYGON 234.760 58.315 234.820 58.315 234.760 58.195 ;
        POLYGON 238.185 58.315 238.185 58.240 238.135 58.240 ;
        RECT 238.185 58.240 240.630 58.315 ;
        POLYGON 238.135 58.240 238.135 58.195 238.110 58.195 ;
        RECT 238.135 58.195 240.630 58.240 ;
        POLYGON 238.110 58.195 238.110 58.190 238.105 58.190 ;
        RECT 238.110 58.190 240.630 58.195 ;
        POLYGON 240.630 58.335 240.745 58.335 240.630 58.190 ;
        POLYGON 242.930 58.335 242.930 58.255 242.840 58.255 ;
        RECT 242.930 58.305 244.900 58.335 ;
        POLYGON 244.900 58.455 245.110 58.455 244.900 58.310 ;
        POLYGON 247.395 58.455 247.395 58.435 247.340 58.435 ;
        RECT 247.395 58.435 253.165 58.455 ;
        POLYGON 247.340 58.435 247.340 58.430 247.335 58.430 ;
        RECT 247.340 58.430 253.165 58.435 ;
        POLYGON 253.165 58.455 253.245 58.430 253.165 58.430 ;
        POLYGON 255.670 58.455 255.710 58.455 255.710 58.430 ;
        RECT 255.710 58.430 257.935 58.455 ;
        POLYGON 257.935 58.495 258.010 58.430 257.935 58.430 ;
        POLYGON 260.560 58.495 260.615 58.495 260.615 58.430 ;
        RECT 260.615 58.430 263.690 58.495 ;
        POLYGON 247.335 58.430 247.335 58.400 247.245 58.400 ;
        RECT 247.335 58.400 253.250 58.430 ;
        POLYGON 247.245 58.400 247.245 58.385 247.195 58.385 ;
        RECT 247.245 58.395 253.250 58.400 ;
        POLYGON 253.250 58.430 253.355 58.395 253.250 58.395 ;
        POLYGON 255.710 58.430 255.735 58.430 255.735 58.415 ;
        RECT 255.735 58.415 258.010 58.430 ;
        POLYGON 255.740 58.415 255.770 58.415 255.770 58.395 ;
        RECT 255.770 58.400 258.010 58.415 ;
        POLYGON 258.010 58.430 258.050 58.400 258.010 58.400 ;
        POLYGON 260.615 58.430 260.640 58.430 260.640 58.405 ;
        RECT 260.640 58.425 263.690 58.430 ;
        POLYGON 263.690 58.610 263.820 58.425 263.690 58.425 ;
        POLYGON 268.250 58.610 268.270 58.610 268.270 58.585 ;
        RECT 268.270 58.585 275.550 58.610 ;
        POLYGON 268.270 58.585 268.355 58.585 268.355 58.425 ;
        RECT 268.355 58.430 275.550 58.585 ;
        POLYGON 275.550 58.610 275.635 58.430 275.550 58.430 ;
        RECT 287.880 58.580 303.120 59.240 ;
        POLYGON 287.880 58.580 287.895 58.580 287.895 58.450 ;
        RECT 287.895 58.430 303.120 58.580 ;
        RECT 268.355 58.425 275.635 58.430 ;
        RECT 260.640 58.400 263.820 58.425 ;
        RECT 255.770 58.395 258.050 58.400 ;
        RECT 247.245 58.385 253.355 58.395 ;
        POLYGON 247.195 58.385 247.195 58.370 247.165 58.370 ;
        RECT 247.195 58.370 253.355 58.385 ;
        POLYGON 253.355 58.395 253.415 58.370 253.355 58.370 ;
        POLYGON 255.770 58.395 255.805 58.395 255.805 58.370 ;
        RECT 255.805 58.370 258.050 58.395 ;
        POLYGON 247.165 58.370 247.165 58.340 247.085 58.340 ;
        RECT 247.165 58.340 253.420 58.370 ;
        POLYGON 247.080 58.340 247.080 58.315 247.010 58.315 ;
        RECT 247.080 58.315 253.420 58.340 ;
        POLYGON 247.010 58.315 247.010 58.310 246.995 58.310 ;
        RECT 247.010 58.310 253.420 58.315 ;
        POLYGON 253.420 58.370 253.580 58.310 253.420 58.310 ;
        POLYGON 255.805 58.370 255.815 58.370 255.815 58.365 ;
        RECT 255.815 58.365 258.050 58.370 ;
        POLYGON 255.815 58.365 255.865 58.365 255.865 58.335 ;
        RECT 255.865 58.335 258.050 58.365 ;
        POLYGON 255.865 58.335 255.900 58.335 255.900 58.310 ;
        RECT 255.900 58.325 258.050 58.335 ;
        POLYGON 258.050 58.400 258.135 58.325 258.050 58.325 ;
        POLYGON 260.640 58.400 260.695 58.400 260.695 58.345 ;
        RECT 260.695 58.395 263.820 58.400 ;
        POLYGON 263.820 58.425 263.840 58.395 263.820 58.395 ;
        POLYGON 268.355 58.425 268.370 58.425 268.370 58.395 ;
        RECT 268.370 58.395 275.635 58.425 ;
        RECT 260.695 58.345 263.840 58.395 ;
        POLYGON 260.695 58.345 260.710 58.345 260.710 58.325 ;
        RECT 260.710 58.325 263.840 58.345 ;
        RECT 255.900 58.310 258.135 58.325 ;
        RECT 242.930 58.265 244.845 58.305 ;
        POLYGON 244.845 58.305 244.900 58.305 244.845 58.265 ;
        POLYGON 246.995 58.310 246.995 58.280 246.920 58.280 ;
        RECT 246.995 58.280 253.580 58.310 ;
        POLYGON 246.920 58.280 246.920 58.265 246.885 58.265 ;
        RECT 246.920 58.270 253.580 58.280 ;
        POLYGON 253.580 58.310 253.670 58.270 253.580 58.270 ;
        POLYGON 255.900 58.310 255.960 58.310 255.960 58.270 ;
        RECT 255.960 58.270 258.135 58.310 ;
        RECT 246.920 58.265 253.670 58.270 ;
        RECT 242.930 58.255 244.795 58.265 ;
        POLYGON 242.840 58.255 242.840 58.245 242.825 58.245 ;
        RECT 242.840 58.245 244.795 58.255 ;
        POLYGON 242.825 58.245 242.825 58.190 242.770 58.190 ;
        RECT 242.825 58.235 244.795 58.245 ;
        POLYGON 244.795 58.265 244.840 58.265 244.795 58.235 ;
        POLYGON 246.885 58.265 246.885 58.235 246.820 58.235 ;
        RECT 246.885 58.235 253.670 58.265 ;
        RECT 242.825 58.190 244.740 58.235 ;
        POLYGON 244.740 58.235 244.795 58.235 244.740 58.190 ;
        POLYGON 246.820 58.235 246.820 58.215 246.775 58.215 ;
        RECT 246.820 58.230 253.670 58.235 ;
        POLYGON 253.670 58.270 253.775 58.230 253.670 58.230 ;
        POLYGON 255.960 58.270 256.005 58.270 256.005 58.240 ;
        RECT 256.005 58.240 258.135 58.270 ;
        POLYGON 256.005 58.240 256.010 58.240 256.010 58.235 ;
        RECT 256.010 58.235 258.135 58.240 ;
        POLYGON 256.015 58.235 256.020 58.235 256.020 58.230 ;
        RECT 256.020 58.230 258.135 58.235 ;
        POLYGON 258.135 58.325 258.245 58.230 258.135 58.230 ;
        POLYGON 260.710 58.325 260.795 58.325 260.795 58.230 ;
        RECT 260.795 58.230 263.840 58.325 ;
        RECT 246.820 58.220 253.775 58.230 ;
        POLYGON 253.775 58.230 253.800 58.220 253.775 58.220 ;
        POLYGON 256.020 58.230 256.035 58.230 256.035 58.220 ;
        RECT 256.035 58.220 258.245 58.230 ;
        RECT 246.820 58.215 253.800 58.220 ;
        POLYGON 246.775 58.215 246.775 58.205 246.750 58.205 ;
        RECT 246.775 58.205 253.800 58.215 ;
        POLYGON 246.750 58.205 246.750 58.190 246.720 58.190 ;
        RECT 246.750 58.190 253.800 58.205 ;
        POLYGON 253.800 58.220 253.860 58.190 253.800 58.190 ;
        POLYGON 256.035 58.220 256.075 58.220 256.075 58.190 ;
        RECT 256.075 58.190 258.245 58.220 ;
        POLYGON 258.245 58.230 258.285 58.190 258.245 58.190 ;
        POLYGON 260.795 58.230 260.830 58.230 260.830 58.190 ;
        RECT 260.830 58.190 263.840 58.230 ;
        POLYGON 263.840 58.395 263.980 58.190 263.840 58.190 ;
        POLYGON 268.370 58.395 268.480 58.395 268.480 58.190 ;
        RECT 268.480 58.295 275.635 58.395 ;
        POLYGON 275.635 58.430 275.695 58.295 275.635 58.295 ;
        POLYGON 287.895 58.430 287.910 58.430 287.910 58.320 ;
        RECT 287.910 58.295 303.120 58.430 ;
        RECT 268.480 58.195 275.695 58.295 ;
        POLYGON 275.695 58.295 275.735 58.195 275.695 58.195 ;
        RECT 268.480 58.190 275.735 58.195 ;
        POLYGON 287.910 58.295 287.925 58.295 287.925 58.190 ;
        RECT 287.925 58.190 303.120 58.295 ;
        POLYGON 230.115 58.185 230.115 58.110 230.090 58.110 ;
        RECT 230.115 58.155 234.740 58.190 ;
        POLYGON 234.740 58.190 234.760 58.190 234.740 58.155 ;
        POLYGON 238.105 58.190 238.105 58.155 238.085 58.155 ;
        RECT 238.105 58.155 240.600 58.190 ;
        POLYGON 240.600 58.190 240.630 58.190 240.600 58.155 ;
        POLYGON 242.770 58.190 242.770 58.155 242.730 58.155 ;
        RECT 242.770 58.155 244.625 58.190 ;
        RECT 230.115 58.110 234.715 58.155 ;
        POLYGON 180.925 57.780 181.025 57.780 181.025 57.535 ;
        RECT 181.025 57.525 195.225 57.780 ;
        RECT 169.420 57.490 173.850 57.525 ;
        POLYGON 164.010 57.490 164.045 57.490 164.045 57.445 ;
        RECT 164.045 57.445 166.390 57.490 ;
        RECT 160.370 57.410 162.025 57.445 ;
        POLYGON 162.025 57.445 162.065 57.410 162.025 57.410 ;
        POLYGON 164.045 57.445 164.080 57.445 164.080 57.410 ;
        RECT 164.080 57.410 166.390 57.445 ;
        RECT 160.370 57.365 162.065 57.410 ;
        RECT 151.910 57.345 154.255 57.365 ;
        POLYGON 154.255 57.365 154.375 57.365 154.255 57.345 ;
        POLYGON 156.245 57.365 156.355 57.365 156.355 57.345 ;
        RECT 156.355 57.345 158.550 57.365 ;
        RECT 151.910 57.335 154.190 57.345 ;
        POLYGON 154.190 57.345 154.255 57.345 154.190 57.335 ;
        POLYGON 156.360 57.345 156.385 57.345 156.385 57.340 ;
        RECT 156.385 57.340 158.550 57.345 ;
        POLYGON 156.390 57.340 156.420 57.340 156.420 57.335 ;
        RECT 156.420 57.335 158.550 57.340 ;
        POLYGON 158.550 57.365 158.615 57.335 158.550 57.335 ;
        POLYGON 160.370 57.365 160.415 57.365 160.415 57.335 ;
        RECT 160.415 57.335 162.065 57.365 ;
        RECT 151.910 57.325 154.130 57.335 ;
        POLYGON 154.130 57.335 154.185 57.335 154.130 57.325 ;
        POLYGON 156.420 57.335 156.450 57.335 156.450 57.330 ;
        RECT 156.450 57.330 158.615 57.335 ;
        POLYGON 156.450 57.330 156.475 57.330 156.475 57.325 ;
        RECT 156.475 57.325 158.615 57.330 ;
        RECT 151.910 57.320 154.110 57.325 ;
        POLYGON 154.110 57.325 154.125 57.325 154.110 57.320 ;
        POLYGON 156.475 57.325 156.500 57.325 156.500 57.320 ;
        RECT 156.500 57.320 158.615 57.325 ;
        RECT 151.910 57.315 153.995 57.320 ;
        RECT 148.760 57.280 150.150 57.315 ;
        POLYGON 148.645 57.280 148.645 57.260 148.625 57.260 ;
        RECT 148.645 57.260 150.150 57.280 ;
        RECT 117.310 57.160 146.785 57.260 ;
        POLYGON 146.785 57.260 146.865 57.260 146.785 57.160 ;
        POLYGON 148.625 57.260 148.625 57.160 148.520 57.160 ;
        RECT 148.625 57.255 150.150 57.260 ;
        POLYGON 150.150 57.315 150.230 57.315 150.150 57.255 ;
        POLYGON 151.705 57.315 151.705 57.300 151.675 57.300 ;
        RECT 151.705 57.300 153.995 57.315 ;
        POLYGON 153.995 57.320 154.110 57.320 153.995 57.300 ;
        POLYGON 156.500 57.320 156.620 57.320 156.620 57.300 ;
        RECT 156.620 57.300 158.615 57.320 ;
        POLYGON 151.670 57.300 151.670 57.255 151.585 57.255 ;
        RECT 151.670 57.285 153.915 57.300 ;
        POLYGON 153.915 57.300 153.995 57.300 153.915 57.285 ;
        POLYGON 156.625 57.300 156.690 57.300 156.690 57.285 ;
        RECT 156.690 57.285 158.615 57.300 ;
        RECT 151.670 57.270 153.840 57.285 ;
        POLYGON 153.840 57.285 153.915 57.285 153.840 57.270 ;
        POLYGON 156.690 57.285 156.735 57.285 156.735 57.275 ;
        RECT 156.735 57.275 158.615 57.285 ;
        POLYGON 156.745 57.275 156.765 57.275 156.765 57.270 ;
        RECT 156.765 57.270 158.615 57.275 ;
        RECT 151.670 57.255 153.755 57.270 ;
        RECT 148.625 57.245 150.135 57.255 ;
        POLYGON 150.135 57.255 150.150 57.255 150.135 57.245 ;
        POLYGON 151.585 57.255 151.585 57.245 151.565 57.245 ;
        RECT 151.585 57.245 153.755 57.255 ;
        POLYGON 153.755 57.270 153.840 57.270 153.755 57.245 ;
        POLYGON 156.765 57.270 156.825 57.270 156.825 57.255 ;
        RECT 156.825 57.255 158.615 57.270 ;
        POLYGON 158.615 57.335 158.770 57.255 158.615 57.255 ;
        POLYGON 160.415 57.335 160.445 57.335 160.445 57.315 ;
        RECT 160.445 57.315 162.065 57.335 ;
        POLYGON 160.445 57.315 160.495 57.315 160.495 57.280 ;
        RECT 160.495 57.280 162.065 57.315 ;
        POLYGON 162.065 57.410 162.210 57.280 162.065 57.280 ;
        POLYGON 164.080 57.410 164.105 57.410 164.105 57.385 ;
        RECT 164.105 57.385 166.390 57.410 ;
        POLYGON 164.105 57.385 164.155 57.385 164.155 57.325 ;
        RECT 164.155 57.325 166.390 57.385 ;
        POLYGON 164.155 57.325 164.190 57.325 164.190 57.285 ;
        RECT 164.190 57.310 166.390 57.325 ;
        POLYGON 166.390 57.490 166.515 57.310 166.390 57.310 ;
        POLYGON 169.420 57.490 169.530 57.490 169.530 57.315 ;
        RECT 169.530 57.380 173.850 57.490 ;
        POLYGON 173.850 57.525 173.920 57.380 173.850 57.380 ;
        POLYGON 181.025 57.525 181.085 57.525 181.085 57.390 ;
        RECT 181.085 57.380 195.225 57.525 ;
        RECT 169.530 57.310 173.920 57.380 ;
        RECT 164.190 57.280 166.515 57.310 ;
        POLYGON 160.495 57.280 160.530 57.280 160.530 57.255 ;
        RECT 160.530 57.255 162.210 57.280 ;
        POLYGON 156.830 57.255 156.870 57.255 156.870 57.245 ;
        RECT 156.870 57.245 158.770 57.255 ;
        RECT 148.625 57.160 150.005 57.245 ;
        RECT 117.310 57.085 146.725 57.160 ;
        POLYGON 146.725 57.160 146.785 57.160 146.725 57.085 ;
        POLYGON 148.520 57.160 148.520 57.095 148.455 57.095 ;
        RECT 148.520 57.150 150.005 57.160 ;
        POLYGON 150.005 57.245 150.135 57.245 150.005 57.150 ;
        POLYGON 151.565 57.245 151.565 57.215 151.510 57.215 ;
        RECT 151.565 57.235 153.705 57.245 ;
        POLYGON 153.705 57.245 153.735 57.245 153.705 57.235 ;
        POLYGON 156.870 57.245 156.910 57.245 156.910 57.235 ;
        RECT 156.910 57.235 158.770 57.245 ;
        RECT 151.565 57.215 153.575 57.235 ;
        POLYGON 151.510 57.215 151.510 57.180 151.445 57.180 ;
        RECT 151.510 57.205 153.575 57.215 ;
        POLYGON 153.575 57.235 153.705 57.235 153.575 57.205 ;
        POLYGON 156.910 57.235 156.990 57.235 156.990 57.215 ;
        RECT 156.990 57.225 158.770 57.235 ;
        POLYGON 158.770 57.255 158.825 57.225 158.770 57.225 ;
        POLYGON 160.530 57.255 160.540 57.255 160.540 57.250 ;
        RECT 160.540 57.250 162.210 57.255 ;
        POLYGON 160.540 57.250 160.570 57.250 160.570 57.225 ;
        RECT 160.570 57.225 162.210 57.250 ;
        POLYGON 162.210 57.280 162.275 57.225 162.210 57.225 ;
        POLYGON 164.190 57.280 164.240 57.280 164.240 57.225 ;
        RECT 164.240 57.225 166.515 57.280 ;
        RECT 156.990 57.215 158.825 57.225 ;
        POLYGON 156.990 57.215 157.015 57.215 157.015 57.205 ;
        RECT 157.015 57.205 158.825 57.215 ;
        RECT 151.510 57.180 153.495 57.205 ;
        POLYGON 153.495 57.205 153.575 57.205 153.495 57.180 ;
        POLYGON 157.015 57.205 157.030 57.205 157.030 57.200 ;
        RECT 157.030 57.200 158.825 57.205 ;
        POLYGON 158.825 57.225 158.885 57.200 158.825 57.200 ;
        POLYGON 160.570 57.225 160.605 57.225 160.605 57.200 ;
        RECT 160.605 57.200 162.275 57.225 ;
        POLYGON 157.030 57.200 157.100 57.200 157.100 57.180 ;
        RECT 157.100 57.180 158.885 57.200 ;
        POLYGON 151.445 57.180 151.445 57.150 151.390 57.150 ;
        RECT 151.445 57.150 153.325 57.180 ;
        RECT 148.520 57.095 149.850 57.150 ;
        POLYGON 148.455 57.095 148.455 57.085 148.445 57.085 ;
        RECT 148.455 57.085 149.850 57.095 ;
        RECT 117.310 56.990 146.650 57.085 ;
        POLYGON 146.650 57.085 146.725 57.085 146.650 56.990 ;
        POLYGON 148.445 57.085 148.445 57.030 148.390 57.030 ;
        RECT 148.445 57.035 149.850 57.085 ;
        POLYGON 149.850 57.150 150.005 57.150 149.850 57.035 ;
        POLYGON 151.390 57.150 151.390 57.095 151.285 57.095 ;
        RECT 151.390 57.135 153.325 57.150 ;
        POLYGON 153.325 57.180 153.480 57.180 153.325 57.135 ;
        POLYGON 157.100 57.180 157.155 57.180 157.155 57.165 ;
        RECT 157.155 57.165 158.885 57.180 ;
        POLYGON 157.155 57.165 157.250 57.165 157.250 57.140 ;
        RECT 157.250 57.155 158.885 57.165 ;
        POLYGON 158.885 57.200 158.965 57.155 158.885 57.155 ;
        POLYGON 160.605 57.200 160.615 57.200 160.615 57.195 ;
        RECT 160.615 57.195 162.275 57.200 ;
        POLYGON 160.615 57.195 160.670 57.195 160.670 57.155 ;
        RECT 160.670 57.155 162.275 57.195 ;
        RECT 157.250 57.140 158.965 57.155 ;
        POLYGON 157.250 57.140 157.265 57.140 157.265 57.135 ;
        RECT 157.265 57.135 158.965 57.140 ;
        RECT 151.390 57.130 153.305 57.135 ;
        POLYGON 153.305 57.135 153.320 57.135 153.305 57.130 ;
        POLYGON 157.265 57.135 157.280 57.135 157.280 57.130 ;
        RECT 157.280 57.130 158.965 57.135 ;
        RECT 151.390 57.105 153.225 57.130 ;
        POLYGON 153.225 57.130 153.305 57.130 153.225 57.105 ;
        POLYGON 157.280 57.130 157.310 57.130 157.310 57.120 ;
        RECT 157.310 57.125 158.965 57.130 ;
        POLYGON 158.965 57.155 159.025 57.125 158.965 57.125 ;
        POLYGON 160.670 57.155 160.695 57.155 160.695 57.140 ;
        RECT 160.695 57.140 162.275 57.155 ;
        POLYGON 160.695 57.140 160.710 57.140 160.710 57.125 ;
        RECT 160.710 57.125 162.275 57.140 ;
        RECT 157.310 57.120 159.025 57.125 ;
        POLYGON 157.315 57.120 157.355 57.120 157.355 57.105 ;
        RECT 157.355 57.105 159.025 57.120 ;
        RECT 151.390 57.095 153.090 57.105 ;
        POLYGON 151.285 57.095 151.285 57.060 151.225 57.060 ;
        RECT 151.285 57.060 153.090 57.095 ;
        POLYGON 153.090 57.105 153.225 57.105 153.090 57.060 ;
        POLYGON 157.355 57.105 157.425 57.105 157.425 57.080 ;
        RECT 157.425 57.080 159.025 57.105 ;
        POLYGON 157.425 57.080 157.485 57.080 157.485 57.060 ;
        RECT 157.485 57.060 159.025 57.080 ;
        POLYGON 151.225 57.060 151.225 57.040 151.195 57.040 ;
        RECT 151.225 57.045 153.040 57.060 ;
        POLYGON 153.040 57.060 153.090 57.060 153.040 57.045 ;
        POLYGON 157.485 57.060 157.530 57.060 157.530 57.045 ;
        RECT 157.530 57.050 159.025 57.060 ;
        POLYGON 159.025 57.125 159.155 57.050 159.025 57.050 ;
        POLYGON 160.710 57.125 160.810 57.125 160.810 57.050 ;
        RECT 160.810 57.065 162.275 57.125 ;
        POLYGON 162.275 57.225 162.440 57.065 162.275 57.065 ;
        POLYGON 164.240 57.225 164.260 57.225 164.260 57.205 ;
        RECT 164.260 57.205 166.515 57.225 ;
        POLYGON 164.260 57.205 164.365 57.205 164.365 57.085 ;
        RECT 164.365 57.095 166.515 57.205 ;
        POLYGON 166.515 57.310 166.665 57.095 166.515 57.095 ;
        POLYGON 169.530 57.310 169.540 57.310 169.540 57.300 ;
        RECT 169.540 57.300 173.920 57.310 ;
        POLYGON 169.540 57.300 169.645 57.300 169.645 57.100 ;
        RECT 169.645 57.155 173.920 57.300 ;
        POLYGON 173.920 57.380 174.025 57.155 173.920 57.155 ;
        POLYGON 181.085 57.380 181.180 57.380 181.180 57.160 ;
        RECT 181.180 57.155 195.225 57.380 ;
        RECT 169.645 57.095 174.025 57.155 ;
        RECT 164.365 57.085 166.665 57.095 ;
        POLYGON 164.365 57.085 164.385 57.085 164.385 57.065 ;
        RECT 164.385 57.065 166.665 57.085 ;
        RECT 160.810 57.050 162.440 57.065 ;
        RECT 157.530 57.045 159.155 57.050 ;
        RECT 151.225 57.040 152.975 57.045 ;
        POLYGON 151.195 57.040 151.195 57.035 151.185 57.035 ;
        RECT 151.195 57.035 152.975 57.040 ;
        RECT 148.445 57.030 149.780 57.035 ;
        POLYGON 148.390 57.030 148.390 56.995 148.360 56.995 ;
        RECT 148.390 56.995 149.780 57.030 ;
        POLYGON 148.360 56.995 148.360 56.990 148.355 56.990 ;
        RECT 148.360 56.990 149.780 56.995 ;
        RECT 117.310 56.920 146.595 56.990 ;
        POLYGON 146.595 56.990 146.650 56.990 146.595 56.920 ;
        POLYGON 148.355 56.990 148.355 56.920 148.290 56.920 ;
        RECT 148.355 56.980 149.780 56.990 ;
        POLYGON 149.780 57.035 149.850 57.035 149.780 56.980 ;
        POLYGON 151.185 57.035 151.185 56.980 151.100 56.980 ;
        RECT 151.185 57.020 152.975 57.035 ;
        POLYGON 152.975 57.045 153.040 57.045 152.975 57.020 ;
        POLYGON 157.530 57.045 157.590 57.045 157.590 57.025 ;
        RECT 157.590 57.025 159.155 57.045 ;
        POLYGON 157.590 57.025 157.600 57.025 157.600 57.020 ;
        RECT 157.600 57.020 159.155 57.025 ;
        RECT 151.185 56.995 152.900 57.020 ;
        POLYGON 152.900 57.020 152.970 57.020 152.900 56.995 ;
        POLYGON 157.600 57.020 157.665 57.020 157.665 56.995 ;
        RECT 157.665 56.995 159.155 57.020 ;
        RECT 151.185 56.980 152.770 56.995 ;
        RECT 148.355 56.930 149.715 56.980 ;
        POLYGON 149.715 56.980 149.780 56.980 149.715 56.930 ;
        POLYGON 151.100 56.980 151.100 56.950 151.050 56.950 ;
        RECT 151.100 56.950 152.770 56.980 ;
        POLYGON 152.770 56.995 152.900 56.995 152.770 56.950 ;
        POLYGON 157.665 56.995 157.690 56.995 157.690 56.985 ;
        RECT 157.690 56.985 159.155 56.995 ;
        POLYGON 157.700 56.985 157.755 56.985 157.755 56.965 ;
        RECT 157.755 56.980 159.155 56.985 ;
        POLYGON 159.155 57.050 159.275 56.980 159.155 56.980 ;
        POLYGON 160.810 57.050 160.860 57.050 160.860 57.015 ;
        RECT 160.860 57.015 162.440 57.050 ;
        POLYGON 160.860 57.015 160.905 57.015 160.905 56.980 ;
        RECT 160.905 56.980 162.440 57.015 ;
        RECT 157.755 56.970 159.275 56.980 ;
        POLYGON 159.275 56.980 159.290 56.970 159.275 56.970 ;
        POLYGON 160.905 56.980 160.915 56.980 160.915 56.970 ;
        RECT 160.915 56.970 162.440 56.980 ;
        RECT 157.755 56.965 159.290 56.970 ;
        POLYGON 157.755 56.965 157.790 56.965 157.790 56.950 ;
        RECT 157.790 56.950 159.290 56.965 ;
        POLYGON 151.050 56.950 151.050 56.930 151.015 56.930 ;
        RECT 151.050 56.930 152.720 56.950 ;
        RECT 148.355 56.920 149.560 56.930 ;
        RECT 117.310 56.810 146.515 56.920 ;
        POLYGON 146.515 56.920 146.595 56.920 146.515 56.810 ;
        POLYGON 148.290 56.920 148.290 56.810 148.185 56.810 ;
        RECT 148.290 56.810 149.560 56.920 ;
        RECT 117.310 56.715 146.445 56.810 ;
        POLYGON 146.445 56.810 146.515 56.810 146.445 56.715 ;
        POLYGON 148.185 56.810 148.185 56.755 148.130 56.755 ;
        RECT 148.185 56.800 149.560 56.810 ;
        POLYGON 149.560 56.930 149.715 56.930 149.560 56.800 ;
        POLYGON 151.015 56.930 151.015 56.890 150.950 56.890 ;
        RECT 151.015 56.925 152.720 56.930 ;
        POLYGON 152.720 56.950 152.770 56.950 152.720 56.925 ;
        POLYGON 157.790 56.950 157.845 56.950 157.845 56.925 ;
        RECT 157.845 56.925 159.290 56.950 ;
        RECT 151.015 56.915 152.690 56.925 ;
        POLYGON 152.690 56.925 152.720 56.925 152.690 56.915 ;
        POLYGON 157.845 56.925 157.860 56.925 157.860 56.920 ;
        RECT 157.860 56.920 159.290 56.925 ;
        POLYGON 159.290 56.970 159.375 56.920 159.290 56.920 ;
        POLYGON 160.915 56.970 160.940 56.970 160.940 56.950 ;
        RECT 160.940 56.950 162.440 56.970 ;
        POLYGON 160.940 56.950 160.975 56.950 160.975 56.920 ;
        RECT 160.975 56.920 162.440 56.950 ;
        POLYGON 157.865 56.920 157.875 56.920 157.875 56.915 ;
        RECT 157.875 56.915 159.375 56.920 ;
        RECT 151.015 56.890 152.505 56.915 ;
        POLYGON 150.950 56.890 150.950 56.865 150.910 56.865 ;
        RECT 150.950 56.865 152.505 56.890 ;
        POLYGON 150.910 56.865 150.910 56.830 150.860 56.830 ;
        RECT 150.910 56.840 152.505 56.865 ;
        POLYGON 152.505 56.915 152.690 56.915 152.505 56.840 ;
        POLYGON 157.875 56.915 157.955 56.915 157.955 56.880 ;
        RECT 157.955 56.895 159.375 56.915 ;
        POLYGON 159.375 56.920 159.420 56.895 159.375 56.895 ;
        POLYGON 160.975 56.920 161.005 56.920 161.005 56.895 ;
        RECT 161.005 56.895 162.440 56.920 ;
        POLYGON 162.440 57.065 162.610 56.895 162.440 56.895 ;
        POLYGON 164.385 57.065 164.435 57.065 164.435 57.000 ;
        RECT 164.435 57.000 166.665 57.065 ;
        POLYGON 164.435 57.000 164.495 57.000 164.495 56.930 ;
        RECT 164.495 56.930 166.665 57.000 ;
        POLYGON 164.495 56.930 164.520 56.930 164.520 56.895 ;
        RECT 164.520 56.895 166.665 56.930 ;
        RECT 157.955 56.880 159.420 56.895 ;
        POLYGON 157.960 56.880 158.005 56.880 158.005 56.860 ;
        RECT 158.005 56.860 159.420 56.880 ;
        POLYGON 158.005 56.860 158.045 56.860 158.045 56.840 ;
        RECT 158.045 56.840 159.420 56.860 ;
        RECT 150.910 56.830 152.485 56.840 ;
        POLYGON 152.485 56.840 152.505 56.840 152.485 56.835 ;
        POLYGON 158.045 56.840 158.055 56.840 158.055 56.835 ;
        RECT 158.055 56.835 159.420 56.840 ;
        POLYGON 150.860 56.830 150.860 56.800 150.815 56.800 ;
        RECT 150.860 56.825 152.470 56.830 ;
        POLYGON 152.470 56.830 152.485 56.830 152.470 56.825 ;
        POLYGON 158.055 56.835 158.075 56.835 158.075 56.825 ;
        RECT 158.075 56.830 159.420 56.835 ;
        POLYGON 159.420 56.895 159.515 56.830 159.420 56.830 ;
        POLYGON 161.005 56.895 161.085 56.895 161.085 56.830 ;
        RECT 161.085 56.830 162.610 56.895 ;
        RECT 158.075 56.825 159.515 56.830 ;
        RECT 150.860 56.800 152.310 56.825 ;
        RECT 148.185 56.775 149.525 56.800 ;
        POLYGON 149.525 56.800 149.560 56.800 149.525 56.775 ;
        POLYGON 150.815 56.800 150.815 56.775 150.780 56.775 ;
        RECT 150.815 56.775 152.310 56.800 ;
        RECT 148.185 56.755 149.435 56.775 ;
        POLYGON 148.130 56.755 148.130 56.715 148.095 56.715 ;
        RECT 148.130 56.715 149.435 56.755 ;
        RECT 117.310 56.660 146.410 56.715 ;
        POLYGON 146.410 56.715 146.445 56.715 146.410 56.660 ;
        POLYGON 148.095 56.715 148.095 56.705 148.085 56.705 ;
        RECT 148.095 56.705 149.435 56.715 ;
        POLYGON 148.085 56.705 148.085 56.660 148.045 56.660 ;
        RECT 148.085 56.690 149.435 56.705 ;
        POLYGON 149.435 56.775 149.525 56.775 149.435 56.690 ;
        POLYGON 150.780 56.775 150.780 56.725 150.705 56.725 ;
        RECT 150.780 56.755 152.310 56.775 ;
        POLYGON 152.310 56.825 152.470 56.825 152.310 56.755 ;
        POLYGON 158.075 56.825 158.125 56.825 158.125 56.800 ;
        RECT 158.125 56.800 159.515 56.825 ;
        POLYGON 158.130 56.800 158.140 56.800 158.140 56.795 ;
        RECT 158.140 56.795 159.515 56.800 ;
        POLYGON 155.150 56.795 155.150 56.790 155.065 56.790 ;
        RECT 155.150 56.790 155.300 56.795 ;
        POLYGON 155.300 56.795 155.485 56.790 155.300 56.790 ;
        POLYGON 158.140 56.795 158.150 56.795 158.150 56.790 ;
        RECT 158.150 56.790 159.515 56.795 ;
        POLYGON 155.000 56.790 155.000 56.785 154.905 56.785 ;
        RECT 155.000 56.785 155.565 56.790 ;
        POLYGON 154.900 56.785 154.900 56.780 154.785 56.780 ;
        RECT 154.900 56.780 155.565 56.785 ;
        POLYGON 155.565 56.790 155.690 56.780 155.565 56.780 ;
        POLYGON 158.150 56.790 158.175 56.790 158.175 56.780 ;
        RECT 158.175 56.780 159.515 56.790 ;
        POLYGON 154.785 56.780 154.785 56.775 154.775 56.775 ;
        RECT 154.785 56.775 155.695 56.780 ;
        POLYGON 155.695 56.780 155.820 56.775 155.695 56.775 ;
        POLYGON 158.175 56.780 158.185 56.780 158.185 56.775 ;
        RECT 158.185 56.775 159.515 56.780 ;
        POLYGON 154.770 56.775 154.770 56.765 154.640 56.765 ;
        RECT 154.770 56.770 155.830 56.775 ;
        POLYGON 155.830 56.775 155.850 56.770 155.830 56.770 ;
        POLYGON 158.185 56.775 158.200 56.775 158.200 56.770 ;
        RECT 158.200 56.770 159.515 56.775 ;
        RECT 154.770 56.765 155.850 56.770 ;
        POLYGON 154.625 56.765 154.625 56.760 154.565 56.760 ;
        RECT 154.625 56.760 155.850 56.765 ;
        POLYGON 155.850 56.770 155.940 56.760 155.850 56.760 ;
        POLYGON 158.200 56.770 158.220 56.770 158.220 56.760 ;
        RECT 158.220 56.760 159.515 56.770 ;
        POLYGON 154.565 56.760 154.565 56.755 154.515 56.755 ;
        RECT 154.565 56.755 155.955 56.760 ;
        RECT 150.780 56.725 152.235 56.755 ;
        POLYGON 152.235 56.755 152.310 56.755 152.235 56.725 ;
        POLYGON 154.515 56.755 154.515 56.735 154.375 56.735 ;
        RECT 154.515 56.745 155.955 56.755 ;
        POLYGON 155.955 56.760 156.085 56.745 155.955 56.745 ;
        POLYGON 158.220 56.760 158.235 56.760 158.235 56.755 ;
        RECT 158.235 56.755 159.515 56.760 ;
        POLYGON 158.235 56.755 158.255 56.755 158.255 56.745 ;
        RECT 158.255 56.745 159.515 56.755 ;
        RECT 154.515 56.740 156.095 56.745 ;
        POLYGON 156.095 56.745 156.155 56.740 156.095 56.740 ;
        POLYGON 158.255 56.745 158.260 56.745 158.260 56.740 ;
        RECT 158.260 56.740 159.515 56.745 ;
        RECT 154.515 56.735 156.155 56.740 ;
        POLYGON 154.345 56.735 154.345 56.725 154.285 56.725 ;
        RECT 154.345 56.730 156.155 56.735 ;
        POLYGON 156.155 56.740 156.215 56.730 156.155 56.730 ;
        POLYGON 158.260 56.740 158.280 56.740 158.280 56.730 ;
        RECT 158.280 56.730 159.515 56.740 ;
        RECT 154.345 56.725 156.220 56.730 ;
        POLYGON 150.705 56.725 150.705 56.690 150.655 56.690 ;
        RECT 150.705 56.715 152.220 56.725 ;
        POLYGON 152.220 56.725 152.235 56.725 152.220 56.715 ;
        POLYGON 154.285 56.725 154.285 56.720 154.255 56.720 ;
        RECT 154.285 56.720 156.220 56.725 ;
        POLYGON 154.250 56.720 154.250 56.715 154.220 56.715 ;
        RECT 154.250 56.715 156.220 56.720 ;
        RECT 150.705 56.690 152.075 56.715 ;
        RECT 148.085 56.660 149.345 56.690 ;
        RECT 117.310 56.435 146.320 56.660 ;
        POLYGON 146.320 56.660 146.410 56.660 146.320 56.525 ;
        POLYGON 148.045 56.660 148.045 56.605 147.995 56.605 ;
        RECT 148.045 56.615 149.345 56.660 ;
        POLYGON 149.345 56.690 149.435 56.690 149.345 56.615 ;
        POLYGON 150.655 56.690 150.655 56.650 150.595 56.650 ;
        RECT 150.655 56.650 152.075 56.690 ;
        POLYGON 150.590 56.650 150.590 56.615 150.545 56.615 ;
        RECT 150.590 56.645 152.075 56.650 ;
        POLYGON 152.075 56.715 152.220 56.715 152.075 56.645 ;
        POLYGON 154.220 56.715 154.220 56.710 154.185 56.710 ;
        RECT 154.220 56.710 156.220 56.715 ;
        POLYGON 156.220 56.730 156.360 56.710 156.220 56.710 ;
        POLYGON 158.280 56.730 158.320 56.730 158.320 56.710 ;
        RECT 158.320 56.710 159.515 56.730 ;
        POLYGON 154.185 56.710 154.185 56.700 154.130 56.700 ;
        RECT 154.185 56.705 156.360 56.710 ;
        POLYGON 156.360 56.710 156.385 56.705 156.360 56.705 ;
        POLYGON 158.320 56.710 158.325 56.710 158.325 56.705 ;
        RECT 158.325 56.705 159.515 56.710 ;
        RECT 154.185 56.700 156.390 56.705 ;
        POLYGON 154.105 56.700 154.105 56.680 153.995 56.680 ;
        RECT 154.105 56.695 156.390 56.700 ;
        POLYGON 156.390 56.705 156.450 56.695 156.390 56.695 ;
        POLYGON 158.325 56.705 158.345 56.705 158.345 56.695 ;
        RECT 158.345 56.695 159.515 56.705 ;
        RECT 154.105 56.690 156.450 56.695 ;
        POLYGON 156.450 56.695 156.475 56.690 156.450 56.690 ;
        POLYGON 158.345 56.695 158.355 56.695 158.355 56.690 ;
        RECT 158.355 56.690 159.515 56.695 ;
        RECT 154.105 56.680 156.475 56.690 ;
        POLYGON 153.995 56.680 153.995 56.665 153.915 56.665 ;
        RECT 153.995 56.665 156.475 56.680 ;
        POLYGON 156.475 56.690 156.625 56.665 156.475 56.665 ;
        POLYGON 158.355 56.690 158.405 56.690 158.405 56.665 ;
        RECT 158.405 56.680 159.515 56.690 ;
        POLYGON 159.515 56.830 159.740 56.680 159.515 56.680 ;
        POLYGON 161.085 56.830 161.180 56.830 161.180 56.755 ;
        RECT 161.180 56.755 162.610 56.830 ;
        POLYGON 161.180 56.755 161.210 56.755 161.210 56.725 ;
        RECT 161.210 56.725 162.610 56.755 ;
        POLYGON 161.210 56.725 161.240 56.725 161.240 56.700 ;
        RECT 161.240 56.705 162.610 56.725 ;
        POLYGON 162.610 56.895 162.790 56.705 162.610 56.705 ;
        POLYGON 164.520 56.895 164.595 56.895 164.595 56.805 ;
        RECT 164.595 56.860 166.665 56.895 ;
        POLYGON 166.665 57.095 166.825 56.860 166.665 56.860 ;
        POLYGON 169.645 57.095 169.690 57.095 169.690 57.015 ;
        RECT 169.690 57.015 174.025 57.095 ;
        POLYGON 169.690 57.015 169.770 57.015 169.770 56.865 ;
        RECT 169.770 56.860 174.025 57.015 ;
        RECT 164.595 56.810 166.825 56.860 ;
        POLYGON 166.825 56.860 166.855 56.810 166.825 56.810 ;
        POLYGON 169.770 56.860 169.800 56.860 169.800 56.810 ;
        RECT 169.800 56.810 174.025 56.860 ;
        RECT 164.595 56.805 166.855 56.810 ;
        POLYGON 164.595 56.805 164.615 56.805 164.615 56.775 ;
        RECT 164.615 56.775 166.855 56.805 ;
        POLYGON 164.615 56.775 164.665 56.775 164.665 56.705 ;
        RECT 164.665 56.705 166.855 56.775 ;
        RECT 161.240 56.700 162.790 56.705 ;
        POLYGON 161.240 56.700 161.260 56.700 161.260 56.680 ;
        RECT 161.260 56.680 162.790 56.700 ;
        RECT 158.405 56.675 159.740 56.680 ;
        POLYGON 159.740 56.680 159.750 56.675 159.740 56.675 ;
        POLYGON 161.260 56.680 161.265 56.680 161.265 56.675 ;
        RECT 161.265 56.675 162.790 56.680 ;
        RECT 158.405 56.665 159.750 56.675 ;
        POLYGON 153.915 56.665 153.915 56.645 153.840 56.645 ;
        RECT 153.915 56.645 156.625 56.665 ;
        RECT 150.590 56.615 151.975 56.645 ;
        RECT 148.045 56.605 149.295 56.615 ;
        POLYGON 147.995 56.600 147.995 56.555 147.955 56.555 ;
        RECT 147.995 56.565 149.295 56.605 ;
        POLYGON 149.295 56.615 149.345 56.615 149.295 56.565 ;
        POLYGON 150.545 56.615 150.545 56.580 150.495 56.580 ;
        RECT 150.545 56.600 151.975 56.615 ;
        POLYGON 151.975 56.645 152.075 56.645 151.975 56.600 ;
        POLYGON 153.840 56.645 153.840 56.630 153.750 56.630 ;
        RECT 153.840 56.640 156.625 56.645 ;
        POLYGON 156.625 56.665 156.735 56.640 156.625 56.640 ;
        POLYGON 158.405 56.665 158.455 56.665 158.455 56.640 ;
        RECT 158.455 56.660 159.750 56.665 ;
        POLYGON 159.750 56.675 159.775 56.660 159.750 56.660 ;
        POLYGON 161.265 56.675 161.280 56.675 161.280 56.660 ;
        RECT 161.280 56.665 162.790 56.675 ;
        POLYGON 162.790 56.705 162.825 56.665 162.790 56.665 ;
        POLYGON 164.665 56.705 164.690 56.705 164.690 56.675 ;
        RECT 164.690 56.695 166.855 56.705 ;
        POLYGON 166.855 56.810 166.930 56.695 166.855 56.695 ;
        POLYGON 169.800 56.810 169.860 56.810 169.860 56.700 ;
        RECT 169.860 56.745 174.025 56.810 ;
        POLYGON 174.025 57.155 174.220 56.745 174.025 56.745 ;
        POLYGON 181.180 57.155 181.215 57.155 181.215 57.075 ;
        RECT 181.215 57.130 195.225 57.155 ;
        POLYGON 195.225 57.930 195.525 57.130 195.225 57.130 ;
        POLYGON 206.230 57.790 206.230 57.130 206.225 57.130 ;
        RECT 206.230 57.505 222.360 58.100 ;
        POLYGON 222.360 58.100 222.435 58.100 222.360 57.515 ;
        POLYGON 230.090 58.100 230.090 58.090 230.085 58.090 ;
        RECT 230.090 58.095 234.715 58.110 ;
        POLYGON 234.715 58.155 234.740 58.155 234.715 58.100 ;
        POLYGON 238.085 58.155 238.085 58.105 238.055 58.105 ;
        RECT 238.085 58.105 240.555 58.155 ;
        RECT 238.055 58.100 240.555 58.105 ;
        POLYGON 240.555 58.155 240.600 58.155 240.555 58.100 ;
        POLYGON 242.730 58.155 242.730 58.100 242.675 58.100 ;
        RECT 242.730 58.100 244.625 58.155 ;
        POLYGON 244.625 58.190 244.740 58.190 244.625 58.100 ;
        POLYGON 246.720 58.190 246.720 58.175 246.685 58.175 ;
        RECT 246.720 58.175 253.860 58.190 ;
        POLYGON 253.860 58.190 253.895 58.175 253.860 58.175 ;
        POLYGON 256.075 58.190 256.100 58.190 256.100 58.175 ;
        RECT 256.100 58.175 258.285 58.190 ;
        POLYGON 246.685 58.175 246.685 58.110 246.545 58.110 ;
        RECT 246.685 58.160 253.900 58.175 ;
        POLYGON 253.900 58.175 253.925 58.160 253.900 58.160 ;
        POLYGON 256.100 58.175 256.120 58.175 256.120 58.160 ;
        RECT 256.120 58.160 258.285 58.175 ;
        RECT 246.685 58.120 253.925 58.160 ;
        POLYGON 253.925 58.160 254.015 58.120 253.925 58.120 ;
        POLYGON 256.120 58.160 256.175 58.160 256.175 58.120 ;
        RECT 256.175 58.120 258.285 58.160 ;
        RECT 246.685 58.115 254.015 58.120 ;
        POLYGON 254.015 58.120 254.030 58.115 254.015 58.115 ;
        POLYGON 256.175 58.120 256.185 58.120 256.185 58.115 ;
        RECT 256.185 58.115 258.285 58.120 ;
        RECT 246.685 58.110 254.030 58.115 ;
        POLYGON 246.540 58.110 246.540 58.105 246.535 58.105 ;
        RECT 246.540 58.105 254.030 58.110 ;
        POLYGON 246.535 58.105 246.535 58.100 246.525 58.100 ;
        RECT 246.535 58.100 254.030 58.105 ;
        POLYGON 254.030 58.115 254.055 58.100 254.030 58.100 ;
        POLYGON 256.185 58.115 256.200 58.115 256.200 58.105 ;
        RECT 256.200 58.105 258.285 58.115 ;
        POLYGON 256.200 58.105 256.205 58.105 256.205 58.100 ;
        RECT 256.205 58.100 258.285 58.105 ;
        POLYGON 258.285 58.190 258.385 58.100 258.285 58.100 ;
        POLYGON 260.830 58.190 260.835 58.190 260.835 58.185 ;
        RECT 260.835 58.185 263.980 58.190 ;
        POLYGON 260.835 58.185 260.850 58.185 260.850 58.165 ;
        RECT 260.850 58.165 263.980 58.185 ;
        POLYGON 260.850 58.165 260.900 58.165 260.900 58.100 ;
        RECT 260.900 58.100 263.980 58.165 ;
        POLYGON 263.980 58.190 264.040 58.100 263.980 58.100 ;
        POLYGON 268.480 58.190 268.530 58.190 268.530 58.100 ;
        RECT 268.530 58.100 275.735 58.190 ;
        POLYGON 275.735 58.190 275.775 58.100 275.735 58.100 ;
        POLYGON 287.925 58.190 287.935 58.190 287.935 58.100 ;
        RECT 230.090 58.090 234.570 58.095 ;
        POLYGON 230.085 58.090 230.085 57.870 230.025 57.870 ;
        RECT 230.085 57.870 234.570 58.090 ;
        POLYGON 230.025 57.870 230.025 57.520 229.935 57.520 ;
        RECT 230.025 57.755 234.570 57.870 ;
        POLYGON 234.570 58.095 234.715 58.095 234.570 57.755 ;
        POLYGON 238.055 58.100 238.055 57.755 237.850 57.755 ;
        RECT 238.055 58.005 240.480 58.100 ;
        POLYGON 240.480 58.100 240.555 58.100 240.480 58.005 ;
        POLYGON 242.675 58.100 242.675 58.015 242.585 58.015 ;
        RECT 242.675 58.070 244.590 58.100 ;
        POLYGON 244.590 58.100 244.625 58.100 244.590 58.070 ;
        POLYGON 246.525 58.100 246.525 58.070 246.460 58.070 ;
        RECT 246.525 58.090 254.055 58.100 ;
        RECT 246.525 58.085 249.915 58.090 ;
        POLYGON 249.915 58.090 250.050 58.090 249.915 58.085 ;
        POLYGON 250.220 58.090 250.345 58.090 250.345 58.085 ;
        RECT 250.345 58.085 254.055 58.090 ;
        RECT 246.525 58.080 249.650 58.085 ;
        POLYGON 249.650 58.085 249.725 58.085 249.650 58.080 ;
        POLYGON 250.465 58.085 250.530 58.085 250.530 58.080 ;
        RECT 250.530 58.080 254.055 58.085 ;
        RECT 246.525 58.070 249.405 58.080 ;
        RECT 242.675 58.015 244.450 58.070 ;
        POLYGON 242.585 58.015 242.585 58.005 242.575 58.005 ;
        RECT 242.585 58.005 244.450 58.015 ;
        RECT 238.055 57.975 240.460 58.005 ;
        POLYGON 240.460 58.005 240.480 58.005 240.460 57.975 ;
        POLYGON 242.575 58.005 242.575 57.975 242.545 57.975 ;
        RECT 242.575 57.975 244.450 58.005 ;
        RECT 238.055 57.805 240.335 57.975 ;
        POLYGON 240.335 57.975 240.460 57.975 240.335 57.805 ;
        POLYGON 242.545 57.975 242.545 57.870 242.440 57.870 ;
        RECT 242.545 57.965 244.450 57.975 ;
        POLYGON 244.450 58.070 244.590 58.070 244.450 57.965 ;
        POLYGON 246.460 58.070 246.460 57.990 246.310 57.990 ;
        RECT 246.460 58.065 249.405 58.070 ;
        POLYGON 249.405 58.080 249.645 58.080 249.405 58.065 ;
        POLYGON 250.530 58.080 250.665 58.080 250.665 58.070 ;
        RECT 250.665 58.070 254.055 58.080 ;
        POLYGON 250.705 58.070 250.785 58.070 250.785 58.065 ;
        RECT 250.785 58.065 254.055 58.070 ;
        RECT 246.460 58.060 249.385 58.065 ;
        POLYGON 249.385 58.065 249.405 58.065 249.385 58.060 ;
        POLYGON 250.785 58.065 250.865 58.065 250.865 58.060 ;
        RECT 250.865 58.060 254.055 58.065 ;
        RECT 246.460 58.055 249.300 58.060 ;
        POLYGON 249.300 58.060 249.380 58.060 249.300 58.055 ;
        POLYGON 250.865 58.060 250.905 58.060 250.905 58.055 ;
        RECT 250.905 58.055 254.055 58.060 ;
        RECT 246.460 58.035 249.120 58.055 ;
        POLYGON 249.120 58.055 249.300 58.055 249.120 58.035 ;
        POLYGON 250.915 58.055 250.955 58.055 250.955 58.050 ;
        RECT 250.955 58.050 254.055 58.055 ;
        POLYGON 250.965 58.050 251.135 58.050 251.135 58.035 ;
        RECT 251.135 58.035 254.055 58.050 ;
        POLYGON 254.055 58.100 254.185 58.035 254.055 58.035 ;
        POLYGON 256.205 58.100 256.215 58.100 256.215 58.090 ;
        RECT 256.215 58.090 258.385 58.100 ;
        POLYGON 256.215 58.090 256.265 58.090 256.265 58.055 ;
        RECT 256.265 58.080 258.385 58.090 ;
        POLYGON 258.385 58.100 258.410 58.080 258.385 58.080 ;
        POLYGON 260.900 58.100 260.920 58.100 260.920 58.080 ;
        RECT 256.265 58.075 258.410 58.080 ;
        POLYGON 258.410 58.080 258.415 58.075 258.410 58.075 ;
        RECT 260.920 58.075 264.040 58.100 ;
        RECT 256.265 58.055 258.415 58.075 ;
        POLYGON 256.265 58.055 256.285 58.055 256.285 58.035 ;
        RECT 256.285 58.035 258.415 58.055 ;
        RECT 246.460 58.030 249.095 58.035 ;
        POLYGON 249.095 58.035 249.120 58.035 249.095 58.030 ;
        POLYGON 251.135 58.035 251.175 58.035 251.175 58.030 ;
        RECT 251.175 58.030 254.185 58.035 ;
        RECT 246.460 58.000 248.875 58.030 ;
        POLYGON 248.875 58.030 249.095 58.030 248.875 58.000 ;
        POLYGON 251.175 58.030 251.220 58.030 251.220 58.025 ;
        RECT 251.220 58.025 254.185 58.030 ;
        POLYGON 251.250 58.025 251.425 58.025 251.425 58.000 ;
        RECT 251.425 58.015 254.185 58.025 ;
        POLYGON 254.185 58.035 254.220 58.015 254.185 58.015 ;
        POLYGON 256.285 58.035 256.315 58.035 256.315 58.015 ;
        RECT 256.315 58.015 258.415 58.035 ;
        RECT 251.425 58.000 254.230 58.015 ;
        RECT 246.460 57.995 248.845 58.000 ;
        POLYGON 248.845 58.000 248.850 58.000 248.845 57.995 ;
        POLYGON 251.425 58.000 251.450 58.000 251.450 57.995 ;
        RECT 251.450 57.995 254.230 58.000 ;
        RECT 246.460 57.990 248.785 57.995 ;
        POLYGON 248.785 57.995 248.840 57.995 248.785 57.990 ;
        POLYGON 251.450 57.995 251.480 57.995 251.480 57.990 ;
        RECT 251.480 57.990 254.230 57.995 ;
        POLYGON 246.310 57.990 246.310 57.965 246.260 57.965 ;
        RECT 246.310 57.965 248.585 57.990 ;
        RECT 242.545 57.945 244.425 57.965 ;
        POLYGON 244.425 57.965 244.450 57.965 244.425 57.945 ;
        POLYGON 246.260 57.965 246.260 57.960 246.250 57.960 ;
        RECT 246.260 57.960 248.585 57.965 ;
        POLYGON 246.245 57.960 246.245 57.955 246.240 57.955 ;
        RECT 246.245 57.955 248.585 57.960 ;
        POLYGON 246.235 57.955 246.235 57.945 246.215 57.945 ;
        RECT 246.235 57.950 248.585 57.955 ;
        POLYGON 248.585 57.990 248.785 57.990 248.585 57.950 ;
        POLYGON 251.485 57.990 251.605 57.990 251.605 57.975 ;
        RECT 251.605 57.985 254.230 57.990 ;
        POLYGON 254.230 58.015 254.280 57.985 254.230 57.985 ;
        POLYGON 256.315 58.015 256.355 58.015 256.355 57.985 ;
        RECT 256.355 57.985 258.415 58.015 ;
        RECT 251.605 57.975 254.280 57.985 ;
        POLYGON 251.605 57.975 251.625 57.975 251.625 57.970 ;
        RECT 251.625 57.970 254.280 57.975 ;
        POLYGON 251.625 57.970 251.740 57.970 251.740 57.950 ;
        RECT 251.740 57.950 254.280 57.970 ;
        RECT 246.235 57.945 248.480 57.950 ;
        RECT 242.545 57.875 244.340 57.945 ;
        POLYGON 244.340 57.945 244.425 57.945 244.340 57.875 ;
        POLYGON 246.215 57.945 246.215 57.875 246.095 57.875 ;
        RECT 246.215 57.930 248.480 57.945 ;
        POLYGON 248.480 57.950 248.585 57.950 248.480 57.930 ;
        POLYGON 251.745 57.950 251.860 57.950 251.860 57.930 ;
        RECT 251.860 57.930 254.280 57.950 ;
        RECT 246.215 57.910 248.395 57.930 ;
        POLYGON 248.395 57.930 248.480 57.930 248.395 57.910 ;
        POLYGON 251.860 57.930 251.920 57.930 251.920 57.920 ;
        RECT 251.920 57.920 254.280 57.930 ;
        POLYGON 251.925 57.920 251.965 57.920 251.965 57.910 ;
        RECT 251.965 57.910 254.280 57.920 ;
        RECT 246.215 57.895 248.320 57.910 ;
        POLYGON 248.320 57.910 248.380 57.910 248.320 57.895 ;
        POLYGON 251.965 57.910 251.990 57.910 251.990 57.905 ;
        RECT 251.990 57.905 254.280 57.910 ;
        POLYGON 252.000 57.905 252.040 57.905 252.040 57.895 ;
        RECT 252.040 57.895 254.280 57.905 ;
        RECT 246.215 57.875 248.185 57.895 ;
        RECT 242.545 57.870 244.260 57.875 ;
        POLYGON 242.440 57.870 242.440 57.805 242.380 57.805 ;
        RECT 242.440 57.810 244.260 57.870 ;
        POLYGON 244.260 57.875 244.340 57.875 244.260 57.810 ;
        POLYGON 246.095 57.875 246.095 57.810 245.980 57.810 ;
        RECT 246.095 57.865 248.185 57.875 ;
        POLYGON 248.185 57.895 248.320 57.895 248.185 57.865 ;
        POLYGON 252.040 57.895 252.060 57.895 252.060 57.890 ;
        RECT 252.060 57.890 254.280 57.895 ;
        POLYGON 252.065 57.890 252.170 57.890 252.170 57.865 ;
        RECT 252.170 57.865 254.280 57.890 ;
        RECT 246.095 57.830 248.050 57.865 ;
        POLYGON 248.050 57.865 248.185 57.865 248.050 57.830 ;
        POLYGON 252.170 57.865 252.255 57.865 252.255 57.845 ;
        RECT 252.255 57.855 254.280 57.865 ;
        POLYGON 254.280 57.985 254.520 57.855 254.280 57.855 ;
        POLYGON 256.355 57.985 256.515 57.985 256.515 57.870 ;
        RECT 256.515 57.955 258.415 57.985 ;
        POLYGON 258.415 58.075 258.545 57.955 258.415 57.955 ;
        POLYGON 260.920 58.075 260.945 58.075 260.945 58.050 ;
        RECT 260.945 58.050 264.040 58.075 ;
        POLYGON 260.945 58.050 261.015 58.050 261.015 57.965 ;
        RECT 261.015 58.010 264.040 58.050 ;
        POLYGON 264.040 58.100 264.105 58.010 264.040 58.010 ;
        POLYGON 268.530 58.100 268.575 58.100 268.575 58.015 ;
        RECT 268.575 58.010 275.775 58.100 ;
        RECT 261.015 57.965 264.105 58.010 ;
        POLYGON 261.015 57.965 261.020 57.965 261.020 57.955 ;
        RECT 261.020 57.955 264.105 57.965 ;
        POLYGON 264.105 58.010 264.140 57.955 264.105 57.955 ;
        POLYGON 268.575 58.010 268.605 58.010 268.605 57.960 ;
        RECT 268.605 57.955 275.775 58.010 ;
        RECT 256.515 57.870 258.545 57.955 ;
        POLYGON 256.515 57.870 256.530 57.870 256.530 57.855 ;
        RECT 256.530 57.855 258.545 57.870 ;
        RECT 252.255 57.845 254.520 57.855 ;
        POLYGON 252.255 57.845 252.305 57.845 252.305 57.830 ;
        RECT 252.305 57.840 254.520 57.845 ;
        POLYGON 254.520 57.855 254.545 57.840 254.520 57.840 ;
        POLYGON 256.530 57.855 256.550 57.855 256.550 57.840 ;
        RECT 256.550 57.840 258.545 57.855 ;
        RECT 252.305 57.830 254.550 57.840 ;
        RECT 246.095 57.810 247.950 57.830 ;
        RECT 242.440 57.805 244.105 57.810 ;
        RECT 238.055 57.795 240.330 57.805 ;
        POLYGON 240.330 57.805 240.335 57.805 240.330 57.795 ;
        POLYGON 242.380 57.805 242.380 57.795 242.370 57.795 ;
        RECT 242.380 57.795 244.105 57.805 ;
        RECT 238.055 57.755 240.230 57.795 ;
        RECT 230.025 57.520 234.430 57.755 ;
        RECT 206.230 57.130 222.255 57.505 ;
        RECT 181.215 57.125 195.525 57.130 ;
        POLYGON 195.525 57.130 195.530 57.125 195.525 57.125 ;
        RECT 181.215 57.075 195.530 57.125 ;
        POLYGON 181.215 57.075 181.330 57.075 181.330 56.745 ;
        RECT 181.330 56.745 195.530 57.075 ;
        RECT 169.860 56.695 174.220 56.745 ;
        RECT 164.690 56.675 166.930 56.695 ;
        POLYGON 164.690 56.675 164.695 56.675 164.695 56.665 ;
        RECT 164.695 56.665 166.930 56.675 ;
        RECT 161.280 56.660 162.825 56.665 ;
        RECT 158.455 56.640 159.775 56.660 ;
        RECT 153.840 56.630 156.745 56.640 ;
        POLYGON 153.750 56.630 153.750 56.625 153.735 56.625 ;
        RECT 153.750 56.625 156.745 56.630 ;
        POLYGON 153.735 56.625 153.735 56.620 153.705 56.620 ;
        RECT 153.735 56.620 156.745 56.625 ;
        POLYGON 156.745 56.640 156.830 56.620 156.745 56.620 ;
        POLYGON 158.455 56.640 158.500 56.640 158.500 56.620 ;
        RECT 158.500 56.620 159.775 56.640 ;
        POLYGON 153.705 56.620 153.705 56.600 153.630 56.600 ;
        RECT 153.705 56.600 156.830 56.620 ;
        RECT 150.545 56.595 151.970 56.600 ;
        POLYGON 151.970 56.600 151.975 56.600 151.970 56.595 ;
        POLYGON 153.630 56.600 153.630 56.595 153.610 56.595 ;
        RECT 153.630 56.595 156.830 56.600 ;
        RECT 150.545 56.580 151.940 56.595 ;
        POLYGON 151.940 56.595 151.970 56.595 151.940 56.580 ;
        POLYGON 153.610 56.595 153.610 56.585 153.575 56.585 ;
        RECT 153.610 56.585 156.830 56.595 ;
        POLYGON 153.575 56.585 153.575 56.580 153.555 56.580 ;
        RECT 153.575 56.580 156.830 56.585 ;
        POLYGON 150.495 56.580 150.495 56.565 150.475 56.565 ;
        RECT 150.495 56.565 151.730 56.580 ;
        RECT 147.995 56.555 149.220 56.565 ;
        POLYGON 147.955 56.555 147.955 56.525 147.925 56.525 ;
        RECT 147.955 56.525 149.220 56.555 ;
        POLYGON 147.925 56.525 147.925 56.515 147.915 56.515 ;
        RECT 147.925 56.515 149.220 56.525 ;
        POLYGON 146.320 56.515 146.345 56.435 146.320 56.435 ;
        RECT 117.310 56.415 146.345 56.435 ;
        POLYGON 147.915 56.515 147.915 56.430 147.840 56.430 ;
        RECT 147.915 56.495 149.220 56.515 ;
        POLYGON 149.220 56.565 149.295 56.565 149.220 56.495 ;
        POLYGON 150.475 56.565 150.475 56.555 150.465 56.555 ;
        RECT 150.475 56.555 151.730 56.565 ;
        POLYGON 150.465 56.555 150.465 56.495 150.390 56.495 ;
        RECT 150.465 56.495 151.730 56.555 ;
        RECT 147.915 56.430 149.140 56.495 ;
        POLYGON 146.345 56.430 146.350 56.415 146.345 56.415 ;
        RECT 117.310 56.390 146.350 56.415 ;
        POLYGON 147.840 56.430 147.840 56.410 147.820 56.410 ;
        RECT 147.840 56.420 149.140 56.430 ;
        POLYGON 149.140 56.495 149.220 56.495 149.140 56.420 ;
        POLYGON 150.390 56.495 150.390 56.420 150.295 56.420 ;
        RECT 150.390 56.470 151.730 56.495 ;
        POLYGON 151.730 56.580 151.940 56.580 151.730 56.470 ;
        POLYGON 153.555 56.580 153.555 56.565 153.495 56.565 ;
        RECT 153.555 56.570 156.830 56.580 ;
        POLYGON 156.830 56.620 157.030 56.570 156.830 56.570 ;
        POLYGON 158.505 56.620 158.550 56.620 158.550 56.590 ;
        RECT 158.550 56.590 159.775 56.620 ;
        POLYGON 158.550 56.590 158.585 56.590 158.585 56.570 ;
        RECT 158.585 56.570 159.775 56.590 ;
        RECT 153.555 56.565 157.030 56.570 ;
        POLYGON 153.480 56.565 153.480 56.515 153.325 56.515 ;
        RECT 153.480 56.535 157.030 56.565 ;
        POLYGON 157.030 56.570 157.155 56.535 157.030 56.535 ;
        POLYGON 158.585 56.570 158.640 56.570 158.640 56.540 ;
        RECT 158.640 56.540 159.775 56.570 ;
        POLYGON 159.775 56.660 159.940 56.540 159.775 56.540 ;
        POLYGON 161.280 56.660 161.305 56.660 161.305 56.640 ;
        RECT 161.305 56.640 162.825 56.660 ;
        POLYGON 161.305 56.640 161.415 56.640 161.415 56.545 ;
        RECT 161.415 56.610 162.825 56.640 ;
        POLYGON 162.825 56.665 162.880 56.610 162.825 56.610 ;
        POLYGON 164.695 56.665 164.705 56.665 164.705 56.655 ;
        RECT 164.705 56.655 166.930 56.665 ;
        POLYGON 164.705 56.655 164.735 56.655 164.735 56.615 ;
        RECT 164.735 56.610 166.930 56.655 ;
        RECT 161.415 56.550 162.880 56.610 ;
        POLYGON 162.880 56.610 162.935 56.550 162.880 56.550 ;
        POLYGON 164.735 56.610 164.785 56.610 164.785 56.550 ;
        RECT 164.785 56.550 166.930 56.610 ;
        RECT 161.415 56.545 162.935 56.550 ;
        POLYGON 161.415 56.545 161.420 56.545 161.420 56.540 ;
        RECT 161.420 56.540 162.935 56.545 ;
        POLYGON 158.640 56.540 158.645 56.540 158.645 56.535 ;
        RECT 158.645 56.535 159.940 56.540 ;
        RECT 153.480 56.515 157.160 56.535 ;
        POLYGON 153.320 56.515 153.320 56.510 153.305 56.510 ;
        RECT 153.320 56.510 157.160 56.515 ;
        POLYGON 157.160 56.535 157.250 56.510 157.160 56.510 ;
        POLYGON 158.645 56.535 158.695 56.535 158.695 56.510 ;
        RECT 158.695 56.510 159.940 56.535 ;
        POLYGON 153.305 56.510 153.305 56.485 153.225 56.485 ;
        RECT 153.305 56.505 157.250 56.510 ;
        POLYGON 157.250 56.510 157.265 56.505 157.250 56.505 ;
        POLYGON 158.695 56.510 158.705 56.510 158.705 56.505 ;
        RECT 158.705 56.505 159.940 56.510 ;
        RECT 153.305 56.490 157.265 56.505 ;
        POLYGON 157.265 56.505 157.315 56.490 157.265 56.490 ;
        POLYGON 158.705 56.505 158.735 56.505 158.735 56.490 ;
        RECT 158.735 56.490 159.940 56.505 ;
        RECT 153.305 56.485 157.315 56.490 ;
        POLYGON 153.225 56.485 153.225 56.470 153.175 56.470 ;
        RECT 153.225 56.470 157.315 56.485 ;
        RECT 150.390 56.440 151.675 56.470 ;
        POLYGON 151.675 56.470 151.725 56.470 151.675 56.440 ;
        POLYGON 153.175 56.470 153.175 56.445 153.090 56.445 ;
        RECT 153.175 56.455 157.315 56.470 ;
        POLYGON 157.315 56.490 157.425 56.455 157.315 56.455 ;
        POLYGON 158.735 56.490 158.745 56.490 158.745 56.485 ;
        RECT 158.745 56.485 159.940 56.490 ;
        POLYGON 158.745 56.485 158.760 56.485 158.760 56.475 ;
        RECT 158.760 56.475 159.940 56.485 ;
        POLYGON 158.765 56.475 158.795 56.475 158.795 56.455 ;
        RECT 158.795 56.455 159.940 56.475 ;
        RECT 153.175 56.445 157.425 56.455 ;
        POLYGON 153.090 56.445 153.090 56.440 153.075 56.440 ;
        RECT 153.090 56.440 157.425 56.445 ;
        RECT 150.390 56.420 151.585 56.440 ;
        RECT 147.840 56.410 149.090 56.420 ;
        RECT 51.940 55.610 111.200 56.390 ;
        POLYGON 111.200 56.390 111.225 55.610 111.200 55.610 ;
        RECT 117.290 56.380 146.350 56.390 ;
        POLYGON 146.350 56.410 146.360 56.380 146.350 56.380 ;
        POLYGON 117.290 56.365 117.290 55.610 117.275 55.610 ;
        RECT 117.290 56.325 146.360 56.380 ;
        POLYGON 147.820 56.410 147.820 56.375 147.790 56.375 ;
        RECT 147.820 56.375 149.090 56.410 ;
        POLYGON 149.090 56.420 149.140 56.420 149.090 56.375 ;
        POLYGON 150.295 56.420 150.295 56.375 150.235 56.375 ;
        RECT 150.295 56.390 151.585 56.420 ;
        POLYGON 151.585 56.440 151.675 56.440 151.585 56.390 ;
        POLYGON 153.075 56.440 153.075 56.430 153.040 56.430 ;
        RECT 153.075 56.430 157.425 56.440 ;
        POLYGON 153.040 56.430 153.040 56.405 152.975 56.405 ;
        RECT 153.040 56.405 157.425 56.430 ;
        POLYGON 152.970 56.405 152.970 56.390 152.935 56.390 ;
        RECT 152.970 56.400 157.425 56.405 ;
        POLYGON 157.425 56.455 157.590 56.400 157.425 56.400 ;
        POLYGON 158.795 56.455 158.885 56.455 158.885 56.400 ;
        RECT 158.885 56.400 159.940 56.455 ;
        POLYGON 159.940 56.540 160.130 56.400 159.940 56.400 ;
        POLYGON 161.420 56.540 161.555 56.540 161.555 56.415 ;
        RECT 161.555 56.410 162.935 56.540 ;
        POLYGON 161.555 56.410 161.565 56.410 161.565 56.400 ;
        RECT 161.565 56.400 162.935 56.410 ;
        RECT 152.970 56.390 157.590 56.400 ;
        RECT 150.295 56.375 151.490 56.390 ;
        POLYGON 146.360 56.375 146.375 56.325 146.360 56.325 ;
        RECT 117.290 56.270 146.375 56.325 ;
        POLYGON 147.790 56.375 147.790 56.320 147.745 56.320 ;
        RECT 147.790 56.320 148.935 56.375 ;
        POLYGON 146.375 56.315 146.390 56.270 146.375 56.270 ;
        RECT 117.290 56.235 146.390 56.270 ;
        POLYGON 147.745 56.315 147.745 56.265 147.700 56.265 ;
        RECT 147.745 56.265 148.935 56.320 ;
        POLYGON 146.390 56.265 146.400 56.235 146.390 56.235 ;
        POLYGON 147.700 56.265 147.700 56.240 147.680 56.240 ;
        RECT 147.700 56.240 148.935 56.265 ;
        RECT 117.290 56.145 146.400 56.235 ;
        POLYGON 146.400 56.235 146.425 56.145 146.400 56.145 ;
        POLYGON 147.680 56.235 147.680 56.145 147.605 56.145 ;
        RECT 147.680 56.220 148.935 56.240 ;
        POLYGON 148.935 56.375 149.090 56.375 148.935 56.220 ;
        POLYGON 150.230 56.375 150.230 56.305 150.150 56.305 ;
        RECT 150.230 56.335 151.490 56.375 ;
        POLYGON 151.490 56.390 151.585 56.390 151.490 56.335 ;
        POLYGON 152.935 56.390 152.935 56.375 152.900 56.375 ;
        RECT 152.935 56.375 157.590 56.390 ;
        POLYGON 152.900 56.375 152.900 56.335 152.785 56.335 ;
        RECT 152.900 56.360 157.590 56.375 ;
        POLYGON 157.590 56.400 157.690 56.360 157.590 56.360 ;
        POLYGON 158.885 56.400 158.945 56.400 158.945 56.360 ;
        RECT 158.945 56.370 160.130 56.400 ;
        POLYGON 160.130 56.400 160.165 56.370 160.130 56.370 ;
        POLYGON 161.565 56.400 161.600 56.400 161.600 56.370 ;
        RECT 161.600 56.370 162.935 56.400 ;
        RECT 158.945 56.360 160.165 56.370 ;
        RECT 152.900 56.355 157.690 56.360 ;
        POLYGON 157.690 56.360 157.700 56.355 157.690 56.355 ;
        POLYGON 158.945 56.360 158.955 56.360 158.955 56.355 ;
        RECT 158.955 56.355 160.165 56.360 ;
        POLYGON 160.165 56.370 160.185 56.355 160.165 56.355 ;
        POLYGON 161.600 56.370 161.620 56.370 161.620 56.355 ;
        RECT 161.620 56.355 162.935 56.370 ;
        RECT 152.900 56.335 157.700 56.355 ;
        RECT 150.230 56.305 151.285 56.335 ;
        POLYGON 150.150 56.305 150.150 56.295 150.135 56.295 ;
        RECT 150.150 56.295 151.285 56.305 ;
        POLYGON 150.135 56.295 150.135 56.220 150.055 56.220 ;
        RECT 150.135 56.220 151.285 56.295 ;
        RECT 147.680 56.210 148.930 56.220 ;
        POLYGON 148.930 56.220 148.935 56.220 148.930 56.210 ;
        POLYGON 150.055 56.220 150.055 56.210 150.045 56.210 ;
        RECT 150.055 56.210 151.285 56.220 ;
        POLYGON 151.285 56.335 151.485 56.335 151.285 56.210 ;
        POLYGON 152.785 56.335 152.785 56.330 152.770 56.330 ;
        RECT 152.785 56.330 157.700 56.335 ;
        POLYGON 152.770 56.330 152.770 56.310 152.720 56.310 ;
        RECT 152.770 56.310 157.700 56.330 ;
        POLYGON 152.720 56.310 152.720 56.300 152.690 56.300 ;
        RECT 152.720 56.300 157.700 56.310 ;
        POLYGON 152.690 56.300 152.690 56.220 152.505 56.220 ;
        RECT 152.690 56.295 157.700 56.300 ;
        POLYGON 157.700 56.355 157.865 56.295 157.700 56.295 ;
        POLYGON 158.955 56.355 158.965 56.355 158.965 56.350 ;
        RECT 158.965 56.350 160.185 56.355 ;
        POLYGON 158.965 56.350 158.990 56.350 158.990 56.340 ;
        RECT 158.990 56.345 160.185 56.350 ;
        POLYGON 160.185 56.355 160.195 56.345 160.185 56.345 ;
        POLYGON 161.620 56.355 161.630 56.355 161.630 56.345 ;
        RECT 161.630 56.345 162.935 56.355 ;
        RECT 158.990 56.340 160.195 56.345 ;
        POLYGON 158.990 56.340 159.015 56.340 159.015 56.320 ;
        RECT 159.015 56.320 160.195 56.340 ;
        POLYGON 159.015 56.320 159.050 56.320 159.050 56.295 ;
        RECT 159.050 56.295 160.195 56.320 ;
        RECT 152.690 56.260 157.865 56.295 ;
        RECT 152.690 56.255 155.045 56.260 ;
        POLYGON 155.045 56.260 155.170 56.260 155.045 56.255 ;
        POLYGON 155.250 56.260 155.265 56.260 155.265 56.255 ;
        RECT 155.265 56.255 157.865 56.260 ;
        POLYGON 157.865 56.295 157.960 56.255 157.865 56.255 ;
        POLYGON 159.050 56.295 159.115 56.295 159.115 56.255 ;
        RECT 159.115 56.255 160.195 56.295 ;
        RECT 152.690 56.250 154.835 56.255 ;
        POLYGON 154.835 56.255 154.910 56.255 154.835 56.250 ;
        POLYGON 155.460 56.255 155.505 56.255 155.505 56.250 ;
        RECT 155.505 56.250 157.960 56.255 ;
        RECT 152.690 56.240 154.645 56.250 ;
        POLYGON 154.645 56.250 154.785 56.250 154.645 56.240 ;
        POLYGON 155.555 56.250 155.625 56.250 155.625 56.245 ;
        RECT 155.625 56.245 157.960 56.250 ;
        POLYGON 155.665 56.245 155.755 56.245 155.755 56.240 ;
        RECT 155.755 56.240 157.960 56.245 ;
        RECT 152.690 56.235 154.570 56.240 ;
        POLYGON 154.570 56.240 154.640 56.240 154.570 56.235 ;
        POLYGON 155.755 56.240 155.850 56.240 155.850 56.235 ;
        RECT 155.850 56.235 157.960 56.240 ;
        POLYGON 157.960 56.255 158.005 56.235 157.960 56.235 ;
        POLYGON 159.115 56.255 159.125 56.255 159.125 56.250 ;
        RECT 159.125 56.250 160.195 56.255 ;
        POLYGON 159.125 56.250 159.145 56.250 159.145 56.235 ;
        RECT 159.145 56.235 160.195 56.250 ;
        RECT 152.690 56.230 154.535 56.235 ;
        POLYGON 154.535 56.235 154.565 56.235 154.535 56.230 ;
        POLYGON 155.850 56.235 155.920 56.235 155.920 56.230 ;
        RECT 155.920 56.230 158.005 56.235 ;
        RECT 152.690 56.220 154.430 56.230 ;
        POLYGON 154.430 56.230 154.505 56.230 154.430 56.220 ;
        POLYGON 155.920 56.230 155.965 56.230 155.965 56.225 ;
        RECT 155.965 56.225 158.005 56.230 ;
        POLYGON 155.970 56.225 156.020 56.225 156.020 56.220 ;
        RECT 156.020 56.220 158.005 56.225 ;
        POLYGON 152.505 56.220 152.505 56.210 152.485 56.210 ;
        RECT 152.505 56.215 154.350 56.220 ;
        POLYGON 154.350 56.220 154.430 56.220 154.350 56.215 ;
        POLYGON 156.020 56.220 156.070 56.220 156.070 56.215 ;
        RECT 156.070 56.215 158.005 56.220 ;
        RECT 152.505 56.210 154.220 56.215 ;
        RECT 147.680 56.165 148.890 56.210 ;
        POLYGON 148.890 56.210 148.930 56.210 148.890 56.165 ;
        POLYGON 150.045 56.210 150.045 56.175 150.005 56.175 ;
        RECT 150.045 56.195 151.265 56.210 ;
        POLYGON 151.265 56.210 151.285 56.210 151.265 56.195 ;
        POLYGON 152.485 56.210 152.485 56.205 152.470 56.205 ;
        RECT 152.485 56.205 154.220 56.210 ;
        POLYGON 152.470 56.205 152.470 56.195 152.445 56.195 ;
        RECT 152.470 56.200 154.220 56.205 ;
        POLYGON 154.220 56.215 154.345 56.215 154.220 56.200 ;
        POLYGON 156.080 56.215 156.125 56.215 156.125 56.210 ;
        RECT 156.125 56.210 158.005 56.215 ;
        POLYGON 156.130 56.210 156.135 56.210 156.135 56.205 ;
        RECT 156.135 56.205 158.005 56.210 ;
        POLYGON 156.155 56.205 156.210 56.205 156.210 56.200 ;
        RECT 156.210 56.200 158.005 56.205 ;
        RECT 152.470 56.195 154.180 56.200 ;
        POLYGON 154.180 56.200 154.215 56.200 154.180 56.195 ;
        POLYGON 156.210 56.200 156.270 56.200 156.270 56.195 ;
        RECT 156.270 56.195 158.005 56.200 ;
        RECT 150.045 56.185 151.245 56.195 ;
        POLYGON 151.245 56.195 151.265 56.195 151.245 56.185 ;
        POLYGON 152.445 56.195 152.445 56.185 152.425 56.185 ;
        RECT 152.445 56.190 154.140 56.195 ;
        POLYGON 154.140 56.195 154.180 56.195 154.140 56.190 ;
        POLYGON 156.270 56.195 156.290 56.195 156.290 56.190 ;
        RECT 156.290 56.190 158.005 56.195 ;
        RECT 152.445 56.185 154.130 56.190 ;
        POLYGON 154.130 56.190 154.140 56.190 154.130 56.185 ;
        POLYGON 156.290 56.190 156.315 56.190 156.315 56.185 ;
        RECT 156.315 56.185 158.005 56.190 ;
        RECT 150.045 56.175 151.040 56.185 ;
        POLYGON 150.005 56.175 150.005 56.165 149.995 56.165 ;
        RECT 150.005 56.165 151.040 56.175 ;
        RECT 147.680 56.145 148.760 56.165 ;
        RECT 117.290 56.110 146.425 56.145 ;
        POLYGON 146.425 56.145 146.435 56.110 146.425 56.110 ;
        RECT 117.290 56.090 146.435 56.110 ;
        POLYGON 147.605 56.145 147.605 56.100 147.565 56.100 ;
        RECT 147.605 56.100 148.760 56.145 ;
        POLYGON 146.435 56.100 146.440 56.090 146.435 56.090 ;
        RECT 117.290 55.985 146.440 56.090 ;
        POLYGON 147.565 56.100 147.565 56.085 147.555 56.085 ;
        RECT 147.565 56.085 148.760 56.100 ;
        POLYGON 147.555 56.085 147.555 56.080 147.550 56.080 ;
        RECT 147.555 56.080 148.760 56.085 ;
        POLYGON 146.440 56.080 146.470 55.985 146.440 55.985 ;
        RECT 117.290 55.875 146.470 55.985 ;
        POLYGON 147.550 56.080 147.550 55.970 147.465 55.970 ;
        RECT 147.550 56.030 148.760 56.080 ;
        POLYGON 148.760 56.165 148.890 56.165 148.760 56.030 ;
        POLYGON 149.995 56.165 149.995 56.045 149.850 56.045 ;
        RECT 149.995 56.050 151.040 56.165 ;
        POLYGON 151.040 56.185 151.245 56.185 151.040 56.050 ;
        POLYGON 152.425 56.185 152.425 56.135 152.310 56.135 ;
        RECT 152.425 56.165 154.010 56.185 ;
        POLYGON 154.010 56.185 154.130 56.185 154.010 56.165 ;
        POLYGON 156.315 56.185 156.435 56.185 156.435 56.165 ;
        RECT 156.435 56.180 158.005 56.185 ;
        POLYGON 158.005 56.235 158.130 56.180 158.005 56.180 ;
        POLYGON 159.145 56.235 159.230 56.235 159.230 56.180 ;
        RECT 159.230 56.180 160.195 56.235 ;
        RECT 156.435 56.165 158.130 56.180 ;
        RECT 152.425 56.150 153.915 56.165 ;
        POLYGON 153.915 56.165 154.005 56.165 153.915 56.150 ;
        POLYGON 156.450 56.165 156.505 56.165 156.505 56.155 ;
        RECT 156.505 56.155 158.130 56.165 ;
        POLYGON 156.510 56.155 156.545 56.155 156.545 56.150 ;
        RECT 156.545 56.150 158.130 56.155 ;
        RECT 152.425 56.145 153.865 56.150 ;
        POLYGON 153.865 56.150 153.915 56.150 153.865 56.145 ;
        POLYGON 156.545 56.150 156.585 56.150 156.585 56.145 ;
        RECT 156.585 56.145 158.130 56.150 ;
        RECT 152.425 56.135 153.795 56.145 ;
        POLYGON 152.310 56.135 152.310 56.095 152.235 56.095 ;
        RECT 152.310 56.130 153.795 56.135 ;
        POLYGON 153.795 56.145 153.865 56.145 153.795 56.130 ;
        POLYGON 156.590 56.145 156.605 56.145 156.605 56.140 ;
        RECT 156.605 56.140 158.130 56.145 ;
        POLYGON 156.605 56.140 156.655 56.140 156.655 56.130 ;
        RECT 156.655 56.130 158.130 56.140 ;
        RECT 152.310 56.120 153.740 56.130 ;
        POLYGON 153.740 56.130 153.790 56.130 153.740 56.120 ;
        POLYGON 156.655 56.130 156.710 56.130 156.710 56.120 ;
        RECT 156.710 56.125 158.130 56.130 ;
        POLYGON 158.130 56.180 158.235 56.125 158.130 56.125 ;
        POLYGON 159.230 56.180 159.260 56.180 159.260 56.160 ;
        RECT 159.260 56.160 160.195 56.180 ;
        POLYGON 159.260 56.160 159.305 56.160 159.305 56.125 ;
        RECT 159.305 56.135 160.195 56.160 ;
        POLYGON 160.195 56.345 160.445 56.135 160.195 56.135 ;
        POLYGON 161.630 56.345 161.645 56.345 161.645 56.330 ;
        RECT 161.645 56.340 162.935 56.345 ;
        POLYGON 162.935 56.550 163.120 56.340 162.935 56.340 ;
        POLYGON 164.785 56.550 164.795 56.550 164.795 56.535 ;
        RECT 164.795 56.545 166.930 56.550 ;
        POLYGON 166.930 56.695 167.020 56.545 166.930 56.545 ;
        POLYGON 169.860 56.695 169.885 56.695 169.885 56.655 ;
        RECT 169.885 56.655 174.220 56.695 ;
        POLYGON 169.885 56.655 169.935 56.655 169.935 56.550 ;
        RECT 169.935 56.545 174.220 56.655 ;
        RECT 164.795 56.535 167.020 56.545 ;
        POLYGON 164.795 56.535 164.855 56.535 164.855 56.460 ;
        RECT 164.855 56.460 167.020 56.535 ;
        POLYGON 164.855 56.460 164.870 56.460 164.870 56.435 ;
        RECT 164.870 56.435 167.020 56.460 ;
        POLYGON 164.870 56.435 164.895 56.435 164.895 56.395 ;
        RECT 164.895 56.400 167.020 56.435 ;
        POLYGON 167.020 56.545 167.110 56.400 167.020 56.400 ;
        POLYGON 169.935 56.545 170.005 56.545 170.005 56.400 ;
        RECT 170.005 56.415 174.220 56.545 ;
        POLYGON 174.220 56.745 174.375 56.415 174.220 56.415 ;
        POLYGON 181.330 56.745 181.445 56.745 181.445 56.420 ;
        RECT 181.445 56.415 195.530 56.745 ;
        RECT 170.005 56.400 174.375 56.415 ;
        RECT 164.895 56.395 167.110 56.400 ;
        POLYGON 164.895 56.395 164.935 56.395 164.935 56.340 ;
        RECT 164.935 56.340 167.110 56.395 ;
        RECT 161.645 56.335 163.120 56.340 ;
        POLYGON 163.120 56.340 163.125 56.335 163.120 56.335 ;
        POLYGON 164.935 56.340 164.940 56.340 164.940 56.335 ;
        RECT 164.940 56.335 167.110 56.340 ;
        RECT 161.645 56.330 163.125 56.335 ;
        POLYGON 161.645 56.330 161.835 56.330 161.835 56.135 ;
        RECT 161.835 56.190 163.125 56.330 ;
        POLYGON 163.125 56.335 163.245 56.190 163.125 56.190 ;
        POLYGON 164.940 56.335 164.955 56.335 164.955 56.315 ;
        RECT 164.955 56.315 167.110 56.335 ;
        POLYGON 164.955 56.315 164.980 56.315 164.980 56.275 ;
        RECT 164.980 56.280 167.110 56.315 ;
        POLYGON 167.110 56.400 167.180 56.280 167.110 56.280 ;
        POLYGON 170.005 56.400 170.060 56.400 170.060 56.285 ;
        RECT 170.060 56.295 174.375 56.400 ;
        POLYGON 174.375 56.415 174.425 56.295 174.375 56.295 ;
        POLYGON 181.445 56.415 181.490 56.415 181.490 56.295 ;
        RECT 181.490 56.295 195.530 56.415 ;
        RECT 170.060 56.280 174.425 56.295 ;
        RECT 164.980 56.275 167.180 56.280 ;
        POLYGON 164.980 56.275 165.035 56.275 165.035 56.190 ;
        RECT 165.035 56.190 167.180 56.275 ;
        RECT 161.835 56.135 163.245 56.190 ;
        POLYGON 163.245 56.190 163.285 56.135 163.245 56.135 ;
        POLYGON 165.035 56.190 165.055 56.190 165.055 56.165 ;
        RECT 165.055 56.165 167.180 56.190 ;
        POLYGON 165.055 56.165 165.080 56.165 165.080 56.135 ;
        RECT 165.080 56.135 167.180 56.165 ;
        RECT 159.305 56.125 160.445 56.135 ;
        RECT 156.710 56.120 158.235 56.125 ;
        POLYGON 158.235 56.125 158.250 56.120 158.235 56.120 ;
        POLYGON 159.305 56.125 159.310 56.125 159.310 56.120 ;
        RECT 159.310 56.120 160.445 56.125 ;
        RECT 152.310 56.110 153.705 56.120 ;
        POLYGON 153.705 56.120 153.740 56.120 153.705 56.110 ;
        POLYGON 156.715 56.120 156.720 56.120 156.720 56.115 ;
        RECT 156.720 56.115 158.255 56.120 ;
        POLYGON 156.720 56.115 156.745 56.115 156.745 56.110 ;
        RECT 156.745 56.110 158.255 56.115 ;
        RECT 152.310 56.095 153.530 56.110 ;
        POLYGON 152.235 56.095 152.235 56.090 152.220 56.090 ;
        RECT 152.235 56.090 153.530 56.095 ;
        POLYGON 152.220 56.085 152.220 56.050 152.150 56.050 ;
        RECT 152.220 56.075 153.530 56.090 ;
        POLYGON 153.530 56.110 153.705 56.110 153.530 56.075 ;
        POLYGON 156.745 56.110 156.840 56.110 156.840 56.090 ;
        RECT 156.840 56.090 158.255 56.110 ;
        POLYGON 156.845 56.090 156.905 56.090 156.905 56.075 ;
        RECT 156.905 56.075 158.255 56.090 ;
        RECT 152.220 56.065 153.495 56.075 ;
        POLYGON 153.495 56.075 153.530 56.075 153.495 56.065 ;
        POLYGON 156.905 56.075 156.925 56.075 156.925 56.070 ;
        RECT 156.925 56.070 158.255 56.075 ;
        POLYGON 156.935 56.070 156.950 56.070 156.950 56.065 ;
        RECT 156.950 56.065 158.255 56.070 ;
        RECT 152.220 56.050 153.365 56.065 ;
        RECT 149.995 56.045 151.010 56.050 ;
        POLYGON 149.850 56.045 149.850 56.030 149.835 56.030 ;
        RECT 149.850 56.030 151.010 56.045 ;
        RECT 147.550 56.010 148.740 56.030 ;
        POLYGON 148.740 56.030 148.760 56.030 148.740 56.010 ;
        POLYGON 149.835 56.030 149.835 56.010 149.815 56.010 ;
        RECT 149.835 56.025 151.010 56.030 ;
        POLYGON 151.010 56.050 151.040 56.050 151.010 56.025 ;
        POLYGON 152.150 56.050 152.150 56.025 152.095 56.025 ;
        RECT 152.150 56.030 153.365 56.050 ;
        POLYGON 153.365 56.065 153.495 56.065 153.365 56.030 ;
        POLYGON 156.950 56.065 156.970 56.065 156.970 56.060 ;
        RECT 156.970 56.060 158.255 56.065 ;
        POLYGON 156.975 56.060 157.030 56.060 157.030 56.045 ;
        RECT 157.030 56.050 158.255 56.060 ;
        POLYGON 158.255 56.120 158.385 56.050 158.255 56.050 ;
        POLYGON 159.310 56.120 159.355 56.120 159.355 56.090 ;
        RECT 159.355 56.095 160.445 56.120 ;
        POLYGON 160.445 56.135 160.495 56.095 160.445 56.095 ;
        POLYGON 161.835 56.135 161.850 56.135 161.850 56.120 ;
        RECT 161.850 56.120 163.285 56.135 ;
        POLYGON 161.850 56.120 161.865 56.120 161.865 56.100 ;
        RECT 161.865 56.100 163.285 56.120 ;
        POLYGON 161.865 56.100 161.870 56.100 161.870 56.095 ;
        RECT 161.870 56.095 163.285 56.100 ;
        RECT 159.355 56.090 160.495 56.095 ;
        POLYGON 159.355 56.090 159.375 56.090 159.375 56.080 ;
        RECT 159.375 56.080 160.495 56.090 ;
        POLYGON 159.375 56.080 159.415 56.080 159.415 56.050 ;
        RECT 159.415 56.055 160.495 56.080 ;
        POLYGON 160.495 56.095 160.540 56.055 160.495 56.055 ;
        POLYGON 161.870 56.095 161.890 56.095 161.890 56.080 ;
        RECT 161.890 56.080 163.285 56.095 ;
        POLYGON 161.890 56.080 161.905 56.080 161.905 56.060 ;
        RECT 161.905 56.055 163.285 56.080 ;
        RECT 159.415 56.050 160.540 56.055 ;
        RECT 157.030 56.045 158.385 56.050 ;
        POLYGON 157.030 56.045 157.075 56.045 157.075 56.030 ;
        RECT 157.075 56.030 158.385 56.045 ;
        RECT 152.150 56.025 153.325 56.030 ;
        RECT 149.835 56.010 150.920 56.025 ;
        RECT 147.550 55.970 148.660 56.010 ;
        POLYGON 146.470 55.970 146.500 55.875 146.470 55.875 ;
        POLYGON 147.465 55.970 147.465 55.880 147.395 55.880 ;
        RECT 147.465 55.915 148.660 55.970 ;
        POLYGON 148.660 56.010 148.740 56.010 148.660 55.915 ;
        POLYGON 149.815 56.010 149.815 55.975 149.780 55.975 ;
        RECT 149.815 55.975 150.920 56.010 ;
        POLYGON 149.780 55.970 149.780 55.915 149.720 55.915 ;
        RECT 149.780 55.965 150.920 55.975 ;
        POLYGON 150.920 56.025 151.010 56.025 150.920 55.965 ;
        POLYGON 152.095 56.025 152.095 56.015 152.075 56.015 ;
        RECT 152.095 56.020 153.325 56.025 ;
        POLYGON 153.325 56.030 153.365 56.030 153.325 56.020 ;
        POLYGON 157.075 56.030 157.110 56.030 157.110 56.020 ;
        RECT 157.110 56.020 158.385 56.030 ;
        RECT 152.095 56.015 153.255 56.020 ;
        POLYGON 152.075 56.015 152.075 55.965 151.985 55.965 ;
        RECT 152.075 56.005 153.255 56.015 ;
        POLYGON 153.255 56.020 153.325 56.020 153.255 56.005 ;
        POLYGON 157.110 56.020 157.150 56.020 157.150 56.010 ;
        RECT 157.150 56.010 158.385 56.020 ;
        POLYGON 157.150 56.010 157.165 56.010 157.165 56.005 ;
        RECT 157.165 56.005 158.385 56.010 ;
        RECT 152.075 55.970 153.150 56.005 ;
        POLYGON 153.150 56.005 153.255 56.005 153.150 55.970 ;
        POLYGON 157.165 56.005 157.235 56.005 157.235 55.985 ;
        RECT 157.235 55.990 158.385 56.005 ;
        POLYGON 158.385 56.050 158.500 55.990 158.385 55.990 ;
        POLYGON 159.415 56.050 159.465 56.050 159.465 56.015 ;
        RECT 159.465 56.015 160.540 56.050 ;
        POLYGON 159.465 56.015 159.495 56.015 159.495 55.995 ;
        RECT 159.495 55.995 160.540 56.015 ;
        POLYGON 159.495 55.995 159.500 55.995 159.500 55.990 ;
        RECT 159.500 55.990 160.540 55.995 ;
        POLYGON 160.540 56.055 160.615 55.990 160.540 55.990 ;
        POLYGON 161.905 56.055 161.965 56.055 161.965 55.990 ;
        RECT 161.965 56.000 163.285 56.055 ;
        POLYGON 163.285 56.135 163.395 56.000 163.285 56.000 ;
        POLYGON 165.080 56.135 165.100 56.135 165.100 56.100 ;
        RECT 165.100 56.100 167.180 56.135 ;
        POLYGON 165.100 56.100 165.125 56.100 165.125 56.060 ;
        RECT 165.125 56.060 167.180 56.100 ;
        POLYGON 165.125 56.060 165.140 56.060 165.140 56.035 ;
        RECT 165.140 56.035 167.180 56.060 ;
        POLYGON 165.140 56.035 165.160 56.035 165.160 56.005 ;
        RECT 165.160 56.000 167.180 56.035 ;
        RECT 161.965 55.990 163.395 56.000 ;
        RECT 157.235 55.985 158.505 55.990 ;
        POLYGON 157.235 55.985 157.280 55.985 157.280 55.970 ;
        RECT 157.280 55.970 158.505 55.985 ;
        RECT 152.075 55.965 153.125 55.970 ;
        POLYGON 153.125 55.970 153.145 55.970 153.125 55.965 ;
        POLYGON 157.280 55.970 157.295 55.970 157.295 55.965 ;
        RECT 157.295 55.965 158.505 55.970 ;
        RECT 149.780 55.955 150.910 55.965 ;
        POLYGON 150.910 55.965 150.920 55.965 150.910 55.955 ;
        POLYGON 151.985 55.965 151.985 55.960 151.975 55.960 ;
        RECT 151.985 55.960 153.090 55.965 ;
        POLYGON 151.970 55.960 151.970 55.955 151.960 55.955 ;
        RECT 151.970 55.955 153.090 55.960 ;
        RECT 149.780 55.915 150.830 55.955 ;
        RECT 147.465 55.880 148.550 55.915 ;
        RECT 117.290 55.855 146.500 55.875 ;
        POLYGON 146.500 55.875 146.505 55.855 146.500 55.855 ;
        RECT 117.290 55.785 146.505 55.855 ;
        POLYGON 147.395 55.875 147.395 55.845 147.370 55.845 ;
        RECT 147.395 55.845 148.550 55.880 ;
        POLYGON 146.505 55.845 146.525 55.785 146.505 55.785 ;
        RECT 117.290 55.730 146.525 55.785 ;
        POLYGON 147.370 55.845 147.370 55.780 147.320 55.780 ;
        RECT 147.370 55.795 148.550 55.845 ;
        POLYGON 148.550 55.915 148.660 55.915 148.550 55.795 ;
        POLYGON 149.720 55.915 149.720 55.795 149.600 55.795 ;
        RECT 149.720 55.900 150.830 55.915 ;
        POLYGON 150.830 55.955 150.910 55.955 150.830 55.900 ;
        POLYGON 151.960 55.955 151.960 55.945 151.940 55.945 ;
        RECT 151.960 55.950 153.090 55.955 ;
        POLYGON 153.090 55.965 153.125 55.965 153.090 55.950 ;
        POLYGON 157.295 55.965 157.315 55.965 157.315 55.960 ;
        RECT 157.315 55.960 158.505 55.965 ;
        POLYGON 157.315 55.960 157.345 55.960 157.345 55.950 ;
        RECT 157.345 55.950 158.505 55.960 ;
        RECT 151.960 55.945 152.960 55.950 ;
        POLYGON 151.940 55.945 151.940 55.900 151.865 55.900 ;
        RECT 151.940 55.915 152.960 55.945 ;
        POLYGON 152.960 55.950 153.090 55.950 152.960 55.915 ;
        POLYGON 157.345 55.950 157.360 55.950 157.360 55.945 ;
        RECT 157.360 55.945 158.505 55.950 ;
        POLYGON 157.365 55.945 157.385 55.945 157.385 55.940 ;
        RECT 157.385 55.935 158.505 55.945 ;
        POLYGON 157.385 55.935 157.445 55.935 157.445 55.915 ;
        RECT 157.445 55.915 158.505 55.935 ;
        POLYGON 158.505 55.990 158.640 55.915 158.505 55.915 ;
        POLYGON 159.500 55.990 159.600 55.990 159.600 55.915 ;
        RECT 159.600 55.915 160.615 55.990 ;
        POLYGON 160.615 55.990 160.695 55.915 160.615 55.915 ;
        POLYGON 161.965 55.990 162.030 55.990 162.030 55.920 ;
        RECT 162.030 55.945 163.395 55.990 ;
        POLYGON 163.395 56.000 163.440 55.945 163.395 55.945 ;
        POLYGON 165.160 56.000 165.190 56.000 165.190 55.960 ;
        RECT 165.190 55.960 167.180 56.000 ;
        POLYGON 165.190 55.960 165.195 55.960 165.195 55.950 ;
        RECT 165.195 55.945 167.180 55.960 ;
        RECT 162.030 55.915 163.440 55.945 ;
        RECT 151.940 55.900 152.930 55.915 ;
        POLYGON 152.930 55.915 152.960 55.915 152.930 55.900 ;
        POLYGON 157.445 55.915 157.490 55.915 157.490 55.900 ;
        RECT 157.490 55.900 158.640 55.915 ;
        RECT 149.720 55.855 150.770 55.900 ;
        POLYGON 150.770 55.900 150.830 55.900 150.770 55.855 ;
        POLYGON 151.865 55.900 151.865 55.855 151.790 55.855 ;
        RECT 151.865 55.855 152.730 55.900 ;
        RECT 149.720 55.795 150.625 55.855 ;
        RECT 147.370 55.780 148.495 55.795 ;
        POLYGON 147.320 55.780 147.320 55.775 147.315 55.775 ;
        RECT 147.320 55.775 148.495 55.780 ;
        POLYGON 146.525 55.770 146.540 55.730 146.525 55.730 ;
        POLYGON 147.315 55.770 147.315 55.730 147.285 55.730 ;
        RECT 147.315 55.730 148.495 55.775 ;
        RECT 117.290 55.675 146.540 55.730 ;
        POLYGON 146.540 55.730 146.555 55.675 146.540 55.675 ;
        RECT 117.290 55.660 146.555 55.675 ;
        POLYGON 147.285 55.730 147.285 55.665 147.240 55.665 ;
        RECT 147.285 55.725 148.495 55.730 ;
        POLYGON 148.495 55.795 148.550 55.795 148.495 55.725 ;
        POLYGON 149.600 55.795 149.600 55.755 149.560 55.755 ;
        RECT 149.600 55.755 150.625 55.795 ;
        POLYGON 149.560 55.755 149.560 55.725 149.525 55.725 ;
        RECT 149.560 55.740 150.625 55.755 ;
        POLYGON 150.625 55.855 150.770 55.855 150.625 55.740 ;
        POLYGON 151.790 55.855 151.790 55.820 151.730 55.820 ;
        RECT 151.790 55.830 152.730 55.855 ;
        POLYGON 152.730 55.900 152.925 55.900 152.730 55.830 ;
        POLYGON 157.490 55.900 157.535 55.900 157.535 55.885 ;
        RECT 157.535 55.885 158.640 55.900 ;
        POLYGON 157.535 55.885 157.590 55.885 157.590 55.860 ;
        RECT 157.590 55.860 158.640 55.885 ;
        POLYGON 157.590 55.860 157.660 55.860 157.660 55.835 ;
        RECT 157.660 55.850 158.640 55.860 ;
        POLYGON 158.640 55.915 158.745 55.850 158.640 55.850 ;
        POLYGON 159.600 55.915 159.690 55.915 159.690 55.850 ;
        RECT 159.690 55.850 160.695 55.915 ;
        RECT 157.660 55.840 158.745 55.850 ;
        POLYGON 158.745 55.850 158.765 55.840 158.745 55.840 ;
        POLYGON 159.690 55.850 159.705 55.850 159.705 55.840 ;
        RECT 159.705 55.840 160.695 55.850 ;
        RECT 157.660 55.835 158.765 55.840 ;
        POLYGON 157.665 55.835 157.670 55.835 157.670 55.830 ;
        RECT 157.670 55.830 158.765 55.835 ;
        RECT 151.790 55.825 152.715 55.830 ;
        POLYGON 152.715 55.830 152.730 55.830 152.715 55.825 ;
        POLYGON 157.670 55.830 157.680 55.830 157.680 55.825 ;
        RECT 157.680 55.825 158.765 55.830 ;
        RECT 151.790 55.820 152.695 55.825 ;
        POLYGON 151.725 55.820 151.725 55.790 151.675 55.790 ;
        RECT 151.725 55.815 152.695 55.820 ;
        POLYGON 152.695 55.825 152.715 55.825 152.695 55.815 ;
        POLYGON 157.680 55.825 157.700 55.825 157.700 55.815 ;
        RECT 157.700 55.815 158.765 55.825 ;
        RECT 151.725 55.810 152.680 55.815 ;
        POLYGON 152.680 55.815 152.690 55.815 152.680 55.810 ;
        POLYGON 157.700 55.815 157.710 55.815 157.710 55.810 ;
        RECT 157.710 55.810 158.765 55.815 ;
        RECT 151.725 55.790 152.535 55.810 ;
        POLYGON 151.675 55.790 151.675 55.740 151.595 55.740 ;
        RECT 151.675 55.750 152.535 55.790 ;
        POLYGON 152.535 55.810 152.680 55.810 152.535 55.750 ;
        POLYGON 157.710 55.810 157.780 55.810 157.780 55.780 ;
        RECT 157.780 55.780 158.765 55.810 ;
        POLYGON 157.780 55.780 157.825 55.780 157.825 55.760 ;
        RECT 157.825 55.765 158.765 55.780 ;
        POLYGON 158.765 55.840 158.885 55.765 158.765 55.765 ;
        POLYGON 159.705 55.840 159.720 55.840 159.720 55.825 ;
        RECT 159.720 55.825 160.695 55.840 ;
        POLYGON 159.720 55.825 159.775 55.825 159.775 55.785 ;
        RECT 159.775 55.785 160.695 55.825 ;
        POLYGON 159.775 55.785 159.800 55.785 159.800 55.765 ;
        RECT 159.800 55.765 160.695 55.785 ;
        POLYGON 160.695 55.915 160.860 55.765 160.695 55.765 ;
        POLYGON 162.030 55.915 162.115 55.915 162.115 55.825 ;
        RECT 162.115 55.825 163.440 55.915 ;
        POLYGON 162.115 55.825 162.170 55.825 162.170 55.770 ;
        RECT 162.170 55.810 163.440 55.825 ;
        POLYGON 163.440 55.945 163.545 55.810 163.440 55.810 ;
        POLYGON 165.195 55.945 165.220 55.945 165.220 55.905 ;
        RECT 165.220 55.935 167.180 55.945 ;
        POLYGON 167.180 56.280 167.375 55.935 167.180 55.935 ;
        POLYGON 170.060 56.280 170.200 56.280 170.200 55.995 ;
        RECT 170.200 55.995 174.425 56.280 ;
        POLYGON 170.200 55.995 170.225 55.995 170.225 55.935 ;
        RECT 170.225 55.935 174.425 55.995 ;
        RECT 165.220 55.905 167.375 55.935 ;
        POLYGON 165.220 55.905 165.280 55.905 165.280 55.815 ;
        RECT 165.280 55.860 167.375 55.905 ;
        POLYGON 167.375 55.935 167.415 55.860 167.375 55.860 ;
        POLYGON 170.225 55.935 170.255 55.935 170.255 55.865 ;
        RECT 170.255 55.860 174.425 55.935 ;
        RECT 165.280 55.810 167.415 55.860 ;
        RECT 162.170 55.765 163.545 55.810 ;
        RECT 157.825 55.760 158.885 55.765 ;
        POLYGON 155.805 55.760 155.805 55.755 155.665 55.755 ;
        RECT 155.805 55.755 155.970 55.760 ;
        POLYGON 155.970 55.760 156.080 55.755 155.970 55.755 ;
        POLYGON 157.825 55.760 157.835 55.760 157.835 55.755 ;
        RECT 157.835 55.755 158.885 55.760 ;
        POLYGON 155.635 55.755 155.635 55.750 155.555 55.750 ;
        RECT 155.635 55.750 156.085 55.755 ;
        POLYGON 156.085 55.755 156.130 55.750 156.085 55.750 ;
        POLYGON 157.835 55.755 157.850 55.755 157.850 55.750 ;
        RECT 157.850 55.750 158.885 55.755 ;
        RECT 151.675 55.740 152.505 55.750 ;
        RECT 149.560 55.730 150.615 55.740 ;
        POLYGON 150.615 55.740 150.625 55.740 150.615 55.730 ;
        POLYGON 151.595 55.740 151.595 55.735 151.585 55.735 ;
        RECT 151.595 55.735 152.505 55.740 ;
        POLYGON 152.505 55.750 152.535 55.750 152.505 55.735 ;
        POLYGON 155.545 55.750 155.545 55.745 155.460 55.745 ;
        RECT 155.545 55.745 156.155 55.750 ;
        POLYGON 155.455 55.745 155.455 55.735 155.370 55.735 ;
        RECT 155.455 55.740 156.155 55.745 ;
        POLYGON 156.155 55.750 156.265 55.740 156.155 55.740 ;
        POLYGON 157.850 55.750 157.865 55.750 157.865 55.745 ;
        RECT 157.865 55.745 158.885 55.750 ;
        POLYGON 157.865 55.745 157.875 55.745 157.875 55.740 ;
        RECT 157.875 55.740 158.885 55.745 ;
        RECT 155.455 55.735 156.295 55.740 ;
        POLYGON 151.585 55.735 151.585 55.730 151.580 55.730 ;
        RECT 151.585 55.730 152.400 55.735 ;
        RECT 149.560 55.725 150.545 55.730 ;
        RECT 147.285 55.665 148.435 55.725 ;
        POLYGON 146.555 55.665 146.560 55.660 146.555 55.660 ;
        RECT 117.290 55.610 146.560 55.660 ;
        POLYGON 147.240 55.665 147.240 55.650 147.230 55.650 ;
        RECT 147.240 55.655 148.435 55.665 ;
        POLYGON 148.435 55.725 148.495 55.725 148.435 55.655 ;
        POLYGON 149.525 55.725 149.525 55.655 149.465 55.655 ;
        RECT 149.525 55.675 150.545 55.725 ;
        POLYGON 150.545 55.730 150.615 55.730 150.545 55.675 ;
        POLYGON 151.580 55.730 151.580 55.675 151.495 55.675 ;
        RECT 151.580 55.695 152.400 55.730 ;
        POLYGON 152.400 55.735 152.505 55.735 152.400 55.695 ;
        POLYGON 155.370 55.735 155.370 55.725 155.280 55.725 ;
        RECT 155.370 55.725 156.295 55.735 ;
        POLYGON 155.250 55.725 155.250 55.715 155.175 55.715 ;
        RECT 155.250 55.720 156.295 55.725 ;
        POLYGON 156.295 55.740 156.440 55.720 156.295 55.720 ;
        POLYGON 157.875 55.740 157.915 55.740 157.915 55.720 ;
        RECT 157.915 55.720 158.885 55.740 ;
        RECT 155.250 55.715 156.450 55.720 ;
        POLYGON 155.170 55.715 155.170 55.695 155.045 55.695 ;
        RECT 155.170 55.710 156.450 55.715 ;
        POLYGON 156.450 55.720 156.510 55.710 156.450 55.710 ;
        POLYGON 157.915 55.720 157.935 55.720 157.935 55.710 ;
        RECT 157.935 55.710 158.885 55.720 ;
        POLYGON 158.885 55.765 158.965 55.710 158.885 55.710 ;
        POLYGON 159.800 55.765 159.860 55.765 159.860 55.710 ;
        RECT 159.860 55.725 160.860 55.765 ;
        POLYGON 160.860 55.765 160.905 55.725 160.860 55.725 ;
        POLYGON 162.170 55.765 162.175 55.765 162.175 55.760 ;
        RECT 162.175 55.760 163.545 55.765 ;
        POLYGON 162.175 55.760 162.205 55.760 162.205 55.725 ;
        RECT 162.205 55.725 163.545 55.760 ;
        RECT 159.860 55.710 160.905 55.725 ;
        RECT 155.170 55.695 156.510 55.710 ;
        POLYGON 156.510 55.710 156.590 55.695 156.510 55.695 ;
        POLYGON 157.935 55.710 157.965 55.710 157.965 55.695 ;
        RECT 157.965 55.700 158.965 55.710 ;
        POLYGON 158.965 55.710 158.990 55.700 158.965 55.700 ;
        POLYGON 159.860 55.710 159.875 55.710 159.875 55.700 ;
        RECT 159.875 55.700 160.905 55.710 ;
        RECT 157.965 55.695 158.990 55.700 ;
        RECT 151.580 55.675 152.290 55.695 ;
        RECT 149.525 55.670 150.540 55.675 ;
        POLYGON 150.540 55.675 150.545 55.675 150.540 55.670 ;
        POLYGON 151.495 55.675 151.495 55.670 151.490 55.670 ;
        RECT 151.495 55.670 152.290 55.675 ;
        RECT 149.525 55.655 150.425 55.670 ;
        RECT 147.240 55.650 148.405 55.655 ;
        RECT 51.940 54.190 111.225 55.610 ;
        POLYGON 111.225 55.610 111.320 54.190 111.225 54.190 ;
        POLYGON 117.275 55.595 117.275 54.260 117.250 54.260 ;
        RECT 117.275 55.515 146.560 55.610 ;
        POLYGON 146.560 55.650 146.600 55.515 146.560 55.515 ;
        RECT 117.275 55.460 146.600 55.515 ;
        POLYGON 147.230 55.650 147.230 55.510 147.130 55.510 ;
        RECT 147.230 55.615 148.405 55.650 ;
        POLYGON 148.405 55.655 148.435 55.655 148.405 55.615 ;
        POLYGON 149.465 55.655 149.465 55.620 149.435 55.620 ;
        RECT 149.465 55.620 150.425 55.655 ;
        POLYGON 149.435 55.620 149.435 55.615 149.430 55.615 ;
        RECT 149.435 55.615 150.425 55.620 ;
        RECT 147.230 55.570 148.370 55.615 ;
        POLYGON 148.370 55.615 148.405 55.615 148.370 55.570 ;
        POLYGON 149.430 55.615 149.430 55.575 149.390 55.575 ;
        RECT 149.430 55.575 150.425 55.615 ;
        POLYGON 150.425 55.670 150.540 55.670 150.425 55.575 ;
        POLYGON 151.485 55.670 151.485 55.575 151.345 55.575 ;
        RECT 151.485 55.640 152.290 55.670 ;
        POLYGON 152.290 55.695 152.400 55.695 152.290 55.640 ;
        POLYGON 155.035 55.695 155.035 55.690 155.010 55.690 ;
        RECT 155.035 55.690 156.605 55.695 ;
        POLYGON 155.000 55.690 155.000 55.680 154.910 55.680 ;
        RECT 155.000 55.680 156.605 55.690 ;
        POLYGON 154.910 55.680 154.910 55.655 154.785 55.655 ;
        RECT 154.910 55.670 156.605 55.680 ;
        POLYGON 156.605 55.695 156.715 55.670 156.605 55.670 ;
        POLYGON 157.965 55.695 158.010 55.695 158.010 55.670 ;
        RECT 158.010 55.680 158.990 55.695 ;
        POLYGON 158.990 55.700 159.015 55.680 158.990 55.680 ;
        POLYGON 159.875 55.700 159.895 55.700 159.895 55.680 ;
        RECT 159.895 55.685 160.905 55.700 ;
        POLYGON 160.905 55.725 160.940 55.685 160.905 55.685 ;
        POLYGON 162.205 55.725 162.210 55.725 162.210 55.720 ;
        RECT 162.210 55.720 163.545 55.725 ;
        POLYGON 162.210 55.720 162.235 55.720 162.235 55.690 ;
        RECT 162.235 55.685 163.545 55.720 ;
        RECT 159.895 55.680 160.940 55.685 ;
        RECT 158.010 55.670 159.015 55.680 ;
        RECT 154.910 55.660 156.725 55.670 ;
        POLYGON 156.725 55.670 156.745 55.660 156.725 55.660 ;
        POLYGON 158.010 55.670 158.030 55.670 158.030 55.660 ;
        RECT 158.030 55.660 159.015 55.670 ;
        RECT 154.910 55.655 156.745 55.660 ;
        POLYGON 154.785 55.655 154.785 55.640 154.715 55.640 ;
        RECT 154.785 55.640 156.745 55.655 ;
        RECT 151.485 55.580 152.165 55.640 ;
        POLYGON 152.165 55.640 152.290 55.640 152.165 55.580 ;
        POLYGON 154.715 55.640 154.715 55.625 154.640 55.625 ;
        RECT 154.715 55.635 156.745 55.640 ;
        POLYGON 156.745 55.660 156.845 55.635 156.745 55.635 ;
        POLYGON 158.030 55.660 158.075 55.660 158.075 55.635 ;
        RECT 158.075 55.635 159.015 55.660 ;
        RECT 154.715 55.625 156.845 55.635 ;
        POLYGON 154.640 55.625 154.640 55.610 154.570 55.610 ;
        RECT 154.640 55.610 156.845 55.625 ;
        POLYGON 156.845 55.635 156.925 55.610 156.845 55.610 ;
        POLYGON 158.075 55.635 158.125 55.635 158.125 55.610 ;
        RECT 158.125 55.610 159.015 55.635 ;
        POLYGON 154.565 55.610 154.565 55.605 154.530 55.605 ;
        RECT 154.565 55.605 156.925 55.610 ;
        POLYGON 156.925 55.610 156.935 55.605 156.925 55.605 ;
        POLYGON 158.130 55.610 158.135 55.610 158.135 55.605 ;
        RECT 158.135 55.605 159.015 55.610 ;
        POLYGON 159.015 55.680 159.125 55.605 159.015 55.605 ;
        POLYGON 159.895 55.680 159.935 55.680 159.935 55.650 ;
        RECT 159.935 55.650 160.940 55.680 ;
        POLYGON 160.940 55.685 160.975 55.650 160.940 55.650 ;
        POLYGON 162.235 55.685 162.265 55.685 162.265 55.650 ;
        RECT 162.265 55.650 163.545 55.685 ;
        POLYGON 163.545 55.810 163.665 55.650 163.545 55.650 ;
        POLYGON 165.280 55.810 165.290 55.810 165.290 55.800 ;
        RECT 165.290 55.800 167.415 55.810 ;
        POLYGON 165.290 55.800 165.300 55.800 165.300 55.785 ;
        RECT 165.300 55.785 167.415 55.800 ;
        POLYGON 165.300 55.785 165.325 55.785 165.325 55.740 ;
        RECT 165.325 55.740 167.415 55.785 ;
        POLYGON 165.325 55.740 165.375 55.740 165.375 55.655 ;
        RECT 165.375 55.650 167.415 55.740 ;
        POLYGON 159.940 55.650 159.985 55.650 159.985 55.605 ;
        RECT 159.985 55.605 160.975 55.650 ;
        POLYGON 154.530 55.605 154.530 55.600 154.505 55.600 ;
        RECT 154.530 55.600 156.940 55.605 ;
        POLYGON 154.500 55.600 154.500 55.580 154.430 55.580 ;
        RECT 154.500 55.595 156.940 55.600 ;
        POLYGON 156.940 55.605 156.975 55.595 156.940 55.595 ;
        POLYGON 158.135 55.605 158.155 55.605 158.155 55.595 ;
        RECT 158.155 55.595 159.125 55.605 ;
        RECT 154.500 55.580 156.975 55.595 ;
        RECT 151.485 55.575 152.135 55.580 ;
        RECT 147.230 55.510 148.195 55.570 ;
        POLYGON 146.600 55.510 146.615 55.460 146.600 55.460 ;
        RECT 117.275 55.385 146.615 55.460 ;
        POLYGON 147.130 55.510 147.130 55.450 147.090 55.450 ;
        RECT 147.130 55.450 148.195 55.510 ;
        POLYGON 146.615 55.450 146.635 55.385 146.615 55.385 ;
        RECT 117.275 55.335 146.635 55.385 ;
        POLYGON 147.090 55.450 147.090 55.385 147.040 55.385 ;
        RECT 147.090 55.385 148.195 55.450 ;
        POLYGON 147.040 55.380 147.040 55.375 147.035 55.375 ;
        RECT 147.040 55.375 148.195 55.385 ;
        POLYGON 146.635 55.375 146.650 55.335 146.635 55.335 ;
        RECT 117.275 55.315 146.650 55.335 ;
        POLYGON 147.035 55.375 147.035 55.320 147.000 55.320 ;
        RECT 147.035 55.340 148.195 55.375 ;
        POLYGON 148.195 55.570 148.370 55.570 148.195 55.340 ;
        POLYGON 149.390 55.570 149.390 55.525 149.345 55.525 ;
        RECT 149.390 55.525 150.325 55.575 ;
        POLYGON 149.345 55.525 149.345 55.465 149.295 55.465 ;
        RECT 149.345 55.485 150.325 55.525 ;
        POLYGON 150.325 55.575 150.425 55.575 150.325 55.485 ;
        POLYGON 151.345 55.575 151.345 55.535 151.285 55.535 ;
        RECT 151.345 55.565 152.135 55.575 ;
        POLYGON 152.135 55.580 152.165 55.580 152.135 55.565 ;
        POLYGON 154.430 55.580 154.430 55.565 154.370 55.565 ;
        RECT 154.430 55.575 156.975 55.580 ;
        POLYGON 156.975 55.595 157.030 55.575 156.975 55.575 ;
        POLYGON 158.155 55.595 158.185 55.595 158.185 55.580 ;
        RECT 158.185 55.580 159.125 55.595 ;
        POLYGON 158.185 55.580 158.190 55.580 158.190 55.575 ;
        RECT 158.190 55.575 159.125 55.580 ;
        RECT 154.430 55.565 157.030 55.575 ;
        RECT 151.345 55.535 151.985 55.565 ;
        POLYGON 151.285 55.535 151.285 55.515 151.265 55.515 ;
        RECT 151.285 55.515 151.985 55.535 ;
        POLYGON 151.265 55.515 151.265 55.505 151.245 55.505 ;
        RECT 151.265 55.505 151.985 55.515 ;
        POLYGON 151.245 55.505 151.245 55.485 151.220 55.485 ;
        RECT 151.245 55.485 151.985 55.505 ;
        POLYGON 151.985 55.565 152.135 55.565 151.985 55.485 ;
        POLYGON 154.370 55.565 154.370 55.560 154.350 55.560 ;
        RECT 154.370 55.560 157.030 55.565 ;
        POLYGON 154.345 55.560 154.345 55.530 154.220 55.530 ;
        RECT 154.345 55.530 157.030 55.560 ;
        POLYGON 157.030 55.575 157.150 55.530 157.030 55.530 ;
        POLYGON 158.190 55.575 158.230 55.575 158.230 55.555 ;
        RECT 158.230 55.555 159.125 55.575 ;
        POLYGON 158.230 55.555 158.245 55.555 158.245 55.545 ;
        RECT 158.245 55.545 159.125 55.555 ;
        POLYGON 158.245 55.545 158.270 55.545 158.270 55.530 ;
        RECT 158.270 55.530 159.125 55.545 ;
        POLYGON 159.125 55.605 159.225 55.530 159.125 55.530 ;
        POLYGON 159.985 55.605 160.005 55.605 160.005 55.590 ;
        RECT 160.005 55.590 160.975 55.605 ;
        POLYGON 160.005 55.590 160.075 55.590 160.075 55.530 ;
        RECT 160.075 55.530 160.975 55.590 ;
        POLYGON 154.215 55.530 154.215 55.520 154.180 55.520 ;
        RECT 154.215 55.520 157.150 55.530 ;
        POLYGON 154.180 55.520 154.180 55.510 154.140 55.510 ;
        RECT 154.180 55.510 157.150 55.520 ;
        POLYGON 154.130 55.510 154.130 55.485 154.050 55.485 ;
        RECT 154.130 55.505 157.150 55.510 ;
        RECT 154.130 55.500 155.465 55.505 ;
        POLYGON 155.465 55.505 155.570 55.505 155.465 55.500 ;
        POLYGON 155.805 55.505 155.820 55.505 155.820 55.500 ;
        RECT 155.820 55.500 157.150 55.505 ;
        RECT 154.130 55.495 155.385 55.500 ;
        POLYGON 155.385 55.500 155.445 55.500 155.385 55.495 ;
        POLYGON 155.875 55.500 155.930 55.500 155.930 55.495 ;
        RECT 155.930 55.495 157.150 55.500 ;
        POLYGON 157.150 55.530 157.235 55.495 157.150 55.495 ;
        POLYGON 158.270 55.530 158.325 55.530 158.325 55.495 ;
        RECT 158.325 55.510 159.230 55.530 ;
        POLYGON 159.230 55.530 159.260 55.510 159.230 55.510 ;
        POLYGON 160.075 55.530 160.095 55.530 160.095 55.510 ;
        RECT 160.095 55.510 160.975 55.530 ;
        RECT 158.325 55.495 159.260 55.510 ;
        RECT 154.130 55.485 155.280 55.495 ;
        RECT 149.345 55.470 150.305 55.485 ;
        POLYGON 150.305 55.485 150.325 55.485 150.305 55.470 ;
        POLYGON 151.220 55.485 151.220 55.470 151.200 55.470 ;
        RECT 151.220 55.470 151.940 55.485 ;
        RECT 149.345 55.465 150.235 55.470 ;
        POLYGON 149.295 55.465 149.295 55.385 149.220 55.385 ;
        RECT 149.295 55.405 150.235 55.465 ;
        POLYGON 150.235 55.470 150.305 55.470 150.235 55.405 ;
        POLYGON 151.200 55.470 151.200 55.405 151.115 55.405 ;
        RECT 151.200 55.460 151.940 55.470 ;
        POLYGON 151.940 55.485 151.985 55.485 151.940 55.460 ;
        POLYGON 154.050 55.485 154.050 55.470 154.005 55.470 ;
        RECT 154.050 55.480 155.280 55.485 ;
        POLYGON 155.280 55.495 155.370 55.495 155.280 55.480 ;
        POLYGON 155.935 55.495 155.950 55.495 155.950 55.490 ;
        RECT 155.950 55.490 157.235 55.495 ;
        POLYGON 155.970 55.490 156.025 55.490 156.025 55.480 ;
        RECT 156.025 55.480 157.235 55.490 ;
        RECT 154.050 55.470 155.205 55.480 ;
        POLYGON 155.205 55.480 155.270 55.480 155.205 55.470 ;
        POLYGON 156.025 55.480 156.085 55.480 156.085 55.470 ;
        RECT 156.085 55.470 157.235 55.480 ;
        POLYGON 154.005 55.470 154.005 55.460 153.970 55.460 ;
        RECT 154.005 55.460 155.130 55.470 ;
        RECT 151.200 55.425 151.880 55.460 ;
        POLYGON 151.880 55.460 151.940 55.460 151.880 55.425 ;
        POLYGON 153.970 55.460 153.970 55.445 153.915 55.445 ;
        RECT 153.970 55.455 155.130 55.460 ;
        POLYGON 155.130 55.470 155.195 55.470 155.130 55.455 ;
        POLYGON 156.085 55.470 156.115 55.470 156.115 55.465 ;
        RECT 156.115 55.465 157.235 55.470 ;
        POLYGON 156.135 55.465 156.180 55.465 156.180 55.455 ;
        RECT 156.180 55.460 157.235 55.465 ;
        POLYGON 157.235 55.495 157.315 55.460 157.235 55.460 ;
        POLYGON 158.325 55.495 158.380 55.495 158.380 55.465 ;
        RECT 158.380 55.465 159.260 55.495 ;
        POLYGON 158.380 55.465 158.385 55.465 158.385 55.460 ;
        RECT 158.385 55.460 159.260 55.465 ;
        RECT 156.180 55.455 157.315 55.460 ;
        RECT 153.970 55.445 155.070 55.455 ;
        POLYGON 153.915 55.445 153.915 55.430 153.865 55.430 ;
        RECT 153.915 55.440 155.070 55.445 ;
        POLYGON 155.070 55.455 155.125 55.455 155.070 55.440 ;
        POLYGON 156.180 55.455 156.225 55.455 156.225 55.445 ;
        RECT 156.225 55.445 157.315 55.455 ;
        POLYGON 156.225 55.445 156.245 55.445 156.245 55.440 ;
        RECT 156.245 55.440 157.315 55.445 ;
        POLYGON 157.315 55.460 157.365 55.440 157.315 55.440 ;
        POLYGON 158.385 55.460 158.415 55.460 158.415 55.440 ;
        RECT 158.415 55.440 159.260 55.460 ;
        RECT 153.915 55.435 155.060 55.440 ;
        POLYGON 155.060 55.440 155.070 55.440 155.060 55.435 ;
        POLYGON 156.245 55.440 156.265 55.440 156.265 55.435 ;
        RECT 156.265 55.435 157.365 55.440 ;
        RECT 153.915 55.430 155.020 55.435 ;
        POLYGON 153.865 55.430 153.865 55.425 153.850 55.425 ;
        RECT 153.865 55.425 155.020 55.430 ;
        POLYGON 155.020 55.435 155.060 55.435 155.020 55.425 ;
        POLYGON 156.265 55.435 156.285 55.435 156.285 55.430 ;
        RECT 156.285 55.430 157.365 55.435 ;
        POLYGON 157.365 55.440 157.385 55.430 157.365 55.430 ;
        POLYGON 158.415 55.440 158.430 55.440 158.430 55.430 ;
        RECT 158.430 55.435 159.260 55.440 ;
        POLYGON 159.260 55.510 159.355 55.435 159.260 55.435 ;
        POLYGON 160.095 55.510 160.145 55.510 160.145 55.470 ;
        RECT 160.145 55.470 160.975 55.510 ;
        POLYGON 160.145 55.470 160.165 55.470 160.165 55.460 ;
        RECT 160.165 55.455 160.975 55.470 ;
        POLYGON 160.165 55.455 160.185 55.455 160.185 55.435 ;
        RECT 160.185 55.440 160.975 55.455 ;
        POLYGON 160.975 55.650 161.180 55.440 160.975 55.440 ;
        POLYGON 162.265 55.650 162.365 55.650 162.365 55.535 ;
        RECT 162.365 55.625 163.665 55.650 ;
        POLYGON 163.665 55.650 163.685 55.625 163.665 55.625 ;
        POLYGON 165.375 55.650 165.385 55.650 165.385 55.640 ;
        RECT 165.385 55.640 167.415 55.650 ;
        POLYGON 165.385 55.640 165.390 55.640 165.390 55.630 ;
        RECT 165.390 55.625 167.415 55.640 ;
        RECT 162.365 55.555 163.685 55.625 ;
        POLYGON 163.685 55.625 163.735 55.555 163.685 55.555 ;
        POLYGON 165.390 55.625 165.400 55.625 165.400 55.610 ;
        RECT 165.400 55.610 167.415 55.625 ;
        POLYGON 165.400 55.610 165.430 55.610 165.430 55.555 ;
        RECT 165.430 55.555 167.415 55.610 ;
        RECT 162.365 55.535 163.735 55.555 ;
        POLYGON 162.365 55.535 162.410 55.535 162.410 55.475 ;
        RECT 162.410 55.475 163.735 55.535 ;
        POLYGON 162.410 55.475 162.435 55.475 162.435 55.440 ;
        RECT 162.435 55.440 163.735 55.475 ;
        RECT 160.185 55.435 161.180 55.440 ;
        RECT 158.430 55.430 159.355 55.435 ;
        POLYGON 156.300 55.430 156.320 55.430 156.320 55.425 ;
        RECT 156.320 55.425 157.385 55.430 ;
        RECT 151.200 55.405 151.810 55.425 ;
        RECT 149.295 55.385 150.190 55.405 ;
        POLYGON 149.220 55.385 149.220 55.340 149.185 55.340 ;
        RECT 149.220 55.365 150.190 55.385 ;
        POLYGON 150.190 55.405 150.235 55.405 150.190 55.365 ;
        POLYGON 151.115 55.405 151.115 55.365 151.060 55.365 ;
        RECT 151.115 55.385 151.810 55.405 ;
        POLYGON 151.810 55.425 151.875 55.425 151.810 55.385 ;
        POLYGON 153.850 55.425 153.850 55.410 153.795 55.410 ;
        RECT 153.850 55.420 155.015 55.425 ;
        POLYGON 155.015 55.425 155.020 55.425 155.015 55.420 ;
        POLYGON 156.320 55.425 156.340 55.425 156.340 55.420 ;
        RECT 156.340 55.420 157.385 55.425 ;
        RECT 153.850 55.410 154.970 55.420 ;
        POLYGON 153.790 55.410 153.790 55.395 153.740 55.395 ;
        RECT 153.790 55.400 154.970 55.410 ;
        POLYGON 154.970 55.420 155.010 55.420 154.970 55.400 ;
        POLYGON 156.340 55.420 156.365 55.420 156.365 55.415 ;
        RECT 156.365 55.415 157.385 55.420 ;
        POLYGON 156.365 55.415 156.410 55.415 156.410 55.400 ;
        RECT 156.410 55.400 157.385 55.415 ;
        RECT 153.790 55.395 154.965 55.400 ;
        POLYGON 154.965 55.400 154.970 55.400 154.965 55.395 ;
        POLYGON 156.410 55.400 156.425 55.400 156.425 55.395 ;
        RECT 156.425 55.395 157.385 55.400 ;
        POLYGON 153.735 55.395 153.735 55.385 153.705 55.385 ;
        RECT 153.735 55.385 154.925 55.395 ;
        RECT 151.115 55.365 151.640 55.385 ;
        RECT 149.220 55.340 150.075 55.365 ;
        RECT 147.035 55.320 148.175 55.340 ;
        POLYGON 146.650 55.320 146.655 55.315 146.650 55.315 ;
        RECT 117.275 55.245 146.655 55.315 ;
        POLYGON 147.000 55.320 147.000 55.305 146.990 55.305 ;
        RECT 147.000 55.315 148.175 55.320 ;
        POLYGON 148.175 55.340 148.195 55.340 148.175 55.315 ;
        POLYGON 149.185 55.340 149.185 55.315 149.165 55.315 ;
        RECT 149.185 55.315 150.075 55.340 ;
        RECT 147.000 55.305 148.130 55.315 ;
        POLYGON 146.655 55.305 146.675 55.245 146.655 55.245 ;
        RECT 117.275 55.150 146.675 55.245 ;
        POLYGON 146.990 55.305 146.990 55.235 146.945 55.235 ;
        RECT 146.990 55.245 148.130 55.305 ;
        POLYGON 148.130 55.315 148.175 55.315 148.130 55.245 ;
        POLYGON 149.165 55.315 149.165 55.280 149.140 55.280 ;
        RECT 149.165 55.280 150.075 55.315 ;
        POLYGON 149.140 55.280 149.140 55.245 149.110 55.245 ;
        RECT 149.140 55.255 150.075 55.280 ;
        POLYGON 150.075 55.365 150.190 55.365 150.075 55.255 ;
        POLYGON 151.060 55.365 151.060 55.350 151.040 55.350 ;
        RECT 151.060 55.350 151.640 55.365 ;
        POLYGON 151.040 55.350 151.040 55.325 151.010 55.325 ;
        RECT 151.040 55.325 151.640 55.350 ;
        POLYGON 151.010 55.325 151.010 55.255 150.920 55.255 ;
        RECT 151.010 55.280 151.640 55.325 ;
        POLYGON 151.640 55.385 151.810 55.385 151.640 55.280 ;
        POLYGON 153.705 55.385 153.705 55.340 153.580 55.340 ;
        RECT 153.705 55.375 154.925 55.385 ;
        POLYGON 154.925 55.395 154.965 55.395 154.925 55.375 ;
        POLYGON 156.425 55.395 156.440 55.395 156.440 55.390 ;
        RECT 156.440 55.390 157.385 55.395 ;
        POLYGON 156.440 55.390 156.480 55.390 156.480 55.380 ;
        RECT 156.480 55.380 157.385 55.390 ;
        POLYGON 156.480 55.380 156.505 55.380 156.505 55.375 ;
        RECT 156.505 55.375 157.385 55.380 ;
        RECT 153.705 55.350 154.900 55.375 ;
        POLYGON 154.900 55.375 154.925 55.375 154.900 55.350 ;
        POLYGON 156.505 55.375 156.585 55.375 156.585 55.350 ;
        RECT 156.585 55.360 157.385 55.375 ;
        POLYGON 157.385 55.430 157.535 55.360 157.385 55.360 ;
        POLYGON 158.430 55.430 158.510 55.430 158.510 55.380 ;
        RECT 158.510 55.425 159.355 55.430 ;
        POLYGON 159.355 55.435 159.375 55.425 159.355 55.425 ;
        POLYGON 160.185 55.435 160.195 55.435 160.195 55.425 ;
        RECT 160.195 55.425 161.180 55.435 ;
        RECT 158.510 55.380 159.375 55.425 ;
        POLYGON 158.510 55.380 158.540 55.380 158.540 55.360 ;
        RECT 158.540 55.360 159.375 55.380 ;
        RECT 156.585 55.350 157.535 55.360 ;
        RECT 153.705 55.340 154.885 55.350 ;
        POLYGON 153.580 55.340 153.580 55.330 153.555 55.330 ;
        RECT 153.580 55.330 154.885 55.340 ;
        POLYGON 154.885 55.350 154.900 55.350 154.885 55.330 ;
        POLYGON 156.590 55.350 156.595 55.350 156.595 55.345 ;
        RECT 156.595 55.345 157.535 55.350 ;
        POLYGON 156.595 55.345 156.650 55.345 156.650 55.330 ;
        RECT 156.650 55.330 157.535 55.345 ;
        POLYGON 157.535 55.360 157.590 55.330 157.535 55.330 ;
        POLYGON 158.540 55.360 158.580 55.360 158.580 55.335 ;
        RECT 158.580 55.335 159.375 55.360 ;
        POLYGON 158.580 55.335 158.585 55.335 158.585 55.330 ;
        RECT 158.585 55.330 159.375 55.335 ;
        POLYGON 153.555 55.330 153.555 55.325 153.530 55.325 ;
        RECT 153.555 55.325 154.880 55.330 ;
        POLYGON 154.880 55.330 154.885 55.330 154.880 55.325 ;
        POLYGON 156.650 55.330 156.660 55.330 156.660 55.325 ;
        RECT 156.660 55.325 157.590 55.330 ;
        POLYGON 153.530 55.325 153.530 55.310 153.495 55.310 ;
        RECT 153.530 55.310 154.870 55.325 ;
        POLYGON 154.870 55.325 154.880 55.325 154.870 55.310 ;
        POLYGON 156.660 55.325 156.700 55.325 156.700 55.310 ;
        RECT 156.700 55.310 157.590 55.325 ;
        POLYGON 153.495 55.310 153.495 55.280 153.415 55.280 ;
        RECT 153.495 55.305 154.870 55.310 ;
        POLYGON 156.700 55.310 156.715 55.310 156.715 55.305 ;
        RECT 156.715 55.305 157.590 55.310 ;
        RECT 153.495 55.280 154.865 55.305 ;
        POLYGON 154.865 55.305 154.870 55.305 154.865 55.295 ;
        POLYGON 156.715 55.305 156.750 55.305 156.750 55.295 ;
        RECT 156.750 55.295 157.590 55.305 ;
        POLYGON 157.590 55.330 157.665 55.295 157.590 55.295 ;
        POLYGON 158.585 55.330 158.630 55.330 158.630 55.295 ;
        RECT 158.630 55.325 159.375 55.330 ;
        POLYGON 159.375 55.425 159.495 55.325 159.375 55.325 ;
        POLYGON 160.195 55.425 160.205 55.425 160.205 55.420 ;
        RECT 160.205 55.420 161.180 55.425 ;
        POLYGON 160.205 55.420 160.305 55.420 160.305 55.325 ;
        RECT 160.305 55.405 161.180 55.420 ;
        POLYGON 161.180 55.440 161.210 55.405 161.180 55.405 ;
        POLYGON 162.435 55.440 162.465 55.440 162.465 55.405 ;
        RECT 162.465 55.415 163.735 55.440 ;
        POLYGON 163.735 55.555 163.830 55.415 163.735 55.415 ;
        POLYGON 165.430 55.555 165.445 55.555 165.445 55.530 ;
        RECT 165.445 55.530 167.415 55.555 ;
        POLYGON 165.445 55.530 165.475 55.530 165.475 55.485 ;
        RECT 165.475 55.485 167.415 55.530 ;
        POLYGON 165.475 55.485 165.485 55.485 165.485 55.465 ;
        RECT 165.485 55.465 167.415 55.485 ;
        POLYGON 167.415 55.860 167.620 55.465 167.415 55.465 ;
        POLYGON 170.255 55.860 170.430 55.860 170.430 55.465 ;
        RECT 170.430 55.465 174.425 55.860 ;
        POLYGON 165.485 55.465 165.490 55.465 165.490 55.460 ;
        RECT 165.490 55.455 167.620 55.465 ;
        POLYGON 165.490 55.455 165.500 55.455 165.500 55.440 ;
        RECT 165.500 55.440 167.620 55.455 ;
        POLYGON 165.500 55.440 165.510 55.440 165.510 55.420 ;
        RECT 165.510 55.430 167.620 55.440 ;
        POLYGON 167.620 55.465 167.635 55.430 167.620 55.430 ;
        POLYGON 170.430 55.465 170.445 55.465 170.445 55.430 ;
        RECT 170.445 55.430 174.425 55.465 ;
        RECT 165.510 55.415 167.635 55.430 ;
        RECT 162.465 55.405 163.830 55.415 ;
        RECT 160.305 55.375 161.210 55.405 ;
        POLYGON 161.210 55.405 161.240 55.375 161.210 55.375 ;
        POLYGON 162.465 55.405 162.485 55.405 162.485 55.380 ;
        RECT 162.485 55.375 163.830 55.405 ;
        RECT 160.305 55.325 161.240 55.375 ;
        RECT 158.630 55.295 159.495 55.325 ;
        RECT 151.010 55.275 151.630 55.280 ;
        POLYGON 151.630 55.280 151.640 55.280 151.630 55.275 ;
        POLYGON 153.415 55.280 153.415 55.275 153.405 55.275 ;
        RECT 153.415 55.275 154.865 55.280 ;
        POLYGON 156.750 55.295 156.795 55.295 156.795 55.275 ;
        RECT 156.795 55.285 157.665 55.295 ;
        POLYGON 157.665 55.295 157.680 55.285 157.665 55.285 ;
        POLYGON 158.630 55.295 158.650 55.295 158.650 55.285 ;
        RECT 158.650 55.285 159.495 55.295 ;
        RECT 156.795 55.275 157.680 55.285 ;
        RECT 151.010 55.255 151.585 55.275 ;
        RECT 149.140 55.245 149.875 55.255 ;
        RECT 146.990 55.235 148.120 55.245 ;
        POLYGON 146.675 55.235 146.700 55.150 146.675 55.150 ;
        POLYGON 146.945 55.235 146.945 55.150 146.890 55.150 ;
        RECT 146.945 55.230 148.120 55.235 ;
        POLYGON 148.120 55.245 148.130 55.245 148.120 55.230 ;
        POLYGON 149.110 55.245 149.110 55.230 149.095 55.230 ;
        RECT 149.110 55.230 149.875 55.245 ;
        RECT 146.945 55.150 148.030 55.230 ;
        RECT 117.275 55.115 146.700 55.150 ;
        POLYGON 146.700 55.150 146.710 55.115 146.700 55.115 ;
        RECT 117.275 55.080 146.710 55.115 ;
        POLYGON 146.890 55.150 146.890 55.110 146.865 55.110 ;
        RECT 146.890 55.110 148.030 55.150 ;
        POLYGON 148.030 55.230 148.120 55.230 148.030 55.110 ;
        POLYGON 149.095 55.230 149.095 55.225 149.090 55.225 ;
        RECT 149.095 55.225 149.875 55.230 ;
        POLYGON 149.090 55.225 149.090 55.110 149.000 55.110 ;
        RECT 149.090 55.110 149.875 55.225 ;
        POLYGON 146.710 55.105 146.720 55.080 146.710 55.080 ;
        RECT 117.275 55.025 146.720 55.080 ;
        POLYGON 146.865 55.105 146.865 55.070 146.840 55.070 ;
        RECT 146.865 55.100 148.025 55.110 ;
        POLYGON 148.025 55.110 148.030 55.110 148.025 55.100 ;
        POLYGON 149.000 55.110 149.000 55.100 148.990 55.100 ;
        RECT 149.000 55.100 149.875 55.110 ;
        RECT 146.865 55.070 147.900 55.100 ;
        POLYGON 146.720 55.070 146.735 55.025 146.720 55.025 ;
        RECT 117.275 54.955 146.735 55.025 ;
        POLYGON 146.840 55.070 146.840 55.015 146.805 55.015 ;
        RECT 146.840 55.015 147.900 55.070 ;
        POLYGON 146.735 55.015 146.755 54.955 146.735 54.955 ;
        RECT 117.275 54.940 146.755 54.955 ;
        POLYGON 146.805 55.015 146.805 54.945 146.765 54.945 ;
        RECT 146.805 54.945 147.900 55.015 ;
        POLYGON 146.765 54.945 146.765 54.940 146.760 54.940 ;
        RECT 146.765 54.940 147.900 54.945 ;
        RECT 117.275 54.910 147.900 54.940 ;
        POLYGON 147.900 55.100 148.025 55.100 147.900 54.910 ;
        POLYGON 148.990 55.100 148.990 55.030 148.935 55.030 ;
        RECT 148.990 55.055 149.875 55.100 ;
        POLYGON 149.875 55.255 150.075 55.255 149.875 55.055 ;
        POLYGON 150.920 55.255 150.920 55.245 150.910 55.245 ;
        RECT 150.920 55.245 151.585 55.255 ;
        POLYGON 151.585 55.275 151.630 55.275 151.585 55.245 ;
        POLYGON 153.405 55.275 153.405 55.245 153.325 55.245 ;
        RECT 153.405 55.245 154.865 55.275 ;
        POLYGON 156.795 55.275 156.840 55.275 156.840 55.260 ;
        RECT 156.840 55.260 157.680 55.275 ;
        POLYGON 156.840 55.260 156.845 55.260 156.845 55.255 ;
        RECT 156.845 55.255 157.680 55.260 ;
        POLYGON 156.845 55.255 156.855 55.255 156.855 55.250 ;
        RECT 156.855 55.250 157.680 55.255 ;
        POLYGON 150.910 55.245 150.910 55.175 150.830 55.175 ;
        RECT 150.910 55.175 151.475 55.245 ;
        POLYGON 150.830 55.175 150.830 55.130 150.770 55.130 ;
        RECT 150.830 55.165 151.475 55.175 ;
        POLYGON 151.475 55.245 151.585 55.245 151.475 55.165 ;
        POLYGON 153.325 55.245 153.325 55.215 153.255 55.215 ;
        RECT 153.325 55.235 154.865 55.245 ;
        POLYGON 154.865 55.250 154.870 55.235 154.865 55.235 ;
        POLYGON 156.855 55.250 156.890 55.250 156.890 55.235 ;
        RECT 156.890 55.235 157.680 55.250 ;
        RECT 153.325 55.220 154.870 55.235 ;
        POLYGON 154.870 55.235 154.880 55.220 154.870 55.220 ;
        POLYGON 156.890 55.235 156.905 55.235 156.905 55.230 ;
        RECT 156.905 55.230 157.680 55.235 ;
        POLYGON 157.680 55.285 157.780 55.230 157.680 55.230 ;
        POLYGON 158.650 55.285 158.720 55.285 158.720 55.230 ;
        RECT 158.720 55.255 159.495 55.285 ;
        POLYGON 159.495 55.325 159.580 55.255 159.495 55.255 ;
        POLYGON 160.305 55.325 160.345 55.325 160.345 55.290 ;
        RECT 160.345 55.300 161.240 55.325 ;
        POLYGON 161.240 55.375 161.305 55.300 161.240 55.300 ;
        POLYGON 162.485 55.375 162.525 55.375 162.525 55.330 ;
        RECT 162.525 55.330 163.830 55.375 ;
        POLYGON 162.525 55.330 162.545 55.330 162.545 55.300 ;
        RECT 162.545 55.300 163.830 55.330 ;
        RECT 160.345 55.290 161.305 55.300 ;
        POLYGON 160.345 55.290 160.380 55.290 160.380 55.255 ;
        RECT 160.380 55.255 161.305 55.290 ;
        RECT 158.720 55.230 159.580 55.255 ;
        POLYGON 156.905 55.230 156.930 55.230 156.930 55.220 ;
        RECT 156.930 55.220 157.780 55.230 ;
        RECT 153.325 55.215 154.880 55.220 ;
        POLYGON 153.255 55.215 153.255 55.165 153.145 55.165 ;
        RECT 153.255 55.205 154.880 55.215 ;
        POLYGON 154.880 55.220 154.885 55.205 154.880 55.205 ;
        POLYGON 156.930 55.220 156.975 55.220 156.975 55.205 ;
        RECT 156.975 55.205 157.780 55.220 ;
        POLYGON 157.780 55.230 157.825 55.205 157.780 55.205 ;
        POLYGON 158.720 55.230 158.750 55.230 158.750 55.205 ;
        RECT 158.750 55.205 159.580 55.230 ;
        RECT 153.255 55.185 154.885 55.205 ;
        POLYGON 154.885 55.205 154.900 55.185 154.885 55.185 ;
        POLYGON 156.975 55.205 157.020 55.205 157.020 55.185 ;
        RECT 157.020 55.185 157.825 55.205 ;
        RECT 153.255 55.175 154.900 55.185 ;
        POLYGON 154.900 55.185 154.905 55.175 154.900 55.175 ;
        POLYGON 157.020 55.185 157.045 55.185 157.045 55.175 ;
        RECT 157.045 55.180 157.825 55.185 ;
        POLYGON 157.825 55.205 157.865 55.180 157.825 55.180 ;
        POLYGON 158.750 55.205 158.785 55.205 158.785 55.180 ;
        RECT 158.785 55.180 159.580 55.205 ;
        RECT 157.045 55.175 157.865 55.180 ;
        RECT 153.255 55.165 154.905 55.175 ;
        RECT 150.830 55.160 151.465 55.165 ;
        POLYGON 151.465 55.165 151.475 55.165 151.465 55.160 ;
        POLYGON 153.145 55.165 153.145 55.160 153.135 55.160 ;
        RECT 153.145 55.160 154.905 55.165 ;
        RECT 150.830 55.130 151.390 55.160 ;
        POLYGON 150.770 55.130 150.770 55.055 150.685 55.055 ;
        RECT 150.770 55.110 151.390 55.130 ;
        POLYGON 151.390 55.160 151.465 55.160 151.390 55.110 ;
        POLYGON 153.135 55.160 153.135 55.155 153.125 55.155 ;
        RECT 153.135 55.155 154.905 55.160 ;
        POLYGON 153.125 55.155 153.125 55.140 153.090 55.140 ;
        RECT 153.125 55.145 154.905 55.155 ;
        POLYGON 154.905 55.175 154.935 55.145 154.905 55.145 ;
        POLYGON 157.045 55.175 157.060 55.175 157.060 55.170 ;
        RECT 157.060 55.170 157.865 55.175 ;
        POLYGON 157.060 55.170 157.090 55.170 157.090 55.155 ;
        RECT 157.090 55.155 157.865 55.170 ;
        POLYGON 157.090 55.155 157.105 55.155 157.105 55.145 ;
        RECT 157.105 55.145 157.865 55.155 ;
        RECT 153.125 55.140 154.935 55.145 ;
        POLYGON 153.090 55.140 153.090 55.110 153.030 55.110 ;
        RECT 153.090 55.120 154.935 55.140 ;
        POLYGON 154.935 55.145 154.965 55.120 154.935 55.120 ;
        POLYGON 157.110 55.145 157.160 55.145 157.160 55.120 ;
        RECT 157.160 55.135 157.865 55.145 ;
        POLYGON 157.865 55.180 157.945 55.135 157.865 55.135 ;
        POLYGON 158.790 55.180 158.850 55.180 158.850 55.135 ;
        RECT 158.850 55.150 159.580 55.180 ;
        POLYGON 159.580 55.255 159.705 55.150 159.580 55.150 ;
        POLYGON 160.380 55.255 160.400 55.255 160.400 55.240 ;
        RECT 160.400 55.240 161.305 55.255 ;
        POLYGON 160.400 55.240 160.490 55.240 160.490 55.150 ;
        RECT 160.490 55.180 161.305 55.240 ;
        POLYGON 161.305 55.300 161.415 55.180 161.305 55.180 ;
        POLYGON 162.545 55.300 162.585 55.300 162.585 55.245 ;
        RECT 162.585 55.290 163.830 55.300 ;
        POLYGON 163.830 55.415 163.915 55.290 163.830 55.290 ;
        POLYGON 165.510 55.415 165.575 55.415 165.575 55.295 ;
        RECT 165.575 55.290 167.635 55.415 ;
        RECT 162.585 55.245 163.915 55.290 ;
        POLYGON 162.585 55.245 162.630 55.245 162.630 55.185 ;
        RECT 162.630 55.180 163.915 55.245 ;
        RECT 160.490 55.150 161.415 55.180 ;
        RECT 158.850 55.135 159.705 55.150 ;
        POLYGON 159.705 55.150 159.720 55.135 159.705 55.135 ;
        POLYGON 160.490 55.150 160.505 55.150 160.505 55.135 ;
        RECT 160.505 55.135 161.415 55.150 ;
        RECT 157.160 55.120 157.945 55.135 ;
        POLYGON 157.945 55.135 157.965 55.120 157.945 55.120 ;
        POLYGON 158.850 55.135 158.870 55.135 158.870 55.120 ;
        RECT 158.870 55.120 159.720 55.135 ;
        RECT 153.090 55.110 154.965 55.120 ;
        POLYGON 154.965 55.120 154.970 55.110 154.965 55.110 ;
        POLYGON 157.160 55.120 157.180 55.120 157.180 55.110 ;
        RECT 157.180 55.110 157.965 55.120 ;
        RECT 150.770 55.055 151.315 55.110 ;
        RECT 148.990 55.030 149.850 55.055 ;
        POLYGON 148.935 55.030 148.935 55.020 148.930 55.020 ;
        RECT 148.935 55.025 149.850 55.030 ;
        POLYGON 149.850 55.055 149.875 55.055 149.850 55.025 ;
        POLYGON 150.685 55.055 150.685 55.025 150.655 55.025 ;
        RECT 150.685 55.050 151.315 55.055 ;
        POLYGON 151.315 55.110 151.390 55.110 151.315 55.050 ;
        POLYGON 153.030 55.110 153.030 55.080 152.965 55.080 ;
        RECT 153.030 55.085 154.970 55.110 ;
        POLYGON 154.970 55.110 155.010 55.085 154.970 55.085 ;
        POLYGON 157.180 55.110 157.195 55.110 157.195 55.105 ;
        RECT 157.195 55.105 157.965 55.110 ;
        POLYGON 157.195 55.105 157.235 55.105 157.235 55.085 ;
        RECT 157.235 55.085 157.965 55.105 ;
        RECT 153.030 55.080 155.010 55.085 ;
        POLYGON 152.960 55.080 152.960 55.065 152.930 55.065 ;
        RECT 152.960 55.075 155.010 55.080 ;
        POLYGON 155.010 55.085 155.020 55.075 155.010 55.075 ;
        POLYGON 157.235 55.085 157.255 55.085 157.255 55.075 ;
        RECT 157.255 55.075 157.965 55.085 ;
        RECT 152.960 55.065 155.020 55.075 ;
        POLYGON 152.930 55.065 152.930 55.060 152.925 55.060 ;
        RECT 152.930 55.060 155.020 55.065 ;
        POLYGON 152.925 55.060 152.925 55.050 152.905 55.050 ;
        RECT 152.925 55.050 155.020 55.060 ;
        POLYGON 155.020 55.075 155.070 55.050 155.020 55.050 ;
        POLYGON 157.255 55.075 157.305 55.075 157.305 55.050 ;
        RECT 157.305 55.050 157.965 55.075 ;
        RECT 150.685 55.025 151.245 55.050 ;
        RECT 148.935 55.020 149.795 55.025 ;
        POLYGON 148.930 55.020 148.930 54.910 148.850 54.910 ;
        RECT 148.930 54.965 149.795 55.020 ;
        POLYGON 149.795 55.025 149.850 55.025 149.795 54.965 ;
        POLYGON 150.655 55.025 150.655 55.000 150.625 55.000 ;
        RECT 150.655 55.000 151.245 55.025 ;
        POLYGON 151.245 55.050 151.310 55.050 151.245 55.000 ;
        POLYGON 152.905 55.050 152.905 55.000 152.815 55.000 ;
        RECT 152.905 55.020 155.070 55.050 ;
        POLYGON 155.070 55.050 155.125 55.020 155.070 55.020 ;
        POLYGON 157.305 55.050 157.365 55.050 157.365 55.020 ;
        RECT 157.365 55.035 157.965 55.050 ;
        POLYGON 157.965 55.120 158.105 55.035 157.965 55.035 ;
        POLYGON 158.870 55.120 158.885 55.120 158.885 55.110 ;
        RECT 158.885 55.110 159.720 55.120 ;
        POLYGON 158.885 55.110 158.915 55.110 158.915 55.085 ;
        RECT 158.915 55.090 159.720 55.110 ;
        POLYGON 159.720 55.135 159.775 55.090 159.720 55.090 ;
        POLYGON 160.505 55.135 160.550 55.135 160.550 55.090 ;
        RECT 160.550 55.090 161.415 55.135 ;
        RECT 158.915 55.085 159.775 55.090 ;
        POLYGON 158.915 55.085 158.950 55.085 158.950 55.055 ;
        RECT 158.950 55.065 159.775 55.085 ;
        POLYGON 159.775 55.090 159.800 55.065 159.775 55.065 ;
        POLYGON 160.550 55.090 160.575 55.090 160.575 55.065 ;
        RECT 160.575 55.065 161.415 55.090 ;
        RECT 158.950 55.055 159.800 55.065 ;
        POLYGON 158.950 55.055 158.970 55.055 158.970 55.035 ;
        RECT 158.970 55.035 159.800 55.055 ;
        RECT 157.365 55.020 158.105 55.035 ;
        POLYGON 158.105 55.035 158.130 55.020 158.105 55.020 ;
        POLYGON 158.970 55.035 158.990 55.035 158.990 55.020 ;
        RECT 158.990 55.020 159.800 55.035 ;
        RECT 152.905 55.015 155.125 55.020 ;
        POLYGON 155.125 55.020 155.130 55.015 155.125 55.015 ;
        POLYGON 157.370 55.020 157.380 55.020 157.380 55.015 ;
        RECT 157.380 55.015 158.130 55.020 ;
        RECT 152.905 55.000 155.130 55.015 ;
        POLYGON 150.625 55.000 150.625 54.965 150.590 54.965 ;
        RECT 150.625 54.965 151.160 55.000 ;
        RECT 148.930 54.910 149.710 54.965 ;
        RECT 117.275 54.800 147.830 54.910 ;
        POLYGON 147.830 54.910 147.900 54.910 147.830 54.800 ;
        POLYGON 148.850 54.910 148.850 54.800 148.775 54.800 ;
        RECT 148.850 54.870 149.710 54.910 ;
        POLYGON 149.710 54.965 149.795 54.965 149.710 54.870 ;
        POLYGON 150.590 54.965 150.590 54.925 150.545 54.925 ;
        RECT 150.590 54.935 151.160 54.965 ;
        POLYGON 151.160 55.000 151.245 55.000 151.160 54.935 ;
        POLYGON 152.815 55.000 152.815 54.955 152.730 54.955 ;
        RECT 152.815 54.985 155.130 55.000 ;
        POLYGON 155.130 55.015 155.195 54.985 155.130 54.985 ;
        POLYGON 157.380 55.015 157.385 55.015 157.385 55.010 ;
        RECT 157.385 55.010 158.130 55.015 ;
        POLYGON 157.390 55.010 157.430 55.010 157.430 54.985 ;
        RECT 157.430 54.985 158.130 55.010 ;
        POLYGON 158.130 55.020 158.185 54.985 158.130 54.985 ;
        POLYGON 158.990 55.020 159.035 55.020 159.035 54.985 ;
        RECT 159.035 54.985 159.800 55.020 ;
        RECT 152.815 54.980 155.200 54.985 ;
        POLYGON 155.200 54.985 155.205 54.980 155.200 54.980 ;
        POLYGON 157.430 54.985 157.440 54.985 157.440 54.980 ;
        RECT 157.440 54.980 158.190 54.985 ;
        RECT 152.815 54.955 155.205 54.980 ;
        POLYGON 155.205 54.980 155.270 54.955 155.205 54.955 ;
        POLYGON 157.440 54.980 157.485 54.980 157.485 54.955 ;
        RECT 157.485 54.955 158.190 54.980 ;
        POLYGON 158.190 54.985 158.230 54.955 158.190 54.955 ;
        POLYGON 159.035 54.985 159.060 54.985 159.060 54.965 ;
        RECT 159.060 54.965 159.800 54.985 ;
        POLYGON 159.060 54.965 159.070 54.965 159.070 54.955 ;
        RECT 159.070 54.955 159.800 54.965 ;
        POLYGON 152.725 54.955 152.725 54.950 152.715 54.950 ;
        RECT 152.725 54.950 155.275 54.955 ;
        POLYGON 157.485 54.955 157.495 54.955 157.495 54.950 ;
        RECT 157.495 54.950 158.230 54.955 ;
        POLYGON 152.715 54.950 152.715 54.935 152.695 54.935 ;
        RECT 152.715 54.935 155.280 54.950 ;
        RECT 150.590 54.925 151.075 54.935 ;
        POLYGON 150.545 54.925 150.545 54.870 150.490 54.870 ;
        RECT 150.545 54.870 151.075 54.925 ;
        RECT 148.850 54.800 149.610 54.870 ;
        RECT 117.275 54.720 147.780 54.800 ;
        POLYGON 147.780 54.800 147.830 54.800 147.780 54.720 ;
        POLYGON 148.775 54.800 148.775 54.780 148.760 54.780 ;
        RECT 148.775 54.780 149.610 54.800 ;
        POLYGON 148.760 54.780 148.760 54.755 148.740 54.755 ;
        RECT 148.760 54.755 149.610 54.780 ;
        POLYGON 149.610 54.870 149.710 54.870 149.610 54.755 ;
        POLYGON 150.490 54.870 150.490 54.810 150.425 54.810 ;
        RECT 150.490 54.860 151.075 54.870 ;
        POLYGON 151.075 54.935 151.160 54.935 151.075 54.860 ;
        POLYGON 152.690 54.935 152.690 54.925 152.680 54.925 ;
        RECT 152.690 54.925 155.280 54.935 ;
        POLYGON 152.680 54.925 152.680 54.860 152.560 54.860 ;
        RECT 152.680 54.920 155.280 54.925 ;
        POLYGON 155.280 54.950 155.370 54.920 155.280 54.920 ;
        POLYGON 157.495 54.950 157.545 54.950 157.545 54.925 ;
        RECT 157.545 54.945 158.230 54.950 ;
        POLYGON 158.230 54.955 158.245 54.945 158.230 54.945 ;
        POLYGON 159.070 54.955 159.080 54.955 159.080 54.945 ;
        RECT 159.080 54.945 159.800 54.955 ;
        RECT 157.545 54.925 158.245 54.945 ;
        POLYGON 157.545 54.925 157.550 54.925 157.550 54.920 ;
        RECT 157.550 54.920 158.245 54.925 ;
        RECT 152.680 54.915 155.370 54.920 ;
        POLYGON 155.370 54.920 155.380 54.915 155.370 54.915 ;
        POLYGON 157.550 54.920 157.560 54.920 157.560 54.915 ;
        RECT 157.560 54.915 158.245 54.920 ;
        RECT 152.680 54.890 155.390 54.915 ;
        POLYGON 155.390 54.915 155.445 54.890 155.390 54.890 ;
        POLYGON 157.560 54.915 157.600 54.915 157.600 54.890 ;
        RECT 157.600 54.890 158.245 54.915 ;
        RECT 152.680 54.885 155.460 54.890 ;
        POLYGON 155.460 54.890 155.465 54.885 155.460 54.885 ;
        POLYGON 157.600 54.890 157.610 54.890 157.610 54.885 ;
        RECT 157.610 54.885 158.245 54.890 ;
        RECT 152.680 54.860 155.465 54.885 ;
        RECT 150.490 54.810 150.945 54.860 ;
        POLYGON 150.425 54.810 150.425 54.755 150.370 54.755 ;
        RECT 150.425 54.755 150.945 54.810 ;
        POLYGON 148.740 54.755 148.740 54.720 148.715 54.720 ;
        RECT 148.740 54.720 149.565 54.755 ;
        RECT 117.275 54.680 147.760 54.720 ;
        POLYGON 147.760 54.720 147.780 54.720 147.760 54.680 ;
        POLYGON 148.715 54.720 148.715 54.685 148.690 54.685 ;
        RECT 148.715 54.695 149.565 54.720 ;
        POLYGON 149.565 54.755 149.610 54.755 149.565 54.695 ;
        POLYGON 150.370 54.755 150.370 54.695 150.310 54.695 ;
        RECT 150.370 54.750 150.945 54.755 ;
        POLYGON 150.945 54.860 151.075 54.860 150.945 54.750 ;
        POLYGON 152.560 54.860 152.560 54.845 152.535 54.845 ;
        RECT 152.560 54.855 155.465 54.860 ;
        POLYGON 155.465 54.885 155.570 54.855 155.465 54.855 ;
        POLYGON 157.610 54.885 157.660 54.885 157.660 54.855 ;
        RECT 157.660 54.855 158.245 54.885 ;
        RECT 152.560 54.845 155.570 54.855 ;
        POLYGON 152.535 54.845 152.535 54.825 152.505 54.825 ;
        RECT 152.535 54.840 155.570 54.845 ;
        POLYGON 155.570 54.855 155.630 54.840 155.570 54.840 ;
        POLYGON 157.665 54.855 157.685 54.855 157.685 54.845 ;
        RECT 157.685 54.850 158.245 54.855 ;
        POLYGON 158.245 54.945 158.380 54.850 158.245 54.850 ;
        POLYGON 159.080 54.945 159.125 54.945 159.125 54.910 ;
        RECT 159.125 54.935 159.800 54.945 ;
        POLYGON 159.800 55.065 159.935 54.935 159.800 54.935 ;
        POLYGON 160.575 55.065 160.640 55.065 160.640 55.000 ;
        RECT 160.640 55.020 161.415 55.065 ;
        POLYGON 161.415 55.180 161.555 55.020 161.415 55.020 ;
        POLYGON 162.630 55.180 162.735 55.180 162.735 55.045 ;
        RECT 162.735 55.150 163.915 55.180 ;
        POLYGON 163.915 55.290 164.010 55.150 163.915 55.150 ;
        POLYGON 165.575 55.290 165.650 55.290 165.650 55.150 ;
        RECT 165.650 55.150 167.635 55.290 ;
        RECT 162.735 55.060 164.010 55.150 ;
        POLYGON 164.010 55.150 164.065 55.060 164.010 55.060 ;
        POLYGON 165.650 55.150 165.675 55.150 165.675 55.105 ;
        RECT 165.675 55.105 167.635 55.150 ;
        POLYGON 165.675 55.105 165.695 55.105 165.695 55.060 ;
        RECT 165.695 55.060 167.635 55.105 ;
        RECT 162.735 55.045 164.065 55.060 ;
        POLYGON 162.735 55.045 162.750 55.045 162.750 55.020 ;
        RECT 162.750 55.020 164.065 55.045 ;
        RECT 160.640 55.000 161.555 55.020 ;
        POLYGON 160.640 55.000 160.695 55.000 160.695 54.935 ;
        RECT 160.695 54.940 161.555 55.000 ;
        POLYGON 161.555 55.020 161.620 54.940 161.555 54.940 ;
        POLYGON 162.750 55.020 162.785 55.020 162.785 54.970 ;
        RECT 162.785 55.000 164.065 55.020 ;
        POLYGON 164.065 55.060 164.105 55.000 164.065 55.000 ;
        POLYGON 165.695 55.060 165.725 55.060 165.725 55.000 ;
        RECT 165.725 55.000 167.635 55.060 ;
        RECT 162.785 54.970 164.105 55.000 ;
        POLYGON 162.785 54.970 162.805 54.970 162.805 54.940 ;
        RECT 162.805 54.940 164.105 54.970 ;
        RECT 160.695 54.935 161.620 54.940 ;
        RECT 159.125 54.910 159.940 54.935 ;
        POLYGON 159.125 54.910 159.130 54.910 159.130 54.905 ;
        RECT 159.130 54.905 159.940 54.910 ;
        POLYGON 159.130 54.905 159.180 54.905 159.180 54.865 ;
        RECT 159.180 54.870 159.940 54.905 ;
        POLYGON 159.940 54.935 160.005 54.870 159.940 54.870 ;
        POLYGON 160.695 54.935 160.760 54.935 160.760 54.870 ;
        RECT 160.760 54.910 161.620 54.935 ;
        POLYGON 161.620 54.940 161.645 54.910 161.620 54.910 ;
        POLYGON 162.805 54.940 162.825 54.940 162.825 54.910 ;
        RECT 162.825 54.920 164.105 54.940 ;
        POLYGON 164.105 55.000 164.155 54.920 164.105 54.920 ;
        POLYGON 165.725 55.000 165.765 55.000 165.765 54.920 ;
        RECT 165.765 54.995 167.635 55.000 ;
        POLYGON 167.635 55.430 167.840 54.995 167.635 54.995 ;
        POLYGON 170.445 55.430 170.455 55.430 170.455 55.410 ;
        RECT 170.455 55.410 174.425 55.430 ;
        POLYGON 170.455 55.410 170.490 55.410 170.490 55.325 ;
        RECT 170.490 55.325 174.425 55.410 ;
        POLYGON 170.490 55.325 170.495 55.325 170.495 55.310 ;
        RECT 170.495 55.310 174.425 55.325 ;
        POLYGON 170.495 55.310 170.610 55.310 170.610 55.005 ;
        RECT 170.610 55.275 174.425 55.310 ;
        POLYGON 174.425 56.295 174.845 55.275 174.425 55.275 ;
        POLYGON 181.490 56.295 181.610 56.295 181.610 55.955 ;
        RECT 181.610 55.955 195.530 56.295 ;
        POLYGON 181.610 55.955 181.675 55.955 181.675 55.765 ;
        RECT 181.675 55.845 195.530 55.955 ;
        POLYGON 195.530 57.125 195.955 55.845 195.530 55.845 ;
        RECT 206.225 57.050 222.255 57.130 ;
        POLYGON 206.225 57.050 206.245 57.050 206.245 56.410 ;
        RECT 206.245 56.410 222.255 57.050 ;
        POLYGON 206.245 56.410 206.265 56.410 206.265 55.870 ;
        RECT 206.265 55.845 222.255 56.410 ;
        RECT 181.675 55.765 195.955 55.845 ;
        POLYGON 181.675 55.765 181.815 55.765 181.815 55.275 ;
        RECT 181.815 55.645 195.955 55.765 ;
        POLYGON 195.955 55.845 196.020 55.645 195.955 55.645 ;
        POLYGON 206.265 55.845 206.270 55.845 206.270 55.735 ;
        RECT 206.270 55.655 222.255 55.845 ;
        POLYGON 222.255 57.505 222.360 57.505 222.255 55.655 ;
        POLYGON 229.935 57.515 229.935 57.425 229.910 57.425 ;
        RECT 229.935 57.425 234.430 57.520 ;
        POLYGON 234.430 57.755 234.570 57.755 234.430 57.425 ;
        POLYGON 237.850 57.755 237.850 57.625 237.775 57.625 ;
        RECT 237.850 57.660 240.230 57.755 ;
        POLYGON 240.230 57.795 240.330 57.795 240.230 57.660 ;
        POLYGON 242.370 57.795 242.370 57.765 242.340 57.765 ;
        RECT 242.370 57.765 244.105 57.795 ;
        POLYGON 242.340 57.765 242.340 57.660 242.240 57.660 ;
        RECT 242.340 57.680 244.105 57.765 ;
        POLYGON 244.105 57.810 244.260 57.810 244.105 57.680 ;
        POLYGON 245.980 57.810 245.980 57.790 245.945 57.790 ;
        RECT 245.980 57.800 247.950 57.810 ;
        POLYGON 247.950 57.830 248.050 57.830 247.950 57.800 ;
        POLYGON 252.305 57.830 252.345 57.830 252.345 57.820 ;
        RECT 252.345 57.820 254.550 57.830 ;
        POLYGON 252.345 57.820 252.410 57.820 252.410 57.805 ;
        RECT 252.410 57.805 254.550 57.820 ;
        RECT 252.415 57.800 254.550 57.805 ;
        RECT 245.980 57.790 247.895 57.800 ;
        POLYGON 245.945 57.790 245.945 57.745 245.875 57.745 ;
        RECT 245.945 57.785 247.895 57.790 ;
        POLYGON 247.895 57.800 247.950 57.800 247.895 57.785 ;
        POLYGON 252.415 57.800 252.470 57.800 252.470 57.785 ;
        RECT 252.470 57.785 254.550 57.800 ;
        RECT 245.945 57.750 247.785 57.785 ;
        POLYGON 247.785 57.785 247.895 57.785 247.785 57.750 ;
        POLYGON 252.470 57.785 252.510 57.785 252.510 57.775 ;
        RECT 252.510 57.775 254.550 57.785 ;
        POLYGON 252.510 57.775 252.525 57.775 252.525 57.770 ;
        RECT 252.525 57.770 254.550 57.775 ;
        POLYGON 252.525 57.770 252.595 57.770 252.595 57.750 ;
        RECT 252.595 57.750 254.550 57.770 ;
        RECT 245.945 57.745 247.610 57.750 ;
        POLYGON 245.875 57.745 245.875 57.710 245.815 57.710 ;
        RECT 245.875 57.710 247.610 57.745 ;
        POLYGON 245.815 57.710 245.815 57.680 245.765 57.680 ;
        RECT 245.815 57.695 247.610 57.710 ;
        POLYGON 247.610 57.750 247.785 57.750 247.610 57.695 ;
        POLYGON 252.595 57.750 252.690 57.750 252.690 57.725 ;
        RECT 252.690 57.725 254.550 57.750 ;
        POLYGON 252.690 57.725 252.760 57.725 252.760 57.700 ;
        RECT 252.760 57.720 254.550 57.725 ;
        POLYGON 254.550 57.840 254.755 57.720 254.550 57.720 ;
        POLYGON 256.550 57.840 256.560 57.840 256.560 57.835 ;
        RECT 256.560 57.835 258.545 57.840 ;
        POLYGON 256.560 57.835 256.570 57.835 256.570 57.825 ;
        RECT 256.570 57.825 258.545 57.835 ;
        POLYGON 256.570 57.825 256.695 57.825 256.695 57.720 ;
        RECT 256.695 57.730 258.545 57.825 ;
        POLYGON 258.545 57.955 258.775 57.730 258.545 57.730 ;
        POLYGON 261.020 57.955 261.085 57.955 261.085 57.875 ;
        RECT 261.085 57.875 264.140 57.955 ;
        POLYGON 261.085 57.875 261.165 57.875 261.165 57.780 ;
        RECT 261.165 57.780 264.140 57.875 ;
        POLYGON 261.165 57.780 261.175 57.780 261.175 57.770 ;
        RECT 261.175 57.770 264.140 57.780 ;
        POLYGON 261.175 57.770 261.205 57.770 261.205 57.730 ;
        RECT 261.205 57.730 264.140 57.770 ;
        RECT 256.695 57.720 258.775 57.730 ;
        RECT 252.760 57.700 254.760 57.720 ;
        POLYGON 252.760 57.700 252.775 57.700 252.775 57.695 ;
        RECT 252.775 57.695 254.760 57.700 ;
        RECT 245.815 57.680 247.515 57.695 ;
        RECT 242.340 57.675 244.100 57.680 ;
        POLYGON 244.100 57.680 244.105 57.680 244.100 57.675 ;
        POLYGON 245.765 57.680 245.765 57.675 245.760 57.675 ;
        RECT 245.765 57.675 247.515 57.680 ;
        RECT 242.340 57.660 244.020 57.675 ;
        RECT 237.850 57.650 240.225 57.660 ;
        POLYGON 240.225 57.660 240.230 57.660 240.225 57.650 ;
        POLYGON 242.240 57.660 242.240 57.650 242.230 57.650 ;
        RECT 242.240 57.650 244.020 57.660 ;
        RECT 237.850 57.625 240.210 57.650 ;
        POLYGON 240.210 57.650 240.225 57.650 240.210 57.625 ;
        POLYGON 242.230 57.650 242.230 57.625 242.210 57.625 ;
        RECT 242.230 57.625 244.020 57.650 ;
        POLYGON 237.775 57.625 237.775 57.550 237.730 57.550 ;
        RECT 237.775 57.550 240.095 57.625 ;
        POLYGON 237.730 57.550 237.730 57.520 237.715 57.520 ;
        RECT 237.730 57.520 240.095 57.550 ;
        POLYGON 237.715 57.520 237.715 57.435 237.670 57.435 ;
        RECT 237.715 57.460 240.095 57.520 ;
        POLYGON 240.095 57.625 240.210 57.625 240.095 57.460 ;
        POLYGON 242.210 57.625 242.210 57.575 242.160 57.575 ;
        RECT 242.210 57.605 244.020 57.625 ;
        POLYGON 244.020 57.675 244.100 57.675 244.020 57.605 ;
        POLYGON 245.760 57.675 245.760 57.615 245.660 57.615 ;
        RECT 245.760 57.665 247.515 57.675 ;
        POLYGON 247.515 57.695 247.610 57.695 247.515 57.665 ;
        POLYGON 252.775 57.695 252.805 57.695 252.805 57.685 ;
        RECT 252.805 57.685 254.760 57.695 ;
        POLYGON 252.810 57.685 252.860 57.685 252.860 57.665 ;
        RECT 252.860 57.665 254.760 57.685 ;
        RECT 245.760 57.660 247.510 57.665 ;
        POLYGON 247.510 57.665 247.515 57.665 247.510 57.660 ;
        POLYGON 252.860 57.665 252.875 57.665 252.875 57.660 ;
        RECT 252.875 57.660 254.760 57.665 ;
        RECT 245.760 57.630 247.425 57.660 ;
        POLYGON 247.425 57.660 247.510 57.660 247.425 57.630 ;
        POLYGON 252.875 57.660 252.890 57.660 252.890 57.655 ;
        RECT 252.890 57.655 254.760 57.660 ;
        POLYGON 254.760 57.720 254.860 57.655 254.760 57.655 ;
        POLYGON 256.695 57.720 256.755 57.720 256.755 57.675 ;
        RECT 256.755 57.715 258.775 57.720 ;
        POLYGON 258.775 57.730 258.790 57.715 258.775 57.715 ;
        POLYGON 261.205 57.730 261.215 57.730 261.215 57.715 ;
        RECT 261.215 57.715 264.140 57.730 ;
        RECT 256.755 57.675 258.790 57.715 ;
        POLYGON 256.755 57.675 256.775 57.675 256.775 57.655 ;
        RECT 256.775 57.670 258.790 57.675 ;
        POLYGON 258.790 57.715 258.830 57.670 258.790 57.670 ;
        POLYGON 261.215 57.715 261.250 57.715 261.250 57.670 ;
        RECT 261.250 57.670 264.140 57.715 ;
        RECT 256.775 57.655 258.830 57.670 ;
        POLYGON 252.895 57.655 252.965 57.655 252.965 57.630 ;
        RECT 252.965 57.630 254.865 57.655 ;
        RECT 245.760 57.615 247.330 57.630 ;
        POLYGON 245.660 57.615 245.660 57.605 245.645 57.605 ;
        RECT 245.660 57.605 247.330 57.615 ;
        RECT 242.210 57.575 243.955 57.605 ;
        POLYGON 242.160 57.575 242.160 57.515 242.105 57.515 ;
        RECT 242.160 57.545 243.955 57.575 ;
        POLYGON 243.955 57.605 244.020 57.605 243.955 57.545 ;
        POLYGON 245.645 57.605 245.645 57.560 245.580 57.560 ;
        RECT 245.645 57.595 247.330 57.605 ;
        POLYGON 247.330 57.630 247.425 57.630 247.330 57.595 ;
        POLYGON 252.965 57.630 253.010 57.630 253.010 57.615 ;
        RECT 253.010 57.615 254.865 57.630 ;
        POLYGON 253.010 57.615 253.030 57.615 253.030 57.605 ;
        RECT 253.030 57.605 254.865 57.615 ;
        POLYGON 253.030 57.605 253.055 57.605 253.055 57.595 ;
        RECT 253.055 57.595 254.865 57.605 ;
        RECT 245.645 57.565 247.250 57.595 ;
        POLYGON 247.250 57.595 247.330 57.595 247.250 57.565 ;
        POLYGON 253.055 57.595 253.085 57.595 253.085 57.585 ;
        RECT 253.085 57.585 254.865 57.595 ;
        POLYGON 253.085 57.585 253.135 57.585 253.135 57.565 ;
        RECT 253.135 57.565 254.865 57.585 ;
        RECT 245.645 57.560 247.195 57.565 ;
        POLYGON 245.580 57.560 245.580 57.545 245.555 57.545 ;
        RECT 245.580 57.545 247.195 57.560 ;
        POLYGON 247.195 57.565 247.250 57.565 247.195 57.545 ;
        POLYGON 253.135 57.565 253.185 57.565 253.185 57.545 ;
        RECT 253.185 57.545 254.865 57.565 ;
        RECT 242.160 57.515 243.870 57.545 ;
        POLYGON 242.105 57.510 242.105 57.460 242.060 57.460 ;
        RECT 242.105 57.465 243.870 57.515 ;
        POLYGON 243.870 57.545 243.955 57.545 243.870 57.465 ;
        POLYGON 245.555 57.545 245.555 57.515 245.510 57.515 ;
        RECT 245.555 57.515 247.075 57.545 ;
        POLYGON 245.510 57.515 245.510 57.465 245.440 57.465 ;
        RECT 245.510 57.495 247.075 57.515 ;
        POLYGON 247.075 57.545 247.195 57.545 247.075 57.495 ;
        POLYGON 253.185 57.545 253.260 57.545 253.260 57.515 ;
        RECT 253.260 57.515 254.865 57.545 ;
        POLYGON 253.260 57.515 253.305 57.515 253.305 57.495 ;
        RECT 253.305 57.495 254.865 57.515 ;
        RECT 245.510 57.465 246.985 57.495 ;
        RECT 242.105 57.460 243.775 57.465 ;
        RECT 237.715 57.435 239.995 57.460 ;
        POLYGON 237.670 57.435 237.670 57.425 237.665 57.425 ;
        RECT 237.670 57.425 239.995 57.435 ;
        POLYGON 229.910 57.425 229.910 57.365 229.895 57.365 ;
        RECT 229.910 57.365 234.390 57.425 ;
        POLYGON 229.895 57.365 229.895 56.780 229.745 56.780 ;
        RECT 229.895 57.330 234.390 57.365 ;
        POLYGON 234.390 57.425 234.430 57.425 234.390 57.330 ;
        POLYGON 237.665 57.425 237.665 57.330 237.615 57.330 ;
        RECT 237.665 57.330 239.995 57.425 ;
        RECT 229.895 57.300 234.380 57.330 ;
        POLYGON 234.380 57.330 234.390 57.330 234.380 57.300 ;
        POLYGON 237.615 57.330 237.615 57.300 237.600 57.300 ;
        RECT 237.615 57.315 239.995 57.330 ;
        POLYGON 239.995 57.460 240.095 57.460 239.995 57.315 ;
        POLYGON 242.060 57.460 242.060 57.315 241.935 57.315 ;
        RECT 242.060 57.380 243.775 57.460 ;
        POLYGON 243.775 57.465 243.870 57.465 243.775 57.380 ;
        POLYGON 245.440 57.465 245.440 57.425 245.380 57.425 ;
        RECT 245.440 57.450 246.985 57.465 ;
        POLYGON 246.985 57.495 247.075 57.495 246.985 57.450 ;
        POLYGON 253.305 57.495 253.355 57.495 253.355 57.475 ;
        RECT 253.355 57.485 254.865 57.495 ;
        POLYGON 254.865 57.655 255.135 57.485 254.865 57.485 ;
        POLYGON 256.775 57.655 256.890 57.655 256.890 57.560 ;
        RECT 256.890 57.590 258.830 57.655 ;
        POLYGON 258.830 57.670 258.905 57.590 258.830 57.590 ;
        POLYGON 261.250 57.670 261.300 57.670 261.300 57.600 ;
        RECT 261.300 57.605 264.140 57.670 ;
        POLYGON 264.140 57.955 264.355 57.605 264.140 57.605 ;
        POLYGON 268.605 57.955 268.705 57.955 268.705 57.775 ;
        RECT 268.705 57.775 275.775 57.955 ;
        POLYGON 268.705 57.775 268.730 57.775 268.730 57.735 ;
        RECT 268.730 57.735 275.775 57.775 ;
        POLYGON 268.730 57.735 268.795 57.735 268.795 57.610 ;
        RECT 268.795 57.605 275.775 57.735 ;
        RECT 261.300 57.600 264.355 57.605 ;
        POLYGON 261.300 57.600 261.305 57.600 261.305 57.590 ;
        RECT 261.305 57.590 264.355 57.600 ;
        RECT 256.890 57.560 258.905 57.590 ;
        POLYGON 256.890 57.560 256.930 57.560 256.930 57.530 ;
        RECT 256.930 57.530 258.905 57.560 ;
        POLYGON 256.930 57.530 256.975 57.530 256.975 57.485 ;
        RECT 256.975 57.485 258.905 57.530 ;
        RECT 253.355 57.475 255.135 57.485 ;
        POLYGON 253.360 57.475 253.410 57.475 253.410 57.450 ;
        RECT 253.410 57.465 255.135 57.475 ;
        POLYGON 255.135 57.485 255.165 57.465 255.135 57.465 ;
        POLYGON 256.975 57.485 256.985 57.485 256.985 57.480 ;
        RECT 256.985 57.480 258.905 57.485 ;
        POLYGON 256.985 57.480 257.000 57.480 257.000 57.465 ;
        RECT 257.000 57.465 258.905 57.480 ;
        RECT 253.410 57.450 255.165 57.465 ;
        RECT 245.440 57.445 246.970 57.450 ;
        POLYGON 246.970 57.450 246.980 57.450 246.970 57.445 ;
        POLYGON 253.410 57.450 253.420 57.450 253.420 57.445 ;
        RECT 253.420 57.445 255.165 57.450 ;
        RECT 245.440 57.425 246.790 57.445 ;
        POLYGON 245.380 57.425 245.380 57.380 245.320 57.380 ;
        RECT 245.380 57.380 246.790 57.425 ;
        RECT 242.060 57.315 243.660 57.380 ;
        RECT 237.615 57.305 239.990 57.315 ;
        POLYGON 239.990 57.315 239.995 57.315 239.990 57.305 ;
        POLYGON 241.935 57.315 241.935 57.310 241.930 57.310 ;
        RECT 241.935 57.310 243.660 57.315 ;
        RECT 237.615 57.300 239.905 57.305 ;
        RECT 229.895 56.780 234.095 57.300 ;
        POLYGON 229.745 56.780 229.745 55.655 229.525 55.655 ;
        RECT 229.745 56.520 234.095 56.780 ;
        POLYGON 234.095 57.300 234.380 57.300 234.095 56.520 ;
        POLYGON 237.600 57.300 237.600 56.785 237.335 56.785 ;
        RECT 237.600 57.170 239.905 57.300 ;
        POLYGON 239.905 57.305 239.990 57.305 239.905 57.170 ;
        POLYGON 241.930 57.305 241.930 57.250 241.880 57.250 ;
        RECT 241.930 57.270 243.660 57.310 ;
        POLYGON 243.660 57.380 243.775 57.380 243.660 57.270 ;
        POLYGON 245.320 57.380 245.320 57.340 245.265 57.340 ;
        RECT 245.320 57.365 246.790 57.380 ;
        POLYGON 246.790 57.445 246.970 57.445 246.790 57.365 ;
        POLYGON 253.420 57.445 253.460 57.445 253.460 57.425 ;
        RECT 253.460 57.425 255.165 57.445 ;
        POLYGON 250.405 57.425 250.405 57.420 250.220 57.420 ;
        RECT 250.405 57.420 250.465 57.425 ;
        POLYGON 250.180 57.420 250.180 57.415 250.060 57.415 ;
        RECT 250.180 57.415 250.465 57.420 ;
        POLYGON 250.465 57.425 250.680 57.415 250.465 57.415 ;
        POLYGON 253.460 57.425 253.480 57.425 253.480 57.415 ;
        RECT 253.480 57.415 255.165 57.425 ;
        POLYGON 250.050 57.415 250.050 57.410 249.915 57.410 ;
        RECT 250.050 57.410 250.705 57.415 ;
        POLYGON 249.890 57.410 249.890 57.400 249.760 57.400 ;
        RECT 249.890 57.400 250.705 57.410 ;
        POLYGON 250.705 57.415 250.855 57.400 250.705 57.400 ;
        POLYGON 253.480 57.415 253.505 57.415 253.505 57.405 ;
        RECT 253.505 57.405 255.165 57.415 ;
        POLYGON 253.505 57.405 253.515 57.405 253.515 57.400 ;
        RECT 253.515 57.400 255.165 57.405 ;
        POLYGON 249.755 57.400 249.755 57.395 249.730 57.395 ;
        RECT 249.755 57.395 250.865 57.400 ;
        POLYGON 250.865 57.400 250.905 57.395 250.865 57.395 ;
        POLYGON 253.515 57.400 253.530 57.400 253.530 57.395 ;
        RECT 253.530 57.395 255.165 57.400 ;
        POLYGON 249.725 57.395 249.725 57.390 249.650 57.390 ;
        RECT 249.725 57.390 250.915 57.395 ;
        POLYGON 250.915 57.395 250.965 57.390 250.915 57.390 ;
        POLYGON 253.530 57.395 253.540 57.395 253.540 57.390 ;
        RECT 253.540 57.390 255.165 57.395 ;
        POLYGON 249.640 57.390 249.640 57.365 249.450 57.365 ;
        RECT 249.640 57.370 250.965 57.390 ;
        POLYGON 250.965 57.390 251.135 57.370 250.965 57.370 ;
        POLYGON 253.540 57.390 253.580 57.390 253.580 57.375 ;
        RECT 253.580 57.375 255.165 57.390 ;
        POLYGON 253.580 57.375 253.590 57.375 253.590 57.370 ;
        RECT 253.590 57.370 255.165 57.375 ;
        RECT 249.640 57.365 251.145 57.370 ;
        RECT 245.320 57.340 246.740 57.365 ;
        POLYGON 246.740 57.365 246.790 57.365 246.740 57.340 ;
        POLYGON 249.450 57.365 249.450 57.360 249.410 57.360 ;
        RECT 249.450 57.360 251.145 57.365 ;
        POLYGON 251.145 57.370 251.225 57.360 251.145 57.360 ;
        POLYGON 253.590 57.370 253.610 57.370 253.610 57.360 ;
        RECT 253.610 57.360 255.165 57.370 ;
        POLYGON 249.405 57.360 249.405 57.355 249.385 57.355 ;
        RECT 249.405 57.355 251.250 57.360 ;
        POLYGON 249.375 57.355 249.375 57.345 249.300 57.345 ;
        RECT 249.375 57.345 251.250 57.355 ;
        POLYGON 249.300 57.345 249.300 57.340 249.270 57.340 ;
        RECT 249.300 57.340 251.250 57.345 ;
        POLYGON 245.265 57.340 245.265 57.335 245.260 57.335 ;
        RECT 245.265 57.335 246.655 57.340 ;
        POLYGON 245.260 57.335 245.260 57.270 245.170 57.270 ;
        RECT 245.260 57.295 246.655 57.335 ;
        POLYGON 246.655 57.340 246.740 57.340 246.655 57.295 ;
        POLYGON 249.270 57.340 249.270 57.315 249.120 57.315 ;
        RECT 249.270 57.330 251.250 57.340 ;
        POLYGON 251.250 57.360 251.425 57.330 251.250 57.330 ;
        POLYGON 253.610 57.360 253.670 57.360 253.670 57.330 ;
        RECT 253.670 57.330 255.165 57.360 ;
        RECT 249.270 57.320 251.425 57.330 ;
        POLYGON 251.425 57.330 251.485 57.320 251.425 57.320 ;
        POLYGON 253.670 57.330 253.685 57.330 253.685 57.325 ;
        RECT 253.685 57.325 255.165 57.330 ;
        POLYGON 253.685 57.325 253.690 57.325 253.690 57.320 ;
        RECT 253.690 57.320 255.165 57.325 ;
        RECT 249.270 57.315 251.485 57.320 ;
        POLYGON 249.120 57.315 249.120 57.295 249.020 57.295 ;
        RECT 249.120 57.295 251.485 57.315 ;
        POLYGON 251.485 57.320 251.605 57.295 251.485 57.295 ;
        POLYGON 253.690 57.320 253.740 57.320 253.740 57.295 ;
        RECT 253.740 57.295 255.165 57.320 ;
        RECT 245.260 57.270 246.540 57.295 ;
        RECT 241.930 57.250 243.630 57.270 ;
        POLYGON 241.880 57.250 241.880 57.170 241.815 57.170 ;
        RECT 241.880 57.240 243.630 57.250 ;
        POLYGON 243.630 57.270 243.660 57.270 243.630 57.240 ;
        POLYGON 245.170 57.270 245.170 57.240 245.130 57.240 ;
        RECT 245.170 57.240 246.540 57.270 ;
        POLYGON 246.540 57.295 246.655 57.295 246.540 57.240 ;
        POLYGON 249.020 57.295 249.020 57.265 248.875 57.265 ;
        RECT 249.020 57.270 251.625 57.295 ;
        POLYGON 251.625 57.295 251.745 57.270 251.625 57.270 ;
        POLYGON 253.740 57.295 253.790 57.295 253.790 57.270 ;
        RECT 253.790 57.290 255.165 57.295 ;
        POLYGON 255.165 57.465 255.420 57.290 255.165 57.290 ;
        POLYGON 257.000 57.465 257.190 57.465 257.190 57.290 ;
        RECT 257.190 57.380 258.905 57.465 ;
        POLYGON 258.905 57.590 259.105 57.380 258.905 57.380 ;
        POLYGON 261.305 57.590 261.425 57.590 261.425 57.435 ;
        RECT 261.425 57.500 264.355 57.590 ;
        POLYGON 264.355 57.605 264.420 57.500 264.355 57.500 ;
        POLYGON 268.795 57.605 268.845 57.605 268.845 57.520 ;
        RECT 268.845 57.520 275.775 57.605 ;
        POLYGON 268.845 57.520 268.850 57.520 268.850 57.505 ;
        RECT 268.850 57.500 275.775 57.520 ;
        RECT 261.425 57.445 264.420 57.500 ;
        POLYGON 264.420 57.500 264.455 57.445 264.420 57.445 ;
        POLYGON 268.850 57.500 268.880 57.500 268.880 57.445 ;
        RECT 268.880 57.445 275.775 57.500 ;
        RECT 261.425 57.435 264.455 57.445 ;
        POLYGON 261.425 57.435 261.460 57.435 261.460 57.385 ;
        RECT 261.460 57.380 264.455 57.435 ;
        RECT 257.190 57.355 259.105 57.380 ;
        POLYGON 259.105 57.380 259.130 57.355 259.105 57.355 ;
        POLYGON 261.460 57.380 261.480 57.380 261.480 57.355 ;
        RECT 261.480 57.355 264.455 57.380 ;
        RECT 257.190 57.330 259.130 57.355 ;
        POLYGON 259.130 57.355 259.150 57.330 259.130 57.330 ;
        POLYGON 261.480 57.355 261.495 57.355 261.495 57.340 ;
        RECT 261.495 57.340 264.455 57.355 ;
        POLYGON 261.495 57.340 261.500 57.340 261.500 57.330 ;
        RECT 261.500 57.330 264.455 57.340 ;
        RECT 257.190 57.290 259.150 57.330 ;
        RECT 253.790 57.270 255.420 57.290 ;
        RECT 249.020 57.265 251.745 57.270 ;
        POLYGON 248.875 57.265 248.875 57.260 248.850 57.260 ;
        RECT 248.875 57.260 251.745 57.265 ;
        POLYGON 248.840 57.260 248.840 57.245 248.785 57.245 ;
        RECT 248.840 57.245 251.745 57.260 ;
        POLYGON 248.785 57.245 248.785 57.240 248.765 57.240 ;
        RECT 248.785 57.240 251.745 57.245 ;
        RECT 241.880 57.170 243.455 57.240 ;
        RECT 237.600 57.045 239.830 57.170 ;
        POLYGON 239.830 57.170 239.905 57.170 239.830 57.045 ;
        POLYGON 241.815 57.170 241.815 57.045 241.715 57.045 ;
        RECT 241.815 57.070 243.455 57.170 ;
        POLYGON 243.455 57.240 243.630 57.240 243.455 57.070 ;
        POLYGON 245.130 57.240 245.130 57.225 245.110 57.225 ;
        RECT 245.130 57.235 246.530 57.240 ;
        POLYGON 246.530 57.240 246.540 57.240 246.530 57.235 ;
        POLYGON 248.765 57.240 248.765 57.235 248.745 57.235 ;
        RECT 248.765 57.235 251.745 57.240 ;
        RECT 245.130 57.225 246.505 57.235 ;
        POLYGON 245.110 57.225 245.110 57.070 244.915 57.070 ;
        RECT 245.110 57.220 246.505 57.225 ;
        POLYGON 246.505 57.235 246.530 57.235 246.505 57.220 ;
        POLYGON 248.745 57.235 248.745 57.220 248.685 57.220 ;
        RECT 248.745 57.225 251.745 57.235 ;
        POLYGON 251.745 57.270 251.925 57.225 251.745 57.225 ;
        POLYGON 253.790 57.270 253.800 57.270 253.800 57.265 ;
        RECT 253.800 57.265 255.420 57.270 ;
        POLYGON 255.420 57.290 255.455 57.265 255.420 57.265 ;
        POLYGON 257.190 57.290 257.200 57.290 257.200 57.285 ;
        RECT 257.200 57.285 259.150 57.290 ;
        POLYGON 257.200 57.285 257.215 57.285 257.215 57.275 ;
        RECT 257.215 57.275 259.150 57.285 ;
        POLYGON 257.215 57.275 257.225 57.275 257.225 57.265 ;
        RECT 257.225 57.265 259.150 57.275 ;
        POLYGON 253.800 57.265 253.870 57.265 253.870 57.225 ;
        RECT 253.870 57.230 255.460 57.265 ;
        POLYGON 255.460 57.265 255.500 57.230 255.460 57.230 ;
        POLYGON 257.225 57.265 257.260 57.265 257.260 57.230 ;
        RECT 257.260 57.230 259.150 57.265 ;
        RECT 253.870 57.225 255.505 57.230 ;
        RECT 248.745 57.220 251.925 57.225 ;
        RECT 245.110 57.095 246.275 57.220 ;
        POLYGON 246.275 57.220 246.505 57.220 246.275 57.095 ;
        POLYGON 248.685 57.220 248.685 57.170 248.485 57.170 ;
        RECT 248.685 57.210 251.925 57.220 ;
        POLYGON 251.925 57.225 251.990 57.210 251.925 57.210 ;
        POLYGON 253.870 57.225 253.900 57.225 253.900 57.210 ;
        RECT 253.900 57.210 255.505 57.225 ;
        RECT 248.685 57.205 251.990 57.210 ;
        POLYGON 251.990 57.210 252.000 57.205 251.990 57.205 ;
        POLYGON 253.900 57.210 253.910 57.210 253.910 57.205 ;
        RECT 253.910 57.205 255.505 57.210 ;
        RECT 248.685 57.190 252.000 57.205 ;
        POLYGON 252.000 57.205 252.065 57.190 252.000 57.190 ;
        POLYGON 253.910 57.205 253.940 57.205 253.940 57.190 ;
        RECT 253.940 57.190 255.505 57.205 ;
        RECT 248.685 57.170 252.065 57.190 ;
        POLYGON 248.480 57.170 248.480 57.145 248.395 57.145 ;
        RECT 248.480 57.145 252.065 57.170 ;
        POLYGON 248.390 57.145 248.390 57.140 248.380 57.140 ;
        RECT 248.390 57.140 252.065 57.145 ;
        POLYGON 248.380 57.140 248.380 57.120 248.320 57.120 ;
        RECT 248.380 57.135 252.065 57.140 ;
        POLYGON 252.065 57.190 252.255 57.135 252.065 57.135 ;
        POLYGON 253.940 57.190 253.995 57.190 253.995 57.165 ;
        RECT 253.995 57.165 255.505 57.190 ;
        POLYGON 253.995 57.165 254.005 57.165 254.005 57.160 ;
        RECT 254.005 57.160 255.505 57.165 ;
        POLYGON 254.005 57.160 254.010 57.160 254.010 57.155 ;
        RECT 254.010 57.155 255.505 57.160 ;
        POLYGON 254.015 57.155 254.045 57.155 254.045 57.135 ;
        RECT 254.045 57.135 255.505 57.155 ;
        RECT 248.380 57.120 252.255 57.135 ;
        POLYGON 248.320 57.120 248.320 57.095 248.235 57.095 ;
        RECT 248.320 57.105 252.255 57.120 ;
        POLYGON 252.255 57.135 252.345 57.105 252.255 57.105 ;
        POLYGON 254.045 57.135 254.095 57.135 254.095 57.105 ;
        RECT 254.095 57.105 255.505 57.135 ;
        RECT 248.320 57.095 252.345 57.105 ;
        RECT 245.110 57.070 246.240 57.095 ;
        POLYGON 246.240 57.095 246.275 57.095 246.240 57.075 ;
        POLYGON 248.235 57.095 248.235 57.080 248.185 57.080 ;
        RECT 248.235 57.080 252.345 57.095 ;
        POLYGON 252.345 57.105 252.415 57.080 252.345 57.080 ;
        POLYGON 254.095 57.105 254.130 57.105 254.130 57.085 ;
        RECT 254.130 57.085 255.505 57.105 ;
        POLYGON 254.130 57.085 254.135 57.085 254.135 57.080 ;
        RECT 254.135 57.080 255.505 57.085 ;
        POLYGON 248.185 57.080 248.185 57.075 248.170 57.075 ;
        RECT 248.185 57.075 252.415 57.080 ;
        POLYGON 248.170 57.075 248.170 57.070 248.155 57.070 ;
        RECT 248.170 57.070 252.415 57.075 ;
        RECT 241.815 57.045 243.375 57.070 ;
        RECT 237.600 56.935 239.760 57.045 ;
        POLYGON 239.760 57.045 239.830 57.045 239.760 56.940 ;
        POLYGON 241.715 57.045 241.715 57.040 241.710 57.040 ;
        RECT 241.715 57.040 243.375 57.045 ;
        POLYGON 241.710 57.040 241.710 56.985 241.670 56.985 ;
        RECT 241.710 56.990 243.375 57.040 ;
        POLYGON 243.375 57.070 243.455 57.070 243.375 56.990 ;
        POLYGON 244.915 57.070 244.915 57.060 244.900 57.060 ;
        RECT 244.915 57.060 246.055 57.070 ;
        POLYGON 244.900 57.060 244.900 57.015 244.845 57.015 ;
        RECT 244.900 57.015 246.055 57.060 ;
        POLYGON 244.845 57.015 244.845 56.990 244.820 56.990 ;
        RECT 244.845 56.990 246.055 57.015 ;
        RECT 241.710 56.985 243.245 56.990 ;
        POLYGON 241.670 56.985 241.670 56.940 241.635 56.940 ;
        RECT 241.670 56.940 243.245 56.985 ;
        RECT 237.600 56.815 239.690 56.935 ;
        POLYGON 239.690 56.935 239.760 56.935 239.690 56.815 ;
        POLYGON 241.635 56.940 241.635 56.870 241.585 56.870 ;
        RECT 241.635 56.870 243.245 56.940 ;
        POLYGON 241.585 56.870 241.585 56.815 241.545 56.815 ;
        RECT 241.585 56.855 243.245 56.870 ;
        POLYGON 243.245 56.990 243.375 56.990 243.245 56.855 ;
        POLYGON 244.820 56.990 244.820 56.970 244.795 56.970 ;
        RECT 244.820 56.970 246.055 56.990 ;
        POLYGON 244.795 56.970 244.795 56.855 244.665 56.855 ;
        RECT 244.795 56.960 246.055 56.970 ;
        POLYGON 246.055 57.070 246.235 57.070 246.055 56.960 ;
        POLYGON 248.155 57.070 248.155 57.035 248.050 57.035 ;
        RECT 248.155 57.050 252.415 57.070 ;
        POLYGON 252.415 57.080 252.510 57.050 252.415 57.050 ;
        POLYGON 254.135 57.080 254.185 57.080 254.185 57.050 ;
        RECT 254.185 57.060 255.505 57.080 ;
        POLYGON 255.505 57.230 255.735 57.060 255.505 57.060 ;
        POLYGON 257.260 57.230 257.275 57.230 257.275 57.215 ;
        RECT 257.275 57.215 259.150 57.230 ;
        POLYGON 257.275 57.215 257.410 57.215 257.410 57.090 ;
        RECT 257.410 57.090 259.150 57.215 ;
        POLYGON 257.410 57.090 257.440 57.090 257.440 57.060 ;
        RECT 257.440 57.080 259.150 57.090 ;
        POLYGON 259.150 57.330 259.370 57.080 259.150 57.080 ;
        POLYGON 261.500 57.330 261.535 57.330 261.535 57.280 ;
        RECT 261.535 57.280 264.455 57.330 ;
        POLYGON 261.535 57.280 261.580 57.280 261.580 57.210 ;
        RECT 261.580 57.210 264.455 57.280 ;
        POLYGON 261.580 57.210 261.635 57.210 261.635 57.135 ;
        RECT 261.635 57.135 264.455 57.210 ;
        POLYGON 261.635 57.135 261.665 57.135 261.665 57.090 ;
        RECT 261.665 57.090 264.455 57.135 ;
        POLYGON 261.665 57.090 261.670 57.090 261.670 57.080 ;
        RECT 261.670 57.080 264.455 57.090 ;
        RECT 257.440 57.060 259.370 57.080 ;
        RECT 254.185 57.055 255.735 57.060 ;
        POLYGON 255.735 57.060 255.740 57.055 255.735 57.055 ;
        POLYGON 257.440 57.060 257.445 57.060 257.445 57.055 ;
        RECT 257.445 57.055 259.370 57.060 ;
        RECT 254.185 57.050 255.740 57.055 ;
        RECT 248.155 57.045 252.510 57.050 ;
        POLYGON 252.510 57.050 252.525 57.045 252.510 57.045 ;
        POLYGON 254.185 57.050 254.195 57.050 254.195 57.045 ;
        RECT 254.195 57.045 255.740 57.050 ;
        RECT 248.155 57.035 252.525 57.045 ;
        POLYGON 248.050 57.035 248.050 57.000 247.950 57.000 ;
        RECT 248.050 57.000 252.525 57.035 ;
        POLYGON 247.945 57.000 247.945 56.980 247.895 56.980 ;
        RECT 247.945 56.985 252.525 57.000 ;
        POLYGON 252.525 57.045 252.690 56.985 252.525 56.985 ;
        POLYGON 254.195 57.045 254.220 57.045 254.220 57.030 ;
        RECT 254.220 57.030 255.740 57.045 ;
        POLYGON 254.220 57.030 254.235 57.030 254.235 57.025 ;
        RECT 254.235 57.025 255.740 57.030 ;
        POLYGON 254.235 57.025 254.295 57.025 254.295 56.985 ;
        RECT 254.295 56.995 255.740 57.025 ;
        POLYGON 255.740 57.055 255.815 56.995 255.740 56.995 ;
        POLYGON 257.445 57.055 257.505 57.055 257.505 56.995 ;
        RECT 257.505 56.995 259.370 57.055 ;
        RECT 254.295 56.985 255.815 56.995 ;
        RECT 247.945 56.980 252.690 56.985 ;
        POLYGON 247.890 56.980 247.890 56.960 247.840 56.960 ;
        RECT 247.890 56.960 252.690 56.980 ;
        RECT 244.795 56.945 246.030 56.960 ;
        POLYGON 246.030 56.960 246.055 56.960 246.030 56.945 ;
        POLYGON 247.840 56.960 247.840 56.945 247.800 56.945 ;
        RECT 247.840 56.955 252.690 56.960 ;
        POLYGON 252.690 56.985 252.760 56.955 252.690 56.955 ;
        POLYGON 254.295 56.985 254.315 56.985 254.315 56.975 ;
        RECT 254.315 56.975 255.815 56.985 ;
        POLYGON 254.315 56.975 254.345 56.975 254.345 56.955 ;
        RECT 254.345 56.960 255.815 56.975 ;
        POLYGON 255.815 56.995 255.860 56.960 255.815 56.960 ;
        POLYGON 257.505 56.995 257.530 56.995 257.530 56.975 ;
        RECT 257.530 56.975 259.370 56.995 ;
        POLYGON 257.530 56.975 257.540 56.975 257.540 56.960 ;
        RECT 257.540 56.960 259.370 56.975 ;
        RECT 254.345 56.955 255.865 56.960 ;
        RECT 247.840 56.945 252.760 56.955 ;
        RECT 244.795 56.890 245.945 56.945 ;
        POLYGON 245.945 56.945 246.030 56.945 245.945 56.890 ;
        POLYGON 247.800 56.945 247.800 56.940 247.785 56.940 ;
        RECT 247.800 56.940 252.760 56.945 ;
        POLYGON 247.785 56.940 247.785 56.890 247.660 56.890 ;
        RECT 247.785 56.935 252.760 56.940 ;
        POLYGON 252.760 56.955 252.810 56.935 252.760 56.935 ;
        POLYGON 254.345 56.955 254.380 56.955 254.380 56.935 ;
        RECT 254.380 56.935 255.865 56.955 ;
        RECT 247.785 56.900 252.810 56.935 ;
        POLYGON 252.810 56.935 252.890 56.900 252.810 56.900 ;
        POLYGON 254.380 56.935 254.430 56.935 254.430 56.900 ;
        RECT 254.430 56.900 255.865 56.935 ;
        RECT 247.785 56.890 252.895 56.900 ;
        RECT 244.795 56.855 245.845 56.890 ;
        RECT 241.585 56.840 243.235 56.855 ;
        POLYGON 243.235 56.855 243.245 56.855 243.235 56.840 ;
        POLYGON 244.665 56.855 244.665 56.840 244.645 56.840 ;
        RECT 244.665 56.840 245.845 56.855 ;
        RECT 241.585 56.815 243.145 56.840 ;
        RECT 237.600 56.785 239.655 56.815 ;
        POLYGON 237.335 56.785 237.335 56.520 237.220 56.520 ;
        RECT 237.335 56.760 239.655 56.785 ;
        POLYGON 239.655 56.815 239.690 56.815 239.655 56.760 ;
        POLYGON 241.545 56.815 241.545 56.760 241.505 56.760 ;
        RECT 241.545 56.760 243.145 56.815 ;
        RECT 237.335 56.750 239.650 56.760 ;
        POLYGON 239.650 56.760 239.655 56.760 239.650 56.750 ;
        POLYGON 241.505 56.760 241.505 56.755 241.500 56.755 ;
        RECT 241.505 56.755 243.145 56.760 ;
        RECT 237.335 56.585 239.560 56.750 ;
        POLYGON 239.560 56.750 239.650 56.750 239.560 56.585 ;
        POLYGON 241.500 56.750 241.500 56.725 241.480 56.725 ;
        RECT 241.500 56.745 243.145 56.755 ;
        POLYGON 243.145 56.840 243.235 56.840 243.145 56.745 ;
        POLYGON 244.645 56.840 244.645 56.790 244.590 56.790 ;
        RECT 244.645 56.820 245.845 56.840 ;
        POLYGON 245.845 56.890 245.945 56.890 245.845 56.820 ;
        POLYGON 247.660 56.890 247.660 56.870 247.610 56.870 ;
        RECT 247.660 56.870 252.895 56.890 ;
        POLYGON 247.610 56.870 247.610 56.835 247.515 56.835 ;
        RECT 247.610 56.850 252.895 56.870 ;
        POLYGON 252.895 56.900 253.010 56.850 252.895 56.850 ;
        POLYGON 254.430 56.900 254.470 56.900 254.470 56.875 ;
        RECT 254.470 56.875 255.865 56.900 ;
        POLYGON 254.475 56.875 254.510 56.875 254.510 56.850 ;
        RECT 254.510 56.850 255.865 56.875 ;
        RECT 247.610 56.845 253.010 56.850 ;
        POLYGON 253.010 56.850 253.030 56.845 253.010 56.845 ;
        POLYGON 254.510 56.850 254.515 56.850 254.515 56.845 ;
        RECT 254.515 56.845 255.865 56.850 ;
        POLYGON 255.865 56.960 256.005 56.845 255.865 56.845 ;
        POLYGON 257.540 56.960 257.625 56.960 257.625 56.875 ;
        RECT 257.625 56.945 259.370 56.960 ;
        POLYGON 259.370 57.080 259.475 56.945 259.370 56.945 ;
        POLYGON 261.670 57.080 261.720 57.080 261.720 57.010 ;
        RECT 261.720 57.035 264.455 57.080 ;
        POLYGON 264.455 57.445 264.690 57.035 264.455 57.035 ;
        POLYGON 268.880 57.445 269.070 57.445 269.070 57.040 ;
        RECT 269.070 57.335 275.775 57.445 ;
        POLYGON 275.775 58.100 276.090 57.335 275.775 57.335 ;
        RECT 269.070 57.275 276.090 57.335 ;
        POLYGON 276.090 57.335 276.115 57.275 276.090 57.275 ;
        RECT 269.070 57.035 276.115 57.275 ;
        RECT 261.720 57.010 264.690 57.035 ;
        POLYGON 261.720 57.010 261.735 57.010 261.735 56.990 ;
        RECT 261.735 56.990 264.690 57.010 ;
        POLYGON 261.735 56.990 261.760 56.990 261.760 56.950 ;
        RECT 261.760 56.980 264.690 56.990 ;
        POLYGON 264.690 57.035 264.720 56.980 264.690 56.980 ;
        POLYGON 269.070 57.035 269.100 57.035 269.100 56.980 ;
        RECT 269.100 56.980 276.115 57.035 ;
        RECT 261.760 56.945 264.720 56.980 ;
        RECT 257.625 56.925 259.475 56.945 ;
        POLYGON 259.475 56.945 259.495 56.925 259.475 56.925 ;
        POLYGON 261.760 56.945 261.775 56.945 261.775 56.925 ;
        RECT 261.775 56.925 264.720 56.945 ;
        RECT 257.625 56.875 259.495 56.925 ;
        POLYGON 257.625 56.875 257.650 56.875 257.650 56.845 ;
        RECT 257.650 56.845 259.495 56.875 ;
        RECT 247.610 56.835 253.030 56.845 ;
        POLYGON 247.515 56.835 247.515 56.830 247.510 56.830 ;
        RECT 247.515 56.830 253.030 56.835 ;
        POLYGON 247.510 56.830 247.510 56.820 247.485 56.820 ;
        RECT 247.510 56.820 253.030 56.830 ;
        POLYGON 253.030 56.845 253.085 56.820 253.030 56.820 ;
        POLYGON 254.515 56.845 254.545 56.845 254.545 56.825 ;
        RECT 254.545 56.840 256.005 56.845 ;
        POLYGON 256.005 56.845 256.015 56.840 256.005 56.840 ;
        POLYGON 257.650 56.845 257.655 56.845 257.655 56.840 ;
        RECT 257.655 56.840 259.495 56.845 ;
        RECT 254.545 56.825 256.015 56.840 ;
        POLYGON 254.545 56.825 254.550 56.825 254.550 56.820 ;
        RECT 254.550 56.820 256.015 56.825 ;
        RECT 244.645 56.790 245.790 56.820 ;
        POLYGON 245.790 56.820 245.840 56.820 245.790 56.790 ;
        POLYGON 247.485 56.820 247.485 56.795 247.425 56.795 ;
        RECT 247.485 56.800 253.085 56.820 ;
        RECT 247.485 56.795 250.290 56.800 ;
        POLYGON 250.290 56.800 250.315 56.800 250.290 56.795 ;
        POLYGON 250.315 56.800 250.370 56.800 250.370 56.795 ;
        RECT 250.370 56.795 253.085 56.800 ;
        POLYGON 247.425 56.795 247.425 56.790 247.415 56.790 ;
        RECT 247.425 56.790 250.055 56.795 ;
        POLYGON 250.055 56.795 250.180 56.795 250.055 56.790 ;
        POLYGON 250.595 56.795 250.640 56.795 250.640 56.790 ;
        RECT 250.640 56.790 253.085 56.795 ;
        POLYGON 244.590 56.790 244.590 56.745 244.540 56.745 ;
        RECT 244.590 56.745 245.660 56.790 ;
        RECT 241.500 56.725 243.100 56.745 ;
        POLYGON 241.480 56.725 241.480 56.710 241.465 56.710 ;
        RECT 241.480 56.710 243.100 56.725 ;
        POLYGON 241.465 56.710 241.465 56.585 241.380 56.585 ;
        RECT 241.465 56.700 243.100 56.710 ;
        POLYGON 243.100 56.745 243.145 56.745 243.100 56.700 ;
        POLYGON 244.540 56.745 244.540 56.700 244.495 56.700 ;
        RECT 244.540 56.700 245.660 56.745 ;
        RECT 241.465 56.630 243.040 56.700 ;
        POLYGON 243.040 56.700 243.100 56.700 243.040 56.630 ;
        POLYGON 244.495 56.700 244.495 56.660 244.450 56.660 ;
        RECT 244.495 56.695 245.660 56.700 ;
        POLYGON 245.660 56.790 245.790 56.790 245.660 56.695 ;
        POLYGON 247.415 56.790 247.415 56.755 247.330 56.755 ;
        RECT 247.415 56.785 249.930 56.790 ;
        POLYGON 249.930 56.790 250.040 56.790 249.930 56.785 ;
        POLYGON 250.640 56.790 250.690 56.790 250.690 56.785 ;
        RECT 250.690 56.785 253.085 56.790 ;
        RECT 247.415 56.780 249.845 56.785 ;
        POLYGON 249.845 56.785 249.915 56.785 249.845 56.780 ;
        POLYGON 250.705 56.785 250.780 56.785 250.780 56.780 ;
        RECT 250.780 56.780 253.085 56.785 ;
        RECT 247.415 56.775 249.785 56.780 ;
        POLYGON 249.785 56.780 249.845 56.780 249.785 56.775 ;
        POLYGON 250.780 56.780 250.860 56.780 250.860 56.775 ;
        RECT 250.860 56.775 253.085 56.780 ;
        RECT 247.415 56.760 249.655 56.775 ;
        POLYGON 249.655 56.775 249.770 56.775 249.655 56.760 ;
        POLYGON 250.860 56.775 250.920 56.775 250.920 56.770 ;
        RECT 250.920 56.770 253.085 56.775 ;
        POLYGON 250.930 56.770 250.960 56.770 250.960 56.765 ;
        RECT 250.960 56.765 253.085 56.770 ;
        POLYGON 250.965 56.765 251.015 56.765 251.015 56.760 ;
        RECT 251.015 56.760 253.085 56.765 ;
        RECT 247.415 56.755 249.515 56.760 ;
        POLYGON 247.330 56.755 247.330 56.720 247.250 56.720 ;
        RECT 247.330 56.745 249.515 56.755 ;
        POLYGON 249.515 56.760 249.650 56.760 249.515 56.745 ;
        POLYGON 251.015 56.760 251.125 56.760 251.125 56.750 ;
        RECT 251.125 56.750 253.085 56.760 ;
        POLYGON 251.135 56.750 251.175 56.750 251.175 56.745 ;
        RECT 251.175 56.745 253.085 56.750 ;
        RECT 247.330 56.730 249.390 56.745 ;
        POLYGON 249.390 56.745 249.495 56.745 249.390 56.730 ;
        POLYGON 251.175 56.745 251.215 56.745 251.215 56.740 ;
        RECT 251.215 56.740 253.085 56.745 ;
        POLYGON 251.220 56.740 251.225 56.740 251.225 56.735 ;
        RECT 251.225 56.735 253.085 56.740 ;
        POLYGON 253.085 56.820 253.260 56.735 253.085 56.735 ;
        POLYGON 254.550 56.820 254.615 56.820 254.615 56.780 ;
        RECT 254.615 56.780 256.015 56.820 ;
        POLYGON 254.615 56.780 254.630 56.780 254.630 56.770 ;
        RECT 254.630 56.770 256.015 56.780 ;
        POLYGON 254.630 56.770 254.680 56.770 254.680 56.735 ;
        RECT 254.680 56.735 256.015 56.770 ;
        POLYGON 251.225 56.735 251.275 56.735 251.275 56.730 ;
        RECT 251.275 56.730 253.260 56.735 ;
        RECT 247.330 56.725 249.385 56.730 ;
        POLYGON 249.385 56.730 249.390 56.730 249.385 56.725 ;
        POLYGON 251.275 56.730 251.305 56.730 251.305 56.725 ;
        RECT 251.305 56.725 253.260 56.730 ;
        RECT 247.330 56.720 249.240 56.725 ;
        POLYGON 247.250 56.720 247.250 56.695 247.205 56.695 ;
        RECT 247.250 56.705 249.240 56.720 ;
        POLYGON 249.240 56.725 249.385 56.725 249.240 56.705 ;
        POLYGON 251.305 56.725 251.395 56.725 251.395 56.710 ;
        RECT 251.395 56.710 253.260 56.725 ;
        POLYGON 251.405 56.710 251.430 56.710 251.430 56.705 ;
        RECT 251.430 56.705 253.260 56.710 ;
        RECT 247.250 56.695 249.190 56.705 ;
        POLYGON 249.190 56.705 249.225 56.705 249.190 56.695 ;
        POLYGON 251.430 56.705 251.485 56.705 251.485 56.695 ;
        RECT 251.485 56.695 253.260 56.705 ;
        RECT 244.495 56.660 245.560 56.695 ;
        POLYGON 244.450 56.660 244.450 56.640 244.425 56.640 ;
        RECT 244.450 56.640 245.560 56.660 ;
        POLYGON 244.425 56.640 244.425 56.630 244.415 56.630 ;
        RECT 244.425 56.630 245.560 56.640 ;
        RECT 241.465 56.585 242.880 56.630 ;
        RECT 237.335 56.575 239.550 56.585 ;
        POLYGON 239.550 56.585 239.560 56.585 239.550 56.575 ;
        POLYGON 241.380 56.585 241.380 56.575 241.375 56.575 ;
        RECT 241.380 56.575 242.880 56.585 ;
        RECT 237.335 56.565 239.545 56.575 ;
        POLYGON 239.545 56.575 239.550 56.575 239.545 56.565 ;
        POLYGON 241.375 56.575 241.375 56.570 241.370 56.570 ;
        RECT 241.375 56.570 242.880 56.575 ;
        RECT 237.335 56.520 239.450 56.565 ;
        RECT 229.745 56.485 234.080 56.520 ;
        POLYGON 234.080 56.520 234.095 56.520 234.080 56.485 ;
        POLYGON 237.220 56.520 237.220 56.485 237.205 56.485 ;
        RECT 237.220 56.485 239.450 56.520 ;
        RECT 229.745 56.245 234.010 56.485 ;
        POLYGON 234.010 56.485 234.080 56.485 234.010 56.245 ;
        POLYGON 237.205 56.485 237.205 56.320 237.135 56.320 ;
        RECT 237.205 56.385 239.450 56.485 ;
        POLYGON 239.450 56.565 239.545 56.565 239.450 56.385 ;
        POLYGON 241.370 56.565 241.370 56.455 241.295 56.455 ;
        RECT 241.370 56.455 242.880 56.570 ;
        POLYGON 241.295 56.455 241.295 56.425 241.270 56.425 ;
        RECT 241.295 56.450 242.880 56.455 ;
        POLYGON 242.880 56.630 243.040 56.630 242.880 56.450 ;
        POLYGON 244.415 56.630 244.415 56.560 244.340 56.560 ;
        RECT 244.415 56.620 245.560 56.630 ;
        POLYGON 245.560 56.695 245.660 56.695 245.560 56.620 ;
        POLYGON 247.205 56.695 247.205 56.690 247.195 56.690 ;
        RECT 247.205 56.690 249.120 56.695 ;
        POLYGON 247.195 56.690 247.195 56.635 247.075 56.635 ;
        RECT 247.195 56.685 249.120 56.690 ;
        POLYGON 249.120 56.695 249.190 56.695 249.120 56.685 ;
        POLYGON 251.485 56.695 251.535 56.695 251.535 56.685 ;
        RECT 251.535 56.690 253.260 56.695 ;
        POLYGON 253.260 56.735 253.355 56.690 253.260 56.690 ;
        POLYGON 254.680 56.735 254.710 56.735 254.710 56.715 ;
        RECT 254.710 56.715 256.015 56.735 ;
        POLYGON 254.710 56.715 254.745 56.715 254.745 56.690 ;
        RECT 254.745 56.690 256.015 56.715 ;
        RECT 251.535 56.685 253.360 56.690 ;
        RECT 247.195 56.655 248.975 56.685 ;
        POLYGON 248.975 56.685 249.120 56.685 248.975 56.655 ;
        POLYGON 251.535 56.685 251.610 56.685 251.610 56.670 ;
        RECT 251.610 56.670 253.360 56.685 ;
        POLYGON 251.610 56.670 251.655 56.670 251.655 56.665 ;
        RECT 251.655 56.665 253.360 56.670 ;
        POLYGON 251.660 56.665 251.700 56.665 251.700 56.655 ;
        RECT 251.700 56.655 253.360 56.665 ;
        RECT 247.195 56.650 248.950 56.655 ;
        POLYGON 248.950 56.655 248.975 56.655 248.950 56.650 ;
        POLYGON 251.700 56.655 251.720 56.655 251.720 56.650 ;
        RECT 251.720 56.650 253.360 56.655 ;
        RECT 247.195 56.635 248.875 56.650 ;
        POLYGON 248.875 56.650 248.945 56.650 248.875 56.635 ;
        POLYGON 251.720 56.650 251.740 56.650 251.740 56.645 ;
        RECT 251.740 56.645 253.360 56.650 ;
        POLYGON 251.745 56.645 251.785 56.645 251.785 56.635 ;
        RECT 251.785 56.635 253.360 56.645 ;
        POLYGON 247.075 56.635 247.075 56.620 247.045 56.620 ;
        RECT 247.075 56.630 248.850 56.635 ;
        POLYGON 248.850 56.635 248.875 56.635 248.850 56.630 ;
        POLYGON 251.785 56.635 251.810 56.635 251.810 56.630 ;
        RECT 251.810 56.630 253.360 56.635 ;
        RECT 247.075 56.620 248.710 56.630 ;
        RECT 244.415 56.560 245.445 56.620 ;
        POLYGON 244.340 56.560 244.340 56.450 244.230 56.450 ;
        RECT 244.340 56.535 245.445 56.560 ;
        POLYGON 245.445 56.620 245.560 56.620 245.445 56.535 ;
        POLYGON 247.045 56.620 247.045 56.590 246.985 56.590 ;
        RECT 247.045 56.595 248.710 56.620 ;
        POLYGON 248.710 56.630 248.850 56.630 248.710 56.595 ;
        POLYGON 251.810 56.630 251.920 56.630 251.920 56.605 ;
        RECT 251.920 56.615 253.360 56.630 ;
        POLYGON 253.360 56.690 253.505 56.615 253.360 56.615 ;
        POLYGON 254.745 56.690 254.850 56.690 254.850 56.615 ;
        RECT 254.850 56.680 256.015 56.690 ;
        POLYGON 256.015 56.840 256.200 56.680 256.015 56.680 ;
        POLYGON 257.655 56.840 257.795 56.840 257.795 56.695 ;
        RECT 257.795 56.770 259.495 56.840 ;
        POLYGON 259.495 56.925 259.620 56.770 259.495 56.770 ;
        POLYGON 261.775 56.925 261.790 56.925 261.790 56.905 ;
        RECT 261.790 56.920 264.720 56.925 ;
        POLYGON 264.720 56.980 264.755 56.920 264.720 56.920 ;
        POLYGON 269.100 56.980 269.125 56.980 269.125 56.925 ;
        RECT 269.125 56.920 276.115 56.980 ;
        RECT 261.790 56.905 264.755 56.920 ;
        POLYGON 261.790 56.905 261.795 56.905 261.795 56.900 ;
        RECT 261.795 56.900 264.755 56.905 ;
        POLYGON 261.795 56.900 261.840 56.900 261.840 56.830 ;
        RECT 261.840 56.830 264.755 56.900 ;
        POLYGON 261.840 56.830 261.850 56.830 261.850 56.810 ;
        RECT 261.850 56.810 264.755 56.830 ;
        POLYGON 261.850 56.810 261.880 56.810 261.880 56.770 ;
        RECT 261.880 56.770 264.755 56.810 ;
        RECT 257.795 56.720 259.620 56.770 ;
        POLYGON 259.620 56.770 259.655 56.720 259.620 56.720 ;
        POLYGON 261.880 56.770 261.910 56.770 261.910 56.720 ;
        RECT 261.910 56.720 264.755 56.770 ;
        RECT 257.795 56.695 259.655 56.720 ;
        POLYGON 257.795 56.695 257.810 56.695 257.810 56.680 ;
        RECT 257.810 56.680 259.655 56.695 ;
        RECT 254.850 56.670 256.200 56.680 ;
        POLYGON 256.200 56.680 256.215 56.670 256.200 56.670 ;
        POLYGON 257.810 56.680 257.820 56.680 257.820 56.670 ;
        RECT 257.820 56.670 259.655 56.680 ;
        RECT 254.850 56.625 256.215 56.670 ;
        POLYGON 256.215 56.670 256.265 56.625 256.215 56.625 ;
        POLYGON 257.820 56.670 257.830 56.670 257.830 56.660 ;
        RECT 257.830 56.660 259.655 56.670 ;
        POLYGON 257.830 56.660 257.860 56.660 257.860 56.625 ;
        RECT 257.860 56.625 259.655 56.660 ;
        RECT 254.850 56.615 256.265 56.625 ;
        POLYGON 256.265 56.625 256.275 56.615 256.265 56.615 ;
        POLYGON 257.860 56.625 257.870 56.625 257.870 56.615 ;
        RECT 257.870 56.615 259.655 56.625 ;
        RECT 251.920 56.605 253.505 56.615 ;
        POLYGON 251.920 56.605 251.935 56.605 251.935 56.600 ;
        RECT 251.935 56.600 253.505 56.605 ;
        POLYGON 251.935 56.600 251.955 56.600 251.955 56.595 ;
        RECT 251.955 56.595 253.505 56.600 ;
        RECT 247.045 56.590 248.665 56.595 ;
        POLYGON 246.980 56.590 246.980 56.585 246.970 56.585 ;
        RECT 246.980 56.585 248.665 56.590 ;
        POLYGON 248.665 56.595 248.710 56.595 248.665 56.585 ;
        POLYGON 251.955 56.595 251.995 56.595 251.995 56.585 ;
        RECT 251.995 56.585 253.505 56.595 ;
        POLYGON 246.970 56.585 246.970 56.535 246.875 56.535 ;
        RECT 246.970 56.565 248.590 56.585 ;
        POLYGON 248.590 56.585 248.665 56.585 248.590 56.565 ;
        RECT 252.000 56.580 253.505 56.585 ;
        POLYGON 252.000 56.580 252.055 56.580 252.055 56.565 ;
        RECT 252.055 56.575 253.505 56.580 ;
        POLYGON 253.505 56.615 253.580 56.575 253.505 56.575 ;
        POLYGON 254.850 56.615 254.860 56.615 254.860 56.605 ;
        RECT 254.860 56.605 256.275 56.615 ;
        POLYGON 254.860 56.605 254.900 56.605 254.900 56.575 ;
        RECT 254.900 56.575 256.275 56.605 ;
        RECT 252.055 56.565 253.580 56.575 ;
        RECT 246.970 56.560 248.585 56.565 ;
        RECT 246.970 56.555 248.565 56.560 ;
        POLYGON 248.565 56.560 248.585 56.560 248.565 56.555 ;
        POLYGON 252.055 56.565 252.095 56.565 252.095 56.555 ;
        RECT 252.095 56.555 253.580 56.565 ;
        RECT 246.970 56.535 248.455 56.555 ;
        RECT 244.340 56.530 245.440 56.535 ;
        POLYGON 245.440 56.535 245.445 56.535 245.440 56.530 ;
        POLYGON 246.875 56.535 246.875 56.530 246.865 56.530 ;
        RECT 246.875 56.530 248.455 56.535 ;
        RECT 244.340 56.485 245.380 56.530 ;
        POLYGON 245.380 56.530 245.440 56.530 245.380 56.485 ;
        POLYGON 246.865 56.530 246.865 56.490 246.790 56.490 ;
        RECT 246.865 56.525 248.455 56.530 ;
        POLYGON 248.455 56.555 248.565 56.555 248.455 56.525 ;
        POLYGON 252.095 56.555 252.175 56.555 252.175 56.535 ;
        RECT 252.175 56.550 253.580 56.555 ;
        POLYGON 253.580 56.575 253.620 56.550 253.580 56.550 ;
        POLYGON 254.900 56.575 254.935 56.575 254.935 56.550 ;
        RECT 254.935 56.550 256.275 56.575 ;
        RECT 252.175 56.535 253.620 56.550 ;
        POLYGON 252.175 56.535 252.205 56.535 252.205 56.525 ;
        RECT 252.205 56.525 253.620 56.535 ;
        RECT 246.865 56.505 248.390 56.525 ;
        POLYGON 248.390 56.525 248.455 56.525 248.390 56.510 ;
        POLYGON 252.205 56.525 252.245 56.525 252.245 56.515 ;
        RECT 252.245 56.515 253.620 56.525 ;
        POLYGON 253.620 56.550 253.685 56.515 253.620 56.515 ;
        POLYGON 254.935 56.550 254.940 56.550 254.940 56.545 ;
        RECT 254.940 56.545 256.275 56.550 ;
        POLYGON 254.940 56.545 254.975 56.545 254.975 56.515 ;
        RECT 254.975 56.515 256.275 56.545 ;
        POLYGON 252.245 56.515 252.250 56.515 252.250 56.510 ;
        RECT 252.250 56.510 253.685 56.515 ;
        RECT 246.865 56.490 248.320 56.505 ;
        POLYGON 246.790 56.490 246.790 56.485 246.780 56.485 ;
        RECT 246.790 56.485 248.320 56.490 ;
        POLYGON 248.320 56.505 248.390 56.505 248.320 56.485 ;
        POLYGON 252.255 56.510 252.330 56.510 252.330 56.485 ;
        RECT 252.330 56.485 253.685 56.510 ;
        RECT 244.340 56.450 245.335 56.485 ;
        RECT 241.295 56.425 242.860 56.450 ;
        POLYGON 242.860 56.450 242.880 56.450 242.860 56.425 ;
        POLYGON 244.230 56.450 244.230 56.425 244.205 56.425 ;
        RECT 244.230 56.445 245.335 56.450 ;
        POLYGON 245.335 56.485 245.380 56.485 245.335 56.445 ;
        POLYGON 246.780 56.485 246.780 56.465 246.740 56.465 ;
        RECT 246.780 56.470 248.265 56.485 ;
        POLYGON 248.265 56.485 248.320 56.485 248.265 56.470 ;
        POLYGON 252.330 56.485 252.375 56.485 252.375 56.470 ;
        RECT 252.375 56.475 253.685 56.485 ;
        POLYGON 253.685 56.515 253.750 56.475 253.685 56.475 ;
        POLYGON 254.975 56.515 255.030 56.515 255.030 56.475 ;
        RECT 255.030 56.475 256.275 56.515 ;
        RECT 252.375 56.470 253.750 56.475 ;
        RECT 246.780 56.465 248.200 56.470 ;
        POLYGON 246.740 56.465 246.740 56.445 246.705 56.445 ;
        RECT 246.740 56.445 248.200 56.465 ;
        POLYGON 248.200 56.470 248.265 56.470 248.200 56.445 ;
        POLYGON 252.375 56.470 252.395 56.470 252.395 56.465 ;
        RECT 252.395 56.465 253.750 56.470 ;
        POLYGON 252.395 56.465 252.430 56.465 252.430 56.450 ;
        RECT 252.430 56.450 253.750 56.465 ;
        POLYGON 253.750 56.475 253.800 56.450 253.750 56.450 ;
        POLYGON 255.030 56.475 255.060 56.475 255.060 56.450 ;
        RECT 255.060 56.450 256.275 56.475 ;
        POLYGON 252.435 56.450 252.450 56.450 252.450 56.445 ;
        RECT 252.450 56.445 253.800 56.450 ;
        RECT 244.230 56.425 245.250 56.445 ;
        POLYGON 241.270 56.425 241.270 56.385 241.245 56.385 ;
        RECT 241.270 56.415 242.850 56.425 ;
        POLYGON 242.850 56.425 242.860 56.425 242.850 56.415 ;
        POLYGON 244.205 56.425 244.205 56.415 244.195 56.415 ;
        RECT 244.205 56.415 245.250 56.425 ;
        RECT 241.270 56.400 242.840 56.415 ;
        POLYGON 242.840 56.415 242.850 56.415 242.840 56.400 ;
        POLYGON 244.195 56.415 244.195 56.400 244.180 56.400 ;
        RECT 244.195 56.400 245.250 56.415 ;
        RECT 241.270 56.385 242.685 56.400 ;
        RECT 237.205 56.320 239.340 56.385 ;
        POLYGON 237.135 56.320 237.135 56.245 237.100 56.245 ;
        RECT 237.135 56.245 239.340 56.320 ;
        RECT 229.745 55.655 233.815 56.245 ;
        RECT 181.815 55.640 196.020 55.645 ;
        POLYGON 196.020 55.645 196.025 55.640 196.020 55.640 ;
        RECT 206.270 55.640 222.225 55.655 ;
        RECT 170.610 55.260 174.845 55.275 ;
        POLYGON 174.845 55.275 174.855 55.260 174.845 55.260 ;
        RECT 181.815 55.260 196.025 55.640 ;
        RECT 170.610 55.060 174.855 55.260 ;
        POLYGON 174.855 55.260 174.925 55.060 174.855 55.060 ;
        POLYGON 181.815 55.260 181.875 55.260 181.875 55.065 ;
        RECT 181.875 55.060 196.025 55.260 ;
        RECT 170.610 54.995 174.925 55.060 ;
        RECT 165.765 54.945 167.840 54.995 ;
        POLYGON 167.840 54.995 167.865 54.945 167.840 54.945 ;
        POLYGON 170.610 54.995 170.630 54.995 170.630 54.955 ;
        RECT 170.630 54.945 174.925 54.995 ;
        RECT 165.765 54.920 167.865 54.945 ;
        RECT 160.760 54.870 161.645 54.910 ;
        RECT 159.180 54.865 160.005 54.870 ;
        POLYGON 159.180 54.865 159.195 54.865 159.195 54.850 ;
        RECT 159.195 54.850 160.005 54.865 ;
        RECT 157.685 54.845 158.385 54.850 ;
        POLYGON 157.685 54.845 157.690 54.845 157.690 54.840 ;
        RECT 157.690 54.840 158.385 54.845 ;
        RECT 152.535 54.835 155.635 54.840 ;
        POLYGON 155.635 54.840 155.650 54.835 155.635 54.835 ;
        POLYGON 157.690 54.840 157.700 54.840 157.700 54.835 ;
        RECT 157.700 54.835 158.385 54.840 ;
        RECT 152.535 54.825 155.650 54.835 ;
        POLYGON 155.650 54.835 155.695 54.825 155.650 54.825 ;
        POLYGON 157.700 54.835 157.715 54.835 157.715 54.825 ;
        RECT 157.715 54.825 158.385 54.835 ;
        POLYGON 152.505 54.825 152.505 54.760 152.400 54.760 ;
        RECT 152.505 54.810 155.695 54.825 ;
        POLYGON 155.695 54.825 155.755 54.810 155.695 54.810 ;
        POLYGON 157.715 54.825 157.735 54.825 157.735 54.810 ;
        RECT 157.735 54.810 158.385 54.825 ;
        RECT 152.505 54.800 155.755 54.810 ;
        POLYGON 155.755 54.810 155.805 54.800 155.755 54.800 ;
        POLYGON 157.735 54.810 157.750 54.810 157.750 54.800 ;
        RECT 157.750 54.800 158.385 54.810 ;
        RECT 152.505 54.795 155.805 54.800 ;
        POLYGON 155.805 54.800 155.815 54.795 155.805 54.795 ;
        POLYGON 157.750 54.800 157.760 54.800 157.760 54.795 ;
        RECT 157.760 54.795 158.385 54.800 ;
        RECT 152.505 54.780 155.820 54.795 ;
        POLYGON 155.820 54.795 155.875 54.780 155.820 54.780 ;
        POLYGON 157.760 54.795 157.785 54.795 157.785 54.780 ;
        RECT 157.785 54.780 158.385 54.795 ;
        RECT 152.505 54.770 155.875 54.780 ;
        POLYGON 155.875 54.780 155.935 54.770 155.875 54.770 ;
        POLYGON 157.785 54.780 157.800 54.780 157.800 54.770 ;
        RECT 157.800 54.770 158.385 54.780 ;
        RECT 152.505 54.765 155.950 54.770 ;
        POLYGON 155.950 54.770 155.970 54.765 155.950 54.765 ;
        POLYGON 157.800 54.770 157.810 54.770 157.810 54.765 ;
        RECT 157.810 54.765 158.385 54.770 ;
        RECT 152.505 54.760 155.970 54.765 ;
        POLYGON 152.400 54.760 152.400 54.750 152.385 54.750 ;
        RECT 152.400 54.750 155.970 54.760 ;
        RECT 150.370 54.730 150.920 54.750 ;
        POLYGON 150.920 54.750 150.945 54.750 150.920 54.730 ;
        POLYGON 152.385 54.750 152.385 54.730 152.355 54.730 ;
        RECT 152.385 54.745 155.970 54.750 ;
        POLYGON 155.970 54.765 156.085 54.745 155.970 54.745 ;
        POLYGON 157.815 54.765 157.845 54.765 157.845 54.745 ;
        RECT 157.845 54.760 158.385 54.765 ;
        POLYGON 158.385 54.850 158.510 54.760 158.385 54.760 ;
        POLYGON 159.195 54.850 159.290 54.850 159.290 54.760 ;
        RECT 159.290 54.760 160.005 54.850 ;
        RECT 157.845 54.745 158.510 54.760 ;
        RECT 152.385 54.740 156.085 54.745 ;
        POLYGON 156.085 54.745 156.115 54.740 156.085 54.740 ;
        POLYGON 157.845 54.745 157.850 54.745 157.850 54.740 ;
        RECT 157.850 54.740 158.510 54.745 ;
        RECT 152.385 54.735 156.120 54.740 ;
        POLYGON 156.120 54.740 156.130 54.735 156.120 54.735 ;
        POLYGON 157.850 54.740 157.860 54.740 157.860 54.735 ;
        RECT 157.860 54.735 158.510 54.740 ;
        RECT 152.385 54.730 156.135 54.735 ;
        RECT 150.370 54.695 150.870 54.730 ;
        RECT 148.715 54.685 149.550 54.695 ;
        RECT 148.690 54.680 149.550 54.685 ;
        POLYGON 149.550 54.695 149.565 54.695 149.550 54.680 ;
        POLYGON 150.310 54.695 150.310 54.680 150.295 54.680 ;
        RECT 150.310 54.680 150.870 54.695 ;
        POLYGON 150.870 54.730 150.920 54.730 150.870 54.680 ;
        POLYGON 152.355 54.730 152.355 54.725 152.350 54.725 ;
        RECT 152.355 54.725 156.135 54.730 ;
        POLYGON 152.350 54.725 152.350 54.695 152.310 54.695 ;
        RECT 152.350 54.720 156.135 54.725 ;
        POLYGON 156.135 54.735 156.225 54.720 156.135 54.720 ;
        POLYGON 157.860 54.735 157.885 54.735 157.885 54.720 ;
        RECT 157.885 54.720 158.510 54.735 ;
        RECT 152.350 54.705 156.225 54.720 ;
        POLYGON 156.225 54.720 156.285 54.705 156.225 54.705 ;
        POLYGON 157.885 54.720 157.905 54.720 157.905 54.705 ;
        RECT 157.905 54.710 158.510 54.720 ;
        POLYGON 158.510 54.760 158.580 54.710 158.510 54.710 ;
        POLYGON 159.290 54.760 159.300 54.760 159.300 54.755 ;
        RECT 159.300 54.755 160.005 54.760 ;
        POLYGON 159.300 54.755 159.345 54.755 159.345 54.710 ;
        RECT 159.345 54.725 160.005 54.755 ;
        POLYGON 160.005 54.870 160.145 54.725 160.005 54.725 ;
        POLYGON 160.760 54.870 160.860 54.870 160.860 54.760 ;
        RECT 160.860 54.760 161.645 54.870 ;
        POLYGON 160.860 54.760 160.880 54.760 160.880 54.735 ;
        RECT 160.880 54.735 161.645 54.760 ;
        POLYGON 160.880 54.735 160.885 54.735 160.885 54.725 ;
        RECT 160.885 54.725 161.645 54.735 ;
        RECT 159.345 54.710 160.145 54.725 ;
        RECT 157.905 54.705 158.580 54.710 ;
        RECT 152.350 54.695 156.300 54.705 ;
        POLYGON 152.310 54.695 152.310 54.685 152.290 54.685 ;
        RECT 152.310 54.690 156.300 54.695 ;
        POLYGON 156.300 54.705 156.365 54.690 156.300 54.690 ;
        POLYGON 157.905 54.705 157.930 54.705 157.930 54.690 ;
        RECT 157.930 54.690 158.580 54.705 ;
        RECT 152.310 54.685 156.365 54.690 ;
        POLYGON 152.290 54.685 152.290 54.680 152.285 54.680 ;
        RECT 152.290 54.680 156.365 54.685 ;
        RECT 117.275 54.605 147.715 54.680 ;
        POLYGON 147.715 54.680 147.760 54.680 147.715 54.605 ;
        POLYGON 148.690 54.680 148.690 54.640 148.660 54.640 ;
        RECT 148.690 54.650 149.525 54.680 ;
        POLYGON 149.525 54.680 149.550 54.680 149.525 54.650 ;
        POLYGON 150.295 54.680 150.295 54.655 150.270 54.655 ;
        RECT 150.295 54.655 150.735 54.680 ;
        RECT 148.690 54.640 149.395 54.650 ;
        POLYGON 148.660 54.640 148.660 54.610 148.640 54.610 ;
        RECT 148.660 54.610 149.395 54.640 ;
        RECT 117.275 54.540 147.675 54.605 ;
        POLYGON 147.675 54.605 147.715 54.605 147.675 54.540 ;
        POLYGON 148.640 54.605 148.640 54.540 148.595 54.540 ;
        RECT 148.640 54.540 149.395 54.610 ;
        RECT 117.275 54.420 147.610 54.540 ;
        POLYGON 147.610 54.540 147.675 54.540 147.610 54.420 ;
        POLYGON 148.595 54.535 148.595 54.465 148.550 54.465 ;
        RECT 148.595 54.485 149.395 54.540 ;
        POLYGON 149.395 54.650 149.525 54.650 149.395 54.485 ;
        POLYGON 150.270 54.650 150.270 54.615 150.235 54.615 ;
        RECT 150.270 54.615 150.735 54.655 ;
        POLYGON 150.235 54.615 150.235 54.565 150.190 54.565 ;
        RECT 150.235 54.565 150.735 54.615 ;
        POLYGON 150.190 54.565 150.190 54.485 150.115 54.485 ;
        RECT 150.190 54.550 150.735 54.565 ;
        POLYGON 150.735 54.680 150.870 54.680 150.735 54.550 ;
        POLYGON 152.285 54.680 152.285 54.580 152.135 54.580 ;
        RECT 152.285 54.670 156.365 54.680 ;
        POLYGON 156.365 54.690 156.440 54.670 156.365 54.670 ;
        POLYGON 157.930 54.690 157.945 54.690 157.945 54.680 ;
        RECT 157.945 54.680 158.580 54.690 ;
        POLYGON 157.945 54.680 157.955 54.680 157.955 54.675 ;
        RECT 157.955 54.675 158.580 54.680 ;
        POLYGON 157.960 54.675 157.965 54.675 157.965 54.670 ;
        RECT 157.965 54.670 158.580 54.675 ;
        RECT 152.285 54.660 156.440 54.670 ;
        POLYGON 156.440 54.670 156.480 54.660 156.440 54.660 ;
        POLYGON 157.965 54.670 157.980 54.670 157.980 54.660 ;
        RECT 157.980 54.665 158.580 54.670 ;
        POLYGON 158.580 54.710 158.640 54.665 158.580 54.665 ;
        POLYGON 159.345 54.710 159.390 54.710 159.390 54.665 ;
        RECT 159.390 54.705 160.145 54.710 ;
        POLYGON 160.145 54.725 160.165 54.705 160.145 54.705 ;
        RECT 159.390 54.665 160.165 54.705 ;
        POLYGON 160.885 54.725 160.910 54.725 160.910 54.700 ;
        RECT 160.910 54.700 161.645 54.725 ;
        RECT 157.980 54.660 158.640 54.665 ;
        RECT 152.285 54.650 156.480 54.660 ;
        POLYGON 156.480 54.660 156.505 54.650 156.480 54.650 ;
        POLYGON 157.980 54.660 157.990 54.660 157.990 54.650 ;
        RECT 157.990 54.655 158.640 54.660 ;
        POLYGON 158.640 54.665 158.650 54.655 158.640 54.655 ;
        POLYGON 159.390 54.665 159.405 54.665 159.405 54.655 ;
        RECT 159.405 54.660 160.165 54.665 ;
        POLYGON 160.165 54.700 160.205 54.660 160.165 54.660 ;
        POLYGON 160.910 54.700 160.925 54.700 160.925 54.685 ;
        RECT 160.925 54.685 161.645 54.700 ;
        POLYGON 160.925 54.685 160.940 54.685 160.940 54.665 ;
        RECT 160.940 54.660 161.645 54.685 ;
        RECT 159.405 54.655 160.205 54.660 ;
        RECT 157.990 54.650 158.650 54.655 ;
        RECT 152.285 54.625 156.505 54.650 ;
        POLYGON 156.505 54.650 156.585 54.625 156.505 54.625 ;
        POLYGON 157.990 54.650 158.025 54.650 158.025 54.625 ;
        RECT 158.025 54.625 158.650 54.650 ;
        RECT 152.285 54.605 156.595 54.625 ;
        POLYGON 156.595 54.625 156.650 54.605 156.595 54.605 ;
        POLYGON 158.025 54.625 158.050 54.625 158.050 54.610 ;
        RECT 158.050 54.610 158.650 54.625 ;
        POLYGON 158.050 54.610 158.055 54.610 158.055 54.605 ;
        RECT 158.055 54.605 158.650 54.610 ;
        RECT 152.285 54.600 156.650 54.605 ;
        POLYGON 156.650 54.605 156.660 54.600 156.650 54.600 ;
        POLYGON 158.055 54.605 158.060 54.605 158.060 54.600 ;
        RECT 158.060 54.600 158.650 54.605 ;
        RECT 152.285 54.585 156.665 54.600 ;
        POLYGON 156.665 54.600 156.715 54.585 156.665 54.585 ;
        POLYGON 158.060 54.600 158.085 54.600 158.085 54.585 ;
        RECT 158.085 54.585 158.650 54.600 ;
        RECT 152.285 54.580 156.715 54.585 ;
        POLYGON 152.135 54.580 152.135 54.550 152.095 54.550 ;
        RECT 152.135 54.570 156.715 54.580 ;
        POLYGON 156.715 54.585 156.750 54.570 156.715 54.570 ;
        POLYGON 158.085 54.585 158.105 54.585 158.105 54.570 ;
        RECT 158.105 54.570 158.650 54.585 ;
        RECT 152.135 54.555 156.750 54.570 ;
        POLYGON 156.750 54.570 156.795 54.555 156.750 54.555 ;
        POLYGON 158.105 54.570 158.125 54.570 158.125 54.555 ;
        RECT 158.125 54.555 158.650 54.570 ;
        RECT 152.135 54.550 156.795 54.555 ;
        RECT 150.190 54.510 150.695 54.550 ;
        POLYGON 150.695 54.550 150.735 54.550 150.695 54.510 ;
        POLYGON 152.095 54.550 152.095 54.510 152.045 54.510 ;
        RECT 152.095 54.535 156.795 54.550 ;
        POLYGON 156.795 54.555 156.840 54.535 156.795 54.535 ;
        POLYGON 158.125 54.555 158.155 54.555 158.155 54.535 ;
        RECT 158.155 54.550 158.650 54.555 ;
        POLYGON 158.650 54.655 158.790 54.550 158.650 54.550 ;
        POLYGON 159.405 54.655 159.440 54.655 159.440 54.625 ;
        RECT 159.440 54.625 160.205 54.655 ;
        POLYGON 159.440 54.625 159.465 54.625 159.465 54.600 ;
        RECT 159.465 54.600 160.205 54.625 ;
        POLYGON 159.465 54.600 159.510 54.600 159.510 54.550 ;
        RECT 159.510 54.550 160.205 54.600 ;
        RECT 158.155 54.535 158.790 54.550 ;
        RECT 152.095 54.510 156.845 54.535 ;
        POLYGON 156.845 54.535 156.905 54.510 156.845 54.510 ;
        POLYGON 158.155 54.535 158.190 54.535 158.190 54.510 ;
        RECT 158.190 54.510 158.790 54.535 ;
        RECT 150.190 54.485 150.615 54.510 ;
        RECT 148.595 54.470 149.385 54.485 ;
        POLYGON 149.385 54.485 149.395 54.485 149.385 54.470 ;
        POLYGON 150.115 54.485 150.115 54.475 150.105 54.475 ;
        RECT 150.115 54.475 150.615 54.485 ;
        RECT 148.595 54.465 149.350 54.470 ;
        POLYGON 148.550 54.465 148.550 54.425 148.525 54.425 ;
        RECT 148.550 54.425 149.350 54.465 ;
        RECT 148.525 54.420 149.350 54.425 ;
        POLYGON 149.350 54.470 149.385 54.470 149.350 54.420 ;
        POLYGON 150.105 54.470 150.105 54.420 150.055 54.420 ;
        RECT 150.105 54.425 150.615 54.475 ;
        POLYGON 150.615 54.510 150.695 54.510 150.615 54.425 ;
        POLYGON 152.045 54.510 152.045 54.465 151.985 54.465 ;
        RECT 152.045 54.480 156.905 54.510 ;
        POLYGON 156.905 54.510 156.975 54.480 156.905 54.480 ;
        POLYGON 158.190 54.510 158.215 54.510 158.215 54.495 ;
        RECT 158.215 54.495 158.790 54.510 ;
        POLYGON 158.215 54.495 158.230 54.495 158.230 54.485 ;
        RECT 158.230 54.485 158.790 54.495 ;
        POLYGON 158.230 54.485 158.240 54.485 158.240 54.480 ;
        RECT 158.240 54.480 158.790 54.485 ;
        RECT 152.045 54.465 156.975 54.480 ;
        POLYGON 151.985 54.465 151.985 54.430 151.940 54.430 ;
        RECT 151.985 54.460 156.975 54.465 ;
        POLYGON 156.975 54.480 157.020 54.460 156.975 54.460 ;
        POLYGON 158.240 54.480 158.265 54.480 158.265 54.460 ;
        RECT 158.265 54.470 158.790 54.480 ;
        POLYGON 158.790 54.550 158.885 54.470 158.790 54.470 ;
        POLYGON 159.510 54.550 159.590 54.550 159.590 54.470 ;
        RECT 159.590 54.505 160.205 54.550 ;
        POLYGON 160.205 54.660 160.345 54.505 160.205 54.505 ;
        POLYGON 160.940 54.660 161.065 54.660 161.065 54.510 ;
        RECT 161.065 54.650 161.645 54.660 ;
        POLYGON 161.645 54.910 161.850 54.650 161.645 54.650 ;
        RECT 162.825 54.905 164.155 54.920 ;
        POLYGON 162.825 54.905 162.960 54.905 162.960 54.700 ;
        RECT 162.960 54.745 164.155 54.905 ;
        POLYGON 164.155 54.920 164.260 54.745 164.155 54.745 ;
        POLYGON 165.765 54.920 165.845 54.920 165.845 54.760 ;
        RECT 165.845 54.760 167.865 54.920 ;
        POLYGON 165.845 54.760 165.850 54.760 165.850 54.745 ;
        RECT 165.850 54.745 167.865 54.760 ;
        RECT 162.960 54.700 164.260 54.745 ;
        POLYGON 162.960 54.700 162.985 54.700 162.985 54.665 ;
        RECT 162.985 54.665 164.260 54.700 ;
        POLYGON 162.985 54.665 162.990 54.665 162.990 54.655 ;
        RECT 162.990 54.650 164.260 54.665 ;
        RECT 161.065 54.625 161.850 54.650 ;
        POLYGON 161.850 54.650 161.865 54.625 161.850 54.625 ;
        POLYGON 162.990 54.650 162.995 54.650 162.995 54.645 ;
        RECT 162.995 54.645 164.260 54.650 ;
        POLYGON 162.995 54.645 163.005 54.645 163.005 54.625 ;
        RECT 163.005 54.625 164.260 54.645 ;
        RECT 161.065 54.595 161.865 54.625 ;
        POLYGON 161.865 54.625 161.890 54.595 161.865 54.595 ;
        POLYGON 163.005 54.625 163.025 54.625 163.025 54.595 ;
        RECT 163.025 54.595 164.260 54.625 ;
        RECT 161.065 54.570 161.890 54.595 ;
        POLYGON 161.890 54.595 161.905 54.570 161.890 54.570 ;
        POLYGON 163.025 54.595 163.040 54.595 163.040 54.570 ;
        RECT 163.040 54.570 164.260 54.595 ;
        RECT 161.065 54.510 161.905 54.570 ;
        POLYGON 161.065 54.510 161.070 54.510 161.070 54.505 ;
        RECT 161.070 54.505 161.905 54.510 ;
        RECT 159.590 54.470 160.345 54.505 ;
        RECT 158.265 54.460 158.885 54.470 ;
        RECT 151.985 54.430 157.020 54.460 ;
        POLYGON 151.940 54.430 151.940 54.425 151.935 54.425 ;
        RECT 151.940 54.425 157.020 54.430 ;
        POLYGON 157.020 54.460 157.090 54.425 157.020 54.425 ;
        POLYGON 158.265 54.460 158.310 54.460 158.310 54.425 ;
        RECT 158.310 54.445 158.885 54.460 ;
        POLYGON 158.885 54.470 158.915 54.445 158.885 54.445 ;
        POLYGON 159.590 54.470 159.615 54.470 159.615 54.445 ;
        RECT 159.615 54.445 160.345 54.470 ;
        RECT 158.310 54.425 158.915 54.445 ;
        RECT 150.105 54.420 150.605 54.425 ;
        RECT 117.275 54.375 147.585 54.420 ;
        POLYGON 147.585 54.420 147.610 54.420 147.585 54.375 ;
        POLYGON 148.525 54.420 148.525 54.375 148.495 54.375 ;
        RECT 148.525 54.375 149.250 54.420 ;
        RECT 117.275 54.345 147.570 54.375 ;
        POLYGON 147.570 54.375 147.585 54.375 147.570 54.345 ;
        POLYGON 148.495 54.375 148.495 54.345 148.475 54.345 ;
        RECT 148.495 54.345 149.250 54.375 ;
        RECT 117.275 54.310 147.550 54.345 ;
        POLYGON 147.550 54.345 147.570 54.345 147.550 54.310 ;
        POLYGON 148.475 54.345 148.475 54.310 148.455 54.310 ;
        RECT 148.475 54.310 149.250 54.345 ;
        RECT 117.275 54.260 147.505 54.310 ;
        RECT 117.250 54.225 147.505 54.260 ;
        POLYGON 147.505 54.310 147.550 54.310 147.505 54.225 ;
        POLYGON 148.455 54.310 148.455 54.235 148.405 54.235 ;
        RECT 148.455 54.290 149.250 54.310 ;
        POLYGON 149.250 54.420 149.350 54.420 149.250 54.290 ;
        POLYGON 150.055 54.420 150.055 54.415 150.050 54.415 ;
        RECT 150.055 54.415 150.605 54.420 ;
        POLYGON 150.605 54.425 150.615 54.425 150.605 54.415 ;
        POLYGON 151.935 54.425 151.935 54.415 151.920 54.415 ;
        RECT 151.935 54.420 157.090 54.425 ;
        POLYGON 157.090 54.425 157.110 54.420 157.090 54.420 ;
        POLYGON 158.310 54.425 158.315 54.425 158.315 54.420 ;
        RECT 158.315 54.420 158.915 54.425 ;
        RECT 151.935 54.415 157.110 54.420 ;
        POLYGON 150.050 54.410 150.050 54.290 149.950 54.290 ;
        RECT 150.050 54.345 150.540 54.415 ;
        POLYGON 150.540 54.415 150.605 54.415 150.540 54.345 ;
        POLYGON 151.920 54.415 151.920 54.380 151.880 54.380 ;
        RECT 151.920 54.380 157.110 54.415 ;
        POLYGON 151.880 54.380 151.880 54.375 151.875 54.375 ;
        RECT 151.880 54.375 157.110 54.380 ;
        POLYGON 157.110 54.420 157.195 54.375 157.110 54.375 ;
        POLYGON 158.315 54.420 158.380 54.420 158.380 54.375 ;
        RECT 158.380 54.415 158.915 54.420 ;
        POLYGON 158.915 54.445 158.950 54.415 158.915 54.415 ;
        POLYGON 159.615 54.445 159.645 54.445 159.645 54.415 ;
        RECT 159.645 54.440 160.345 54.445 ;
        POLYGON 160.345 54.505 160.400 54.440 160.345 54.440 ;
        POLYGON 161.070 54.505 161.080 54.505 161.080 54.495 ;
        RECT 161.080 54.495 161.905 54.505 ;
        POLYGON 161.080 54.495 161.120 54.495 161.120 54.440 ;
        RECT 161.120 54.440 161.905 54.495 ;
        RECT 159.645 54.430 160.400 54.440 ;
        POLYGON 160.400 54.440 160.410 54.430 160.400 54.430 ;
        POLYGON 161.120 54.440 161.125 54.440 161.125 54.435 ;
        RECT 161.125 54.430 161.905 54.440 ;
        RECT 159.645 54.415 160.410 54.430 ;
        RECT 158.380 54.375 158.950 54.415 ;
        POLYGON 151.875 54.375 151.875 54.345 151.835 54.345 ;
        RECT 151.875 54.370 157.195 54.375 ;
        POLYGON 157.195 54.375 157.215 54.370 157.195 54.370 ;
        POLYGON 158.380 54.375 158.385 54.375 158.385 54.370 ;
        RECT 158.385 54.370 158.950 54.375 ;
        RECT 151.875 54.345 157.215 54.370 ;
        RECT 150.050 54.290 150.485 54.345 ;
        RECT 148.455 54.235 149.170 54.290 ;
        POLYGON 148.405 54.235 148.405 54.225 148.400 54.225 ;
        RECT 148.405 54.225 149.170 54.235 ;
        RECT 51.940 54.005 111.320 54.190 ;
        POLYGON 51.940 54.005 51.955 54.005 51.955 53.955 ;
        RECT 51.955 53.955 111.320 54.005 ;
        POLYGON 51.955 53.955 53.295 53.955 53.295 50.000 ;
        RECT 53.295 53.515 111.320 53.955 ;
        POLYGON 111.320 54.190 111.390 53.515 111.320 53.515 ;
        POLYGON 117.250 54.190 117.250 53.515 117.235 53.515 ;
        RECT 117.250 54.100 147.440 54.225 ;
        POLYGON 147.440 54.225 147.505 54.225 147.440 54.100 ;
        POLYGON 148.400 54.225 148.400 54.165 148.370 54.165 ;
        RECT 148.400 54.170 149.170 54.225 ;
        POLYGON 149.170 54.290 149.250 54.290 149.170 54.170 ;
        POLYGON 149.950 54.290 149.950 54.200 149.875 54.200 ;
        RECT 149.950 54.285 150.485 54.290 ;
        POLYGON 150.485 54.345 150.540 54.345 150.485 54.285 ;
        POLYGON 151.835 54.345 151.835 54.325 151.810 54.325 ;
        RECT 151.835 54.325 157.215 54.345 ;
        POLYGON 151.810 54.325 151.810 54.285 151.765 54.285 ;
        RECT 151.810 54.285 157.215 54.325 ;
        POLYGON 157.215 54.370 157.365 54.285 157.215 54.285 ;
        POLYGON 158.385 54.370 158.495 54.370 158.495 54.285 ;
        RECT 158.495 54.325 158.950 54.370 ;
        POLYGON 158.950 54.415 159.060 54.325 158.950 54.325 ;
        POLYGON 159.645 54.415 159.700 54.415 159.700 54.360 ;
        RECT 159.700 54.360 160.410 54.415 ;
        POLYGON 159.700 54.360 159.730 54.360 159.730 54.325 ;
        RECT 159.730 54.325 160.410 54.360 ;
        RECT 158.495 54.285 159.060 54.325 ;
        RECT 149.950 54.200 150.370 54.285 ;
        POLYGON 149.875 54.200 149.875 54.170 149.855 54.170 ;
        RECT 149.875 54.170 150.370 54.200 ;
        RECT 148.400 54.165 149.155 54.170 ;
        POLYGON 148.370 54.165 148.370 54.100 148.335 54.100 ;
        RECT 148.370 54.150 149.155 54.165 ;
        POLYGON 149.155 54.170 149.170 54.170 149.155 54.150 ;
        POLYGON 149.855 54.170 149.855 54.150 149.835 54.150 ;
        RECT 149.855 54.150 150.370 54.170 ;
        POLYGON 150.370 54.285 150.485 54.285 150.370 54.150 ;
        POLYGON 151.765 54.285 151.765 54.180 151.640 54.180 ;
        RECT 151.765 54.275 157.370 54.285 ;
        POLYGON 157.370 54.285 157.380 54.275 157.370 54.275 ;
        POLYGON 158.495 54.285 158.510 54.285 158.510 54.275 ;
        RECT 151.765 54.200 157.390 54.275 ;
        POLYGON 157.390 54.275 157.515 54.200 157.390 54.200 ;
        RECT 158.510 54.270 159.060 54.285 ;
        POLYGON 158.510 54.270 158.545 54.270 158.545 54.245 ;
        RECT 158.545 54.265 159.060 54.270 ;
        POLYGON 159.060 54.325 159.125 54.265 159.060 54.265 ;
        POLYGON 159.730 54.325 159.770 54.325 159.770 54.280 ;
        RECT 159.770 54.280 160.410 54.325 ;
        POLYGON 159.770 54.280 159.780 54.280 159.780 54.265 ;
        RECT 159.780 54.275 160.410 54.280 ;
        POLYGON 160.410 54.430 160.535 54.275 160.410 54.275 ;
        POLYGON 161.125 54.430 161.190 54.430 161.190 54.350 ;
        RECT 161.190 54.350 161.905 54.430 ;
        POLYGON 161.190 54.350 161.225 54.350 161.225 54.305 ;
        RECT 161.225 54.305 161.905 54.350 ;
        POLYGON 161.225 54.305 161.240 54.305 161.240 54.280 ;
        RECT 161.240 54.275 161.905 54.305 ;
        POLYGON 161.905 54.570 162.115 54.275 161.905 54.275 ;
        POLYGON 163.040 54.570 163.115 54.570 163.115 54.445 ;
        RECT 163.115 54.565 164.260 54.570 ;
        POLYGON 164.260 54.745 164.365 54.565 164.260 54.565 ;
        POLYGON 165.850 54.745 165.930 54.745 165.930 54.565 ;
        RECT 165.930 54.740 167.865 54.745 ;
        POLYGON 167.865 54.945 167.950 54.740 167.865 54.740 ;
        POLYGON 170.630 54.945 170.710 54.945 170.710 54.745 ;
        RECT 170.710 54.740 174.925 54.945 ;
        RECT 165.930 54.565 167.950 54.740 ;
        RECT 163.115 54.535 164.365 54.565 ;
        POLYGON 164.365 54.565 164.385 54.535 164.365 54.535 ;
        POLYGON 165.930 54.565 165.940 54.565 165.940 54.545 ;
        RECT 165.940 54.550 167.950 54.565 ;
        POLYGON 167.950 54.740 168.030 54.550 167.950 54.550 ;
        POLYGON 170.710 54.740 170.750 54.740 170.750 54.640 ;
        RECT 170.750 54.640 174.925 54.740 ;
        POLYGON 170.750 54.640 170.775 54.640 170.775 54.560 ;
        RECT 170.775 54.570 174.925 54.640 ;
        POLYGON 174.925 55.060 175.105 54.570 174.925 54.570 ;
        POLYGON 181.875 55.060 182.015 55.060 182.015 54.575 ;
        RECT 182.015 54.570 196.025 55.060 ;
        RECT 170.775 54.555 175.105 54.570 ;
        POLYGON 175.105 54.570 175.110 54.555 175.105 54.555 ;
        POLYGON 182.015 54.570 182.020 54.570 182.020 54.555 ;
        RECT 182.020 54.555 196.025 54.570 ;
        RECT 170.775 54.550 175.110 54.555 ;
        RECT 165.940 54.535 168.030 54.550 ;
        RECT 163.115 54.445 164.385 54.535 ;
        POLYGON 163.115 54.445 163.120 54.445 163.120 54.440 ;
        RECT 163.120 54.440 164.385 54.445 ;
        POLYGON 163.120 54.440 163.145 54.440 163.145 54.400 ;
        RECT 163.145 54.435 164.385 54.440 ;
        POLYGON 164.385 54.535 164.435 54.435 164.385 54.435 ;
        POLYGON 165.940 54.535 165.990 54.535 165.990 54.435 ;
        RECT 165.990 54.505 168.030 54.535 ;
        POLYGON 168.030 54.550 168.050 54.505 168.030 54.505 ;
        POLYGON 170.775 54.550 170.790 54.550 170.790 54.515 ;
        RECT 170.790 54.505 175.110 54.550 ;
        RECT 165.990 54.435 168.050 54.505 ;
        RECT 163.145 54.400 164.435 54.435 ;
        POLYGON 163.145 54.400 163.215 54.400 163.215 54.280 ;
        RECT 163.215 54.330 164.435 54.400 ;
        POLYGON 164.435 54.435 164.495 54.330 164.435 54.330 ;
        POLYGON 165.990 54.435 166.015 54.435 166.015 54.380 ;
        RECT 166.015 54.380 168.050 54.435 ;
        POLYGON 166.015 54.380 166.030 54.380 166.030 54.340 ;
        RECT 166.030 54.330 168.050 54.380 ;
        RECT 163.215 54.275 164.495 54.330 ;
        RECT 159.780 54.265 160.535 54.275 ;
        POLYGON 160.535 54.275 160.540 54.265 160.535 54.265 ;
        POLYGON 161.240 54.275 161.250 54.275 161.250 54.265 ;
        RECT 161.250 54.265 162.115 54.275 ;
        RECT 158.545 54.260 159.125 54.265 ;
        POLYGON 159.125 54.265 159.130 54.260 159.125 54.260 ;
        POLYGON 159.780 54.265 159.785 54.265 159.785 54.260 ;
        RECT 159.785 54.260 160.540 54.265 ;
        RECT 158.545 54.245 159.130 54.260 ;
        POLYGON 158.545 54.245 158.595 54.245 158.595 54.200 ;
        RECT 158.595 54.215 159.130 54.245 ;
        POLYGON 159.130 54.260 159.180 54.215 159.130 54.215 ;
        POLYGON 159.785 54.260 159.795 54.260 159.795 54.250 ;
        RECT 159.795 54.250 160.540 54.260 ;
        POLYGON 159.800 54.250 159.830 54.250 159.830 54.215 ;
        RECT 159.830 54.215 160.540 54.250 ;
        RECT 158.595 54.200 159.180 54.215 ;
        RECT 151.765 54.180 157.515 54.200 ;
        POLYGON 157.515 54.200 157.545 54.180 157.515 54.180 ;
        POLYGON 158.595 54.200 158.620 54.200 158.620 54.180 ;
        RECT 158.620 54.180 159.180 54.200 ;
        POLYGON 151.640 54.180 151.640 54.175 151.630 54.175 ;
        RECT 151.640 54.175 157.545 54.180 ;
        POLYGON 151.630 54.175 151.630 54.150 151.605 54.150 ;
        RECT 151.630 54.150 157.545 54.175 ;
        RECT 148.370 54.100 149.115 54.150 ;
        RECT 117.250 54.050 147.415 54.100 ;
        POLYGON 147.415 54.100 147.440 54.100 147.415 54.050 ;
        POLYGON 148.335 54.100 148.335 54.050 148.305 54.050 ;
        RECT 148.335 54.090 149.115 54.100 ;
        POLYGON 149.115 54.150 149.155 54.150 149.115 54.090 ;
        POLYGON 149.835 54.145 149.835 54.100 149.795 54.100 ;
        RECT 149.835 54.125 150.350 54.150 ;
        POLYGON 150.350 54.150 150.370 54.150 150.350 54.125 ;
        POLYGON 151.605 54.150 151.605 54.125 151.580 54.125 ;
        RECT 151.605 54.125 157.545 54.150 ;
        RECT 149.835 54.115 150.340 54.125 ;
        POLYGON 150.340 54.125 150.350 54.125 150.340 54.115 ;
        POLYGON 151.580 54.125 151.580 54.115 151.570 54.115 ;
        RECT 151.580 54.115 157.545 54.125 ;
        RECT 149.835 54.100 150.325 54.115 ;
        POLYGON 149.795 54.100 149.795 54.095 149.790 54.095 ;
        RECT 149.795 54.095 150.325 54.100 ;
        RECT 149.790 54.090 150.325 54.095 ;
        POLYGON 150.325 54.115 150.340 54.115 150.325 54.090 ;
        POLYGON 151.570 54.115 151.570 54.090 151.540 54.090 ;
        RECT 151.570 54.105 157.545 54.115 ;
        POLYGON 157.545 54.180 157.665 54.105 157.545 54.105 ;
        POLYGON 158.620 54.180 158.630 54.180 158.630 54.175 ;
        RECT 158.630 54.175 159.180 54.180 ;
        POLYGON 158.630 54.175 158.705 54.175 158.705 54.105 ;
        RECT 158.705 54.110 159.180 54.175 ;
        POLYGON 159.180 54.215 159.300 54.110 159.180 54.110 ;
        POLYGON 159.830 54.215 159.910 54.215 159.910 54.125 ;
        RECT 159.910 54.210 160.540 54.215 ;
        POLYGON 160.540 54.265 160.585 54.210 160.540 54.210 ;
        POLYGON 161.250 54.265 161.260 54.265 161.260 54.255 ;
        RECT 161.260 54.255 162.115 54.265 ;
        POLYGON 161.260 54.255 161.290 54.255 161.290 54.210 ;
        RECT 161.290 54.210 162.115 54.255 ;
        RECT 159.910 54.135 160.585 54.210 ;
        POLYGON 160.585 54.210 160.640 54.135 160.585 54.135 ;
        POLYGON 161.290 54.210 161.325 54.210 161.325 54.160 ;
        RECT 161.325 54.190 162.115 54.210 ;
        POLYGON 162.115 54.275 162.170 54.190 162.115 54.190 ;
        POLYGON 163.215 54.275 163.245 54.275 163.245 54.220 ;
        RECT 163.245 54.220 164.495 54.275 ;
        POLYGON 163.245 54.220 163.260 54.220 163.260 54.190 ;
        RECT 163.260 54.190 164.495 54.220 ;
        RECT 161.325 54.180 162.170 54.190 ;
        POLYGON 162.170 54.190 162.175 54.180 162.170 54.180 ;
        POLYGON 163.260 54.190 163.265 54.190 163.265 54.180 ;
        RECT 163.265 54.180 164.495 54.190 ;
        RECT 161.325 54.160 162.175 54.180 ;
        POLYGON 161.325 54.160 161.340 54.160 161.340 54.135 ;
        RECT 161.340 54.135 162.175 54.160 ;
        RECT 159.910 54.125 160.640 54.135 ;
        POLYGON 159.910 54.125 159.925 54.125 159.925 54.110 ;
        RECT 159.925 54.110 160.640 54.125 ;
        RECT 158.705 54.105 159.300 54.110 ;
        RECT 151.570 54.095 157.665 54.105 ;
        POLYGON 157.665 54.105 157.685 54.095 157.665 54.095 ;
        POLYGON 158.705 54.105 158.720 54.105 158.720 54.095 ;
        RECT 158.720 54.095 159.300 54.105 ;
        RECT 151.570 54.090 157.685 54.095 ;
        RECT 148.335 54.050 148.985 54.090 ;
        RECT 117.250 53.990 147.390 54.050 ;
        POLYGON 147.390 54.050 147.415 54.050 147.390 53.990 ;
        POLYGON 148.305 54.045 148.305 53.990 148.275 53.990 ;
        RECT 148.305 53.990 148.985 54.050 ;
        RECT 117.250 53.905 147.350 53.990 ;
        POLYGON 147.350 53.990 147.390 53.990 147.350 53.905 ;
        POLYGON 148.275 53.990 148.275 53.910 148.230 53.910 ;
        RECT 148.275 53.910 148.985 53.990 ;
        RECT 117.250 53.845 147.320 53.905 ;
        POLYGON 147.320 53.905 147.350 53.905 147.320 53.845 ;
        POLYGON 148.230 53.905 148.230 53.845 148.195 53.845 ;
        RECT 148.230 53.885 148.985 53.910 ;
        POLYGON 148.985 54.090 149.115 54.090 148.985 53.885 ;
        POLYGON 149.790 54.090 149.790 53.975 149.710 53.975 ;
        RECT 149.790 54.015 150.265 54.090 ;
        POLYGON 150.265 54.090 150.325 54.090 150.265 54.015 ;
        POLYGON 151.540 54.090 151.540 54.030 151.475 54.030 ;
        RECT 151.540 54.070 157.685 54.090 ;
        POLYGON 157.685 54.095 157.715 54.070 157.685 54.070 ;
        POLYGON 158.720 54.095 158.745 54.095 158.745 54.070 ;
        RECT 158.745 54.090 159.300 54.095 ;
        POLYGON 159.300 54.110 159.320 54.090 159.300 54.090 ;
        POLYGON 159.925 54.110 159.945 54.110 159.945 54.090 ;
        RECT 159.945 54.090 160.640 54.110 ;
        RECT 158.745 54.070 159.320 54.090 ;
        RECT 151.540 54.030 157.715 54.070 ;
        POLYGON 151.475 54.030 151.475 54.025 151.465 54.025 ;
        RECT 151.475 54.025 157.715 54.030 ;
        POLYGON 151.465 54.025 151.465 54.015 151.455 54.015 ;
        RECT 151.465 54.015 157.715 54.025 ;
        RECT 149.790 53.975 150.175 54.015 ;
        POLYGON 149.710 53.975 149.710 53.885 149.645 53.885 ;
        RECT 149.710 53.900 150.175 53.975 ;
        POLYGON 150.175 54.015 150.265 54.015 150.175 53.900 ;
        POLYGON 151.455 54.015 151.455 53.900 151.340 53.900 ;
        RECT 151.455 54.005 157.715 54.015 ;
        POLYGON 157.715 54.070 157.815 54.005 157.715 54.005 ;
        POLYGON 158.745 54.070 158.760 54.070 158.760 54.060 ;
        RECT 158.760 54.060 159.320 54.070 ;
        POLYGON 158.760 54.060 158.790 54.060 158.790 54.035 ;
        RECT 158.790 54.050 159.320 54.060 ;
        POLYGON 159.320 54.090 159.355 54.050 159.320 54.050 ;
        POLYGON 159.945 54.090 159.960 54.090 159.960 54.075 ;
        RECT 159.960 54.075 160.640 54.090 ;
        POLYGON 159.960 54.075 159.975 54.075 159.975 54.055 ;
        RECT 159.975 54.050 160.640 54.075 ;
        RECT 158.790 54.035 159.355 54.050 ;
        POLYGON 158.790 54.035 158.815 54.035 158.815 54.015 ;
        RECT 158.815 54.015 159.355 54.035 ;
        POLYGON 158.815 54.015 158.825 54.015 158.825 54.005 ;
        RECT 158.825 54.005 159.355 54.015 ;
        RECT 151.455 53.955 157.815 54.005 ;
        POLYGON 157.815 54.005 157.885 53.955 157.815 53.955 ;
        POLYGON 158.825 54.005 158.875 54.005 158.875 53.955 ;
        RECT 158.875 53.970 159.355 54.005 ;
        POLYGON 159.355 54.050 159.440 53.970 159.355 53.970 ;
        POLYGON 159.975 54.050 160.005 54.050 160.005 54.015 ;
        RECT 160.005 54.040 160.640 54.050 ;
        POLYGON 160.640 54.135 160.710 54.040 160.640 54.040 ;
        POLYGON 161.340 54.135 161.360 54.135 161.360 54.110 ;
        RECT 161.360 54.125 162.175 54.135 ;
        POLYGON 162.175 54.180 162.210 54.125 162.175 54.125 ;
        POLYGON 163.265 54.180 163.270 54.180 163.270 54.175 ;
        RECT 163.270 54.175 164.495 54.180 ;
        POLYGON 163.270 54.175 163.295 54.175 163.295 54.125 ;
        RECT 163.295 54.145 164.495 54.175 ;
        POLYGON 164.495 54.330 164.595 54.145 164.495 54.145 ;
        POLYGON 166.030 54.330 166.095 54.330 166.095 54.170 ;
        RECT 166.095 54.170 168.050 54.330 ;
        POLYGON 166.095 54.170 166.105 54.170 166.105 54.145 ;
        RECT 166.105 54.145 168.050 54.170 ;
        RECT 163.295 54.125 164.595 54.145 ;
        RECT 161.360 54.110 162.210 54.125 ;
        POLYGON 161.360 54.110 161.410 54.110 161.410 54.040 ;
        RECT 161.410 54.040 162.210 54.110 ;
        RECT 160.005 54.015 160.710 54.040 ;
        POLYGON 160.005 54.015 160.010 54.015 160.010 54.010 ;
        RECT 160.010 54.010 160.710 54.015 ;
        POLYGON 160.010 54.010 160.045 54.010 160.045 53.970 ;
        RECT 160.045 53.975 160.710 54.010 ;
        POLYGON 160.710 54.040 160.760 53.975 160.710 53.975 ;
        POLYGON 161.410 54.040 161.445 54.040 161.445 53.995 ;
        RECT 161.445 53.995 162.210 54.040 ;
        POLYGON 161.445 53.995 161.455 53.995 161.455 53.980 ;
        RECT 161.455 53.975 162.210 53.995 ;
        RECT 160.045 53.970 160.760 53.975 ;
        RECT 158.875 53.955 159.440 53.970 ;
        RECT 151.455 53.910 157.885 53.955 ;
        POLYGON 157.885 53.955 157.945 53.910 157.885 53.910 ;
        POLYGON 158.875 53.955 158.925 53.955 158.925 53.910 ;
        RECT 158.925 53.910 159.440 53.955 ;
        RECT 151.455 53.900 157.945 53.910 ;
        POLYGON 157.945 53.910 157.960 53.900 157.945 53.900 ;
        POLYGON 158.925 53.910 158.935 53.910 158.935 53.900 ;
        RECT 158.935 53.900 159.440 53.910 ;
        RECT 149.710 53.885 150.165 53.900 ;
        POLYGON 150.165 53.900 150.175 53.900 150.165 53.885 ;
        POLYGON 151.340 53.900 151.340 53.885 151.325 53.885 ;
        RECT 151.340 53.885 157.960 53.900 ;
        POLYGON 157.960 53.900 157.980 53.885 157.960 53.885 ;
        POLYGON 158.935 53.900 158.950 53.900 158.950 53.885 ;
        RECT 158.950 53.885 159.440 53.900 ;
        RECT 148.230 53.880 148.980 53.885 ;
        POLYGON 148.980 53.885 148.985 53.885 148.980 53.880 ;
        POLYGON 149.645 53.885 149.645 53.880 149.640 53.880 ;
        RECT 149.645 53.880 150.075 53.885 ;
        RECT 148.230 53.850 148.965 53.880 ;
        POLYGON 148.965 53.880 148.980 53.880 148.965 53.850 ;
        POLYGON 149.640 53.880 149.640 53.850 149.615 53.850 ;
        RECT 149.640 53.850 150.075 53.880 ;
        RECT 148.230 53.845 148.930 53.850 ;
        RECT 117.250 53.815 147.310 53.845 ;
        POLYGON 147.310 53.845 147.320 53.845 147.310 53.815 ;
        POLYGON 148.195 53.845 148.195 53.820 148.180 53.820 ;
        RECT 148.195 53.820 148.930 53.845 ;
        RECT 117.250 53.805 147.305 53.815 ;
        POLYGON 148.180 53.815 148.180 53.810 148.175 53.810 ;
        RECT 148.180 53.810 148.930 53.820 ;
        RECT 117.250 53.760 147.285 53.805 ;
        POLYGON 147.285 53.805 147.305 53.805 147.285 53.760 ;
        POLYGON 148.175 53.810 148.175 53.765 148.155 53.765 ;
        RECT 148.175 53.795 148.930 53.810 ;
        POLYGON 148.930 53.850 148.965 53.850 148.930 53.795 ;
        POLYGON 149.615 53.845 149.615 53.840 149.610 53.840 ;
        RECT 149.615 53.840 150.075 53.850 ;
        POLYGON 149.610 53.840 149.610 53.795 149.580 53.795 ;
        RECT 149.610 53.795 150.075 53.840 ;
        RECT 148.175 53.765 148.860 53.795 ;
        RECT 117.250 53.660 147.240 53.760 ;
        POLYGON 147.240 53.760 147.285 53.760 147.240 53.660 ;
        POLYGON 148.155 53.760 148.155 53.660 148.105 53.660 ;
        RECT 148.155 53.675 148.860 53.765 ;
        POLYGON 148.860 53.795 148.930 53.795 148.860 53.675 ;
        POLYGON 149.580 53.795 149.580 53.775 149.565 53.775 ;
        RECT 149.580 53.775 150.075 53.795 ;
        POLYGON 149.565 53.775 149.565 53.750 149.550 53.750 ;
        RECT 149.565 53.755 150.075 53.775 ;
        POLYGON 150.075 53.885 150.165 53.885 150.075 53.755 ;
        POLYGON 151.325 53.885 151.325 53.875 151.315 53.875 ;
        RECT 151.325 53.875 157.980 53.885 ;
        POLYGON 151.310 53.875 151.310 53.805 151.245 53.805 ;
        RECT 151.310 53.825 157.980 53.875 ;
        POLYGON 157.980 53.885 158.050 53.825 157.980 53.825 ;
        POLYGON 158.950 53.885 158.995 53.885 158.995 53.845 ;
        RECT 158.995 53.845 159.440 53.885 ;
        POLYGON 158.995 53.845 159.015 53.845 159.015 53.825 ;
        RECT 159.015 53.830 159.440 53.845 ;
        POLYGON 159.440 53.970 159.580 53.830 159.440 53.830 ;
        POLYGON 160.045 53.970 160.155 53.970 160.155 53.835 ;
        RECT 160.155 53.835 160.760 53.970 ;
        POLYGON 160.155 53.835 160.160 53.835 160.160 53.830 ;
        RECT 160.160 53.830 160.760 53.835 ;
        POLYGON 160.760 53.975 160.860 53.830 160.760 53.830 ;
        POLYGON 161.455 53.975 161.490 53.975 161.490 53.925 ;
        RECT 161.490 53.925 162.210 53.975 ;
        POLYGON 161.490 53.925 161.545 53.925 161.545 53.835 ;
        RECT 161.545 53.890 162.210 53.925 ;
        POLYGON 162.210 54.125 162.365 53.890 162.210 53.890 ;
        POLYGON 163.295 54.125 163.350 54.125 163.350 54.020 ;
        RECT 163.350 54.100 164.595 54.125 ;
        POLYGON 164.595 54.145 164.615 54.100 164.595 54.100 ;
        POLYGON 166.105 54.145 166.120 54.145 166.120 54.105 ;
        RECT 166.120 54.100 168.050 54.145 ;
        POLYGON 168.050 54.505 168.205 54.100 168.050 54.100 ;
        POLYGON 170.790 54.505 170.925 54.505 170.925 54.110 ;
        RECT 170.925 54.100 175.110 54.505 ;
        RECT 163.350 54.020 164.615 54.100 ;
        POLYGON 163.350 54.020 163.370 54.020 163.370 53.980 ;
        RECT 163.370 53.980 164.615 54.020 ;
        POLYGON 163.370 53.980 163.395 53.980 163.395 53.935 ;
        RECT 163.395 53.945 164.615 53.980 ;
        POLYGON 164.615 54.100 164.690 53.945 164.615 53.945 ;
        POLYGON 166.120 54.100 166.165 54.100 166.165 54.000 ;
        RECT 166.165 54.015 168.205 54.100 ;
        POLYGON 168.205 54.100 168.240 54.015 168.205 54.015 ;
        POLYGON 170.925 54.100 170.955 54.100 170.955 54.020 ;
        RECT 170.955 54.015 175.110 54.100 ;
        RECT 166.165 54.000 168.240 54.015 ;
        POLYGON 166.165 54.000 166.180 54.000 166.180 53.955 ;
        RECT 166.180 53.945 168.240 54.000 ;
        RECT 163.395 53.935 164.690 53.945 ;
        POLYGON 163.395 53.935 163.415 53.935 163.415 53.895 ;
        RECT 163.415 53.915 164.690 53.935 ;
        POLYGON 164.690 53.945 164.705 53.915 164.690 53.915 ;
        POLYGON 166.180 53.945 166.190 53.945 166.190 53.925 ;
        RECT 166.190 53.915 168.240 53.945 ;
        RECT 163.415 53.890 164.705 53.915 ;
        RECT 161.545 53.830 162.365 53.890 ;
        RECT 159.015 53.825 159.580 53.830 ;
        RECT 151.310 53.805 158.050 53.825 ;
        POLYGON 151.245 53.805 151.245 53.755 151.200 53.755 ;
        RECT 151.245 53.755 158.050 53.805 ;
        RECT 149.565 53.750 150.050 53.755 ;
        POLYGON 149.550 53.750 149.550 53.720 149.525 53.720 ;
        RECT 149.550 53.720 150.050 53.750 ;
        POLYGON 150.050 53.755 150.075 53.755 150.050 53.720 ;
        POLYGON 151.200 53.755 151.200 53.720 151.165 53.720 ;
        RECT 151.200 53.720 158.050 53.755 ;
        POLYGON 149.525 53.720 149.525 53.675 149.495 53.675 ;
        RECT 149.525 53.675 150.010 53.720 ;
        RECT 148.155 53.660 148.770 53.675 ;
        RECT 117.250 53.580 147.210 53.660 ;
        POLYGON 147.210 53.660 147.240 53.660 147.210 53.580 ;
        POLYGON 148.105 53.660 148.105 53.580 148.065 53.580 ;
        RECT 148.105 53.580 148.770 53.660 ;
        RECT 117.250 53.560 147.200 53.580 ;
        POLYGON 147.200 53.580 147.210 53.580 147.200 53.560 ;
        POLYGON 148.065 53.580 148.065 53.560 148.055 53.560 ;
        RECT 148.065 53.560 148.770 53.580 ;
        RECT 117.250 53.535 147.195 53.560 ;
        POLYGON 147.195 53.560 147.200 53.560 147.195 53.545 ;
        POLYGON 147.195 53.545 147.200 53.535 147.195 53.535 ;
        RECT 117.250 53.520 147.200 53.535 ;
        POLYGON 148.055 53.560 148.055 53.530 148.040 53.530 ;
        RECT 148.055 53.530 148.770 53.560 ;
        POLYGON 147.200 53.525 147.205 53.520 147.200 53.520 ;
        RECT 117.250 53.515 147.205 53.520 ;
        RECT 53.295 52.805 111.390 53.515 ;
        POLYGON 111.390 53.515 111.460 52.805 111.390 52.805 ;
        RECT 117.235 53.500 147.205 53.515 ;
        POLYGON 148.040 53.525 148.040 53.510 148.030 53.510 ;
        RECT 148.040 53.510 148.770 53.530 ;
        POLYGON 148.770 53.675 148.860 53.675 148.770 53.510 ;
        POLYGON 149.495 53.670 149.495 53.510 149.395 53.510 ;
        RECT 149.495 53.660 150.010 53.675 ;
        POLYGON 150.010 53.720 150.050 53.720 150.010 53.660 ;
        POLYGON 151.165 53.720 151.165 53.715 151.160 53.715 ;
        RECT 151.165 53.715 158.050 53.720 ;
        POLYGON 151.160 53.715 151.160 53.660 151.115 53.660 ;
        RECT 151.160 53.695 158.050 53.715 ;
        POLYGON 158.050 53.825 158.215 53.695 158.050 53.695 ;
        POLYGON 159.015 53.825 159.060 53.825 159.060 53.785 ;
        RECT 159.060 53.785 159.580 53.825 ;
        POLYGON 159.580 53.830 159.620 53.785 159.580 53.785 ;
        POLYGON 160.160 53.830 160.165 53.830 160.165 53.825 ;
        RECT 160.165 53.825 160.860 53.830 ;
        POLYGON 160.165 53.825 160.190 53.825 160.190 53.790 ;
        RECT 160.190 53.795 160.860 53.825 ;
        POLYGON 160.860 53.830 160.880 53.795 160.860 53.795 ;
        POLYGON 161.545 53.830 161.555 53.830 161.555 53.820 ;
        RECT 161.555 53.820 162.365 53.830 ;
        POLYGON 161.555 53.820 161.570 53.820 161.570 53.795 ;
        RECT 161.570 53.800 162.365 53.820 ;
        POLYGON 162.365 53.890 162.410 53.800 162.365 53.800 ;
        POLYGON 163.415 53.890 163.420 53.890 163.420 53.885 ;
        RECT 163.420 53.885 164.705 53.890 ;
        POLYGON 163.420 53.885 163.450 53.885 163.450 53.825 ;
        RECT 163.450 53.825 164.705 53.885 ;
        POLYGON 163.450 53.825 163.460 53.825 163.460 53.800 ;
        RECT 163.460 53.800 164.705 53.825 ;
        RECT 161.570 53.795 162.410 53.800 ;
        RECT 160.190 53.785 160.880 53.795 ;
        POLYGON 159.060 53.785 159.070 53.785 159.070 53.775 ;
        RECT 159.070 53.775 159.620 53.785 ;
        POLYGON 159.070 53.775 159.140 53.775 159.140 53.695 ;
        RECT 159.140 53.700 159.620 53.775 ;
        POLYGON 159.620 53.785 159.700 53.700 159.620 53.700 ;
        POLYGON 160.190 53.785 160.205 53.785 160.205 53.770 ;
        RECT 160.205 53.770 160.880 53.785 ;
        POLYGON 160.205 53.770 160.260 53.770 160.260 53.700 ;
        RECT 160.260 53.760 160.880 53.770 ;
        POLYGON 160.880 53.795 160.905 53.760 160.880 53.760 ;
        POLYGON 161.570 53.795 161.590 53.795 161.590 53.760 ;
        RECT 161.590 53.760 162.410 53.795 ;
        RECT 160.260 53.730 160.905 53.760 ;
        POLYGON 160.905 53.760 160.925 53.730 160.905 53.730 ;
        POLYGON 161.590 53.760 161.605 53.760 161.605 53.740 ;
        RECT 161.605 53.740 162.410 53.760 ;
        POLYGON 161.605 53.740 161.610 53.740 161.610 53.730 ;
        RECT 161.610 53.730 162.410 53.740 ;
        RECT 160.260 53.700 160.925 53.730 ;
        RECT 159.140 53.695 159.700 53.700 ;
        RECT 151.160 53.685 158.215 53.695 ;
        POLYGON 158.215 53.695 158.230 53.685 158.215 53.685 ;
        POLYGON 159.140 53.695 159.150 53.695 159.150 53.685 ;
        RECT 159.150 53.685 159.700 53.695 ;
        RECT 151.160 53.675 158.230 53.685 ;
        POLYGON 158.230 53.685 158.240 53.675 158.230 53.675 ;
        POLYGON 159.150 53.685 159.160 53.685 159.160 53.675 ;
        RECT 159.160 53.675 159.700 53.685 ;
        RECT 151.160 53.660 158.240 53.675 ;
        RECT 149.495 53.630 149.995 53.660 ;
        POLYGON 149.995 53.660 150.010 53.660 149.995 53.630 ;
        POLYGON 151.115 53.660 151.115 53.635 151.090 53.635 ;
        RECT 151.115 53.655 158.240 53.660 ;
        POLYGON 158.240 53.675 158.265 53.655 158.240 53.655 ;
        POLYGON 159.160 53.675 159.180 53.675 159.180 53.655 ;
        RECT 159.180 53.655 159.700 53.675 ;
        RECT 151.115 53.635 158.265 53.655 ;
        RECT 149.495 53.515 149.920 53.630 ;
        POLYGON 149.920 53.630 149.995 53.630 149.920 53.515 ;
        POLYGON 151.090 53.630 151.090 53.615 151.075 53.615 ;
        RECT 151.090 53.615 158.265 53.635 ;
        POLYGON 151.075 53.615 151.075 53.545 151.010 53.545 ;
        RECT 151.075 53.550 158.265 53.615 ;
        POLYGON 158.265 53.655 158.380 53.550 158.265 53.550 ;
        POLYGON 159.180 53.655 159.250 53.655 159.250 53.585 ;
        RECT 159.250 53.625 159.700 53.655 ;
        POLYGON 159.700 53.700 159.770 53.625 159.700 53.625 ;
        POLYGON 160.260 53.700 160.280 53.700 160.280 53.675 ;
        RECT 160.280 53.675 160.925 53.700 ;
        POLYGON 160.280 53.675 160.295 53.675 160.295 53.655 ;
        RECT 160.295 53.655 160.925 53.675 ;
        POLYGON 160.295 53.655 160.315 53.655 160.315 53.625 ;
        RECT 160.315 53.625 160.925 53.655 ;
        RECT 159.250 53.595 159.770 53.625 ;
        POLYGON 159.770 53.625 159.795 53.595 159.770 53.595 ;
        POLYGON 160.315 53.625 160.340 53.625 160.340 53.595 ;
        RECT 160.340 53.595 160.925 53.625 ;
        RECT 159.250 53.585 159.800 53.595 ;
        POLYGON 159.250 53.585 159.275 53.585 159.275 53.555 ;
        RECT 159.275 53.550 159.800 53.585 ;
        RECT 151.075 53.545 158.380 53.550 ;
        POLYGON 151.010 53.545 151.010 53.515 150.985 53.515 ;
        RECT 151.010 53.515 158.380 53.545 ;
        RECT 149.495 53.510 149.860 53.515 ;
        POLYGON 147.205 53.510 147.210 53.500 147.205 53.500 ;
        POLYGON 148.030 53.510 148.030 53.500 148.025 53.500 ;
        RECT 148.030 53.500 148.745 53.510 ;
        POLYGON 117.235 53.460 117.235 52.930 117.225 52.930 ;
        RECT 117.235 53.310 147.210 53.500 ;
        POLYGON 147.210 53.500 147.270 53.310 147.210 53.310 ;
        RECT 117.235 53.295 147.270 53.310 ;
        POLYGON 148.025 53.500 148.025 53.300 147.940 53.300 ;
        RECT 148.025 53.465 148.745 53.500 ;
        POLYGON 148.745 53.510 148.770 53.510 148.745 53.465 ;
        POLYGON 149.395 53.510 149.395 53.495 149.385 53.495 ;
        RECT 149.395 53.495 149.860 53.510 ;
        POLYGON 149.385 53.495 149.385 53.470 149.370 53.470 ;
        RECT 149.385 53.470 149.860 53.495 ;
        RECT 148.025 53.375 148.700 53.465 ;
        POLYGON 148.700 53.465 148.745 53.465 148.700 53.375 ;
        POLYGON 149.370 53.465 149.370 53.435 149.350 53.435 ;
        RECT 149.370 53.435 149.860 53.470 ;
        POLYGON 149.350 53.435 149.350 53.375 149.315 53.375 ;
        RECT 149.350 53.415 149.860 53.435 ;
        POLYGON 149.860 53.515 149.920 53.515 149.860 53.415 ;
        POLYGON 150.985 53.515 150.985 53.465 150.945 53.465 ;
        RECT 150.985 53.465 158.380 53.515 ;
        POLYGON 150.945 53.465 150.945 53.440 150.920 53.440 ;
        RECT 150.945 53.440 158.380 53.465 ;
        POLYGON 150.920 53.440 150.920 53.415 150.900 53.415 ;
        RECT 150.920 53.435 158.380 53.440 ;
        POLYGON 158.380 53.550 158.510 53.435 158.380 53.435 ;
        POLYGON 159.275 53.550 159.305 53.550 159.305 53.520 ;
        RECT 159.305 53.520 159.800 53.550 ;
        POLYGON 159.310 53.520 159.320 53.520 159.320 53.510 ;
        RECT 159.320 53.510 159.800 53.520 ;
        RECT 150.920 53.415 158.510 53.435 ;
        POLYGON 159.320 53.510 159.380 53.510 159.380 53.430 ;
        RECT 159.380 53.455 159.800 53.510 ;
        POLYGON 159.800 53.595 159.910 53.455 159.800 53.455 ;
        POLYGON 160.340 53.595 160.380 53.595 160.380 53.540 ;
        RECT 160.380 53.540 160.925 53.595 ;
        POLYGON 160.925 53.730 161.040 53.540 160.925 53.540 ;
        POLYGON 161.610 53.730 161.615 53.730 161.615 53.725 ;
        RECT 161.615 53.725 162.410 53.730 ;
        POLYGON 161.615 53.725 161.675 53.725 161.675 53.620 ;
        RECT 161.675 53.705 162.410 53.725 ;
        POLYGON 162.410 53.800 162.465 53.705 162.410 53.705 ;
        POLYGON 163.460 53.800 163.495 53.800 163.495 53.725 ;
        RECT 163.495 53.735 164.705 53.800 ;
        POLYGON 164.705 53.915 164.785 53.735 164.705 53.735 ;
        POLYGON 166.190 53.915 166.255 53.915 166.255 53.740 ;
        RECT 166.255 53.770 168.240 53.915 ;
        POLYGON 168.240 54.015 168.325 53.770 168.240 53.770 ;
        POLYGON 170.955 54.015 170.980 54.015 170.980 53.945 ;
        RECT 170.980 53.950 175.110 54.015 ;
        POLYGON 175.110 54.555 175.305 53.950 175.110 53.950 ;
        POLYGON 182.020 54.555 182.060 54.555 182.060 54.420 ;
        RECT 182.060 54.420 196.025 54.555 ;
        POLYGON 182.060 54.420 182.165 54.420 182.165 53.960 ;
        RECT 182.165 54.135 196.025 54.420 ;
        POLYGON 196.025 55.640 196.465 54.135 196.025 54.135 ;
        POLYGON 206.270 55.640 206.275 55.640 206.275 55.605 ;
        RECT 206.275 55.605 222.225 55.640 ;
        POLYGON 206.275 55.605 206.370 55.605 206.370 54.185 ;
        RECT 206.370 54.185 222.225 55.605 ;
        POLYGON 206.370 54.185 206.375 54.185 206.375 54.135 ;
        RECT 182.165 54.130 196.465 54.135 ;
        POLYGON 196.465 54.135 196.470 54.130 196.465 54.130 ;
        RECT 206.375 54.130 222.225 54.185 ;
        RECT 182.165 53.950 196.470 54.130 ;
        RECT 170.980 53.945 175.305 53.950 ;
        POLYGON 170.980 53.945 171.025 53.945 171.025 53.785 ;
        RECT 171.025 53.900 175.305 53.945 ;
        POLYGON 175.305 53.950 175.315 53.900 175.305 53.900 ;
        POLYGON 182.165 53.950 182.175 53.950 182.175 53.915 ;
        RECT 182.175 53.900 196.470 53.950 ;
        RECT 171.025 53.770 175.315 53.900 ;
        RECT 166.255 53.735 168.325 53.770 ;
        RECT 163.495 53.725 164.785 53.735 ;
        POLYGON 163.495 53.725 163.505 53.725 163.505 53.705 ;
        RECT 163.505 53.705 164.785 53.725 ;
        RECT 161.675 53.620 162.465 53.705 ;
        POLYGON 161.675 53.620 161.710 53.620 161.710 53.560 ;
        RECT 161.710 53.605 162.465 53.620 ;
        POLYGON 162.465 53.705 162.525 53.605 162.465 53.605 ;
        POLYGON 163.505 53.705 163.540 53.705 163.540 53.635 ;
        RECT 163.540 53.635 164.785 53.705 ;
        POLYGON 163.540 53.635 163.545 53.635 163.545 53.615 ;
        RECT 163.545 53.615 164.785 53.635 ;
        POLYGON 163.545 53.615 163.550 53.615 163.550 53.605 ;
        RECT 163.550 53.605 164.785 53.615 ;
        RECT 161.710 53.560 162.525 53.605 ;
        POLYGON 161.710 53.560 161.720 53.560 161.720 53.540 ;
        RECT 161.720 53.540 162.525 53.560 ;
        POLYGON 160.380 53.540 160.385 53.540 160.385 53.535 ;
        RECT 160.385 53.535 161.040 53.540 ;
        POLYGON 160.385 53.535 160.400 53.535 160.400 53.510 ;
        RECT 160.400 53.510 161.040 53.535 ;
        POLYGON 160.400 53.510 160.440 53.510 160.440 53.455 ;
        RECT 160.440 53.500 161.040 53.510 ;
        POLYGON 161.040 53.540 161.065 53.500 161.040 53.500 ;
        POLYGON 161.720 53.540 161.740 53.540 161.740 53.505 ;
        RECT 161.740 53.500 162.525 53.540 ;
        RECT 160.440 53.475 161.065 53.500 ;
        POLYGON 161.065 53.500 161.080 53.475 161.065 53.475 ;
        POLYGON 161.740 53.500 161.755 53.500 161.755 53.480 ;
        RECT 161.755 53.495 162.525 53.500 ;
        POLYGON 162.525 53.605 162.585 53.495 162.525 53.495 ;
        POLYGON 163.550 53.605 163.605 53.605 163.605 53.495 ;
        RECT 163.605 53.560 164.785 53.605 ;
        POLYGON 164.785 53.735 164.855 53.560 164.785 53.560 ;
        POLYGON 166.255 53.735 166.300 53.735 166.300 53.620 ;
        RECT 166.300 53.620 168.325 53.735 ;
        POLYGON 166.300 53.620 166.315 53.620 166.315 53.570 ;
        RECT 166.315 53.560 168.325 53.620 ;
        RECT 163.605 53.495 164.855 53.560 ;
        RECT 161.755 53.475 162.585 53.495 ;
        RECT 160.440 53.455 161.080 53.475 ;
        RECT 159.380 53.430 159.910 53.455 ;
        RECT 149.350 53.400 149.855 53.415 ;
        POLYGON 149.855 53.415 149.860 53.415 149.855 53.410 ;
        POLYGON 150.900 53.415 150.900 53.410 150.895 53.410 ;
        RECT 150.900 53.410 158.510 53.415 ;
        RECT 149.350 53.375 149.800 53.400 ;
        RECT 148.025 53.300 148.660 53.375 ;
        POLYGON 147.270 53.300 147.275 53.295 147.270 53.295 ;
        RECT 117.235 53.250 147.275 53.295 ;
        POLYGON 147.275 53.295 147.290 53.250 147.275 53.250 ;
        RECT 117.235 53.215 147.290 53.250 ;
        POLYGON 147.940 53.295 147.940 53.240 147.915 53.240 ;
        RECT 147.940 53.290 148.660 53.300 ;
        POLYGON 148.660 53.375 148.700 53.375 148.660 53.290 ;
        POLYGON 149.315 53.375 149.315 53.290 149.265 53.290 ;
        RECT 149.315 53.305 149.800 53.375 ;
        POLYGON 149.800 53.400 149.855 53.400 149.800 53.305 ;
        POLYGON 150.895 53.410 150.895 53.375 150.870 53.375 ;
        RECT 150.895 53.395 158.510 53.410 ;
        POLYGON 158.510 53.430 158.545 53.395 158.510 53.395 ;
        POLYGON 159.380 53.430 159.415 53.430 159.415 53.395 ;
        RECT 159.415 53.400 159.910 53.430 ;
        POLYGON 159.910 53.455 159.960 53.400 159.910 53.400 ;
        POLYGON 160.440 53.455 160.455 53.455 160.455 53.435 ;
        RECT 160.455 53.435 161.080 53.455 ;
        POLYGON 160.455 53.435 160.475 53.435 160.475 53.405 ;
        RECT 160.475 53.400 161.080 53.435 ;
        RECT 159.415 53.395 159.960 53.400 ;
        RECT 150.895 53.375 158.545 53.395 ;
        POLYGON 150.870 53.375 150.870 53.305 150.815 53.305 ;
        RECT 150.870 53.315 158.545 53.375 ;
        POLYGON 158.545 53.395 158.630 53.315 158.545 53.315 ;
        POLYGON 159.415 53.395 159.480 53.395 159.480 53.315 ;
        RECT 159.480 53.345 159.960 53.395 ;
        POLYGON 159.960 53.400 160.005 53.345 159.960 53.345 ;
        POLYGON 160.475 53.400 160.515 53.400 160.515 53.350 ;
        RECT 160.515 53.345 161.080 53.400 ;
        RECT 159.480 53.335 160.005 53.345 ;
        POLYGON 160.005 53.345 160.010 53.335 160.005 53.335 ;
        POLYGON 160.515 53.345 160.520 53.345 160.520 53.340 ;
        RECT 160.520 53.335 161.080 53.345 ;
        RECT 159.480 53.315 160.010 53.335 ;
        RECT 150.870 53.305 158.630 53.315 ;
        RECT 149.315 53.300 149.795 53.305 ;
        POLYGON 149.795 53.305 149.800 53.305 149.795 53.300 ;
        POLYGON 150.815 53.305 150.815 53.300 150.810 53.300 ;
        RECT 150.815 53.300 158.630 53.305 ;
        RECT 149.315 53.290 149.755 53.300 ;
        RECT 147.940 53.240 148.595 53.290 ;
        POLYGON 147.290 53.240 147.300 53.215 147.290 53.215 ;
        RECT 117.235 53.135 147.300 53.215 ;
        POLYGON 147.915 53.240 147.915 53.205 147.900 53.205 ;
        RECT 147.915 53.205 148.595 53.240 ;
        POLYGON 147.300 53.205 147.325 53.135 147.300 53.135 ;
        POLYGON 147.900 53.205 147.900 53.140 147.875 53.140 ;
        RECT 147.900 53.160 148.595 53.205 ;
        POLYGON 148.595 53.290 148.660 53.290 148.595 53.160 ;
        POLYGON 149.265 53.285 149.265 53.260 149.250 53.260 ;
        RECT 149.265 53.260 149.755 53.290 ;
        POLYGON 149.250 53.260 149.250 53.205 149.220 53.205 ;
        RECT 149.250 53.225 149.755 53.260 ;
        POLYGON 149.755 53.300 149.795 53.300 149.755 53.225 ;
        POLYGON 150.810 53.300 150.810 53.225 150.750 53.225 ;
        RECT 150.810 53.225 158.630 53.300 ;
        RECT 149.250 53.205 149.705 53.225 ;
        POLYGON 149.220 53.205 149.220 53.160 149.195 53.160 ;
        RECT 149.220 53.160 149.705 53.205 ;
        RECT 147.900 53.145 148.590 53.160 ;
        POLYGON 148.590 53.160 148.595 53.160 148.590 53.145 ;
        POLYGON 149.195 53.160 149.195 53.145 149.185 53.145 ;
        RECT 149.195 53.145 149.705 53.160 ;
        RECT 147.900 53.140 148.550 53.145 ;
        RECT 117.235 53.120 147.325 53.135 ;
        POLYGON 147.325 53.135 147.330 53.120 147.325 53.120 ;
        RECT 117.235 53.025 147.330 53.120 ;
        POLYGON 147.875 53.135 147.875 53.115 147.865 53.115 ;
        RECT 147.875 53.115 148.550 53.140 ;
        POLYGON 147.330 53.115 147.360 53.025 147.330 53.025 ;
        POLYGON 147.865 53.115 147.865 53.025 147.830 53.025 ;
        RECT 147.865 53.065 148.550 53.115 ;
        POLYGON 148.550 53.145 148.590 53.145 148.550 53.065 ;
        POLYGON 149.185 53.140 149.185 53.115 149.170 53.115 ;
        RECT 149.185 53.125 149.705 53.145 ;
        POLYGON 149.705 53.225 149.755 53.225 149.705 53.125 ;
        POLYGON 150.750 53.225 150.750 53.205 150.735 53.205 ;
        RECT 150.750 53.205 158.630 53.225 ;
        POLYGON 150.735 53.205 150.735 53.150 150.695 53.150 ;
        RECT 150.735 53.175 158.630 53.205 ;
        POLYGON 158.630 53.315 158.760 53.175 158.630 53.175 ;
        POLYGON 159.480 53.315 159.490 53.315 159.490 53.305 ;
        RECT 159.490 53.305 160.010 53.315 ;
        POLYGON 159.490 53.305 159.525 53.305 159.525 53.265 ;
        RECT 159.525 53.295 160.010 53.305 ;
        POLYGON 160.010 53.335 160.045 53.295 160.010 53.295 ;
        POLYGON 160.520 53.335 160.525 53.335 160.525 53.330 ;
        RECT 160.525 53.330 161.080 53.335 ;
        POLYGON 160.525 53.330 160.545 53.330 160.545 53.295 ;
        RECT 160.545 53.295 161.080 53.330 ;
        RECT 159.525 53.265 160.045 53.295 ;
        POLYGON 159.525 53.265 159.560 53.265 159.560 53.220 ;
        RECT 159.560 53.220 160.045 53.265 ;
        POLYGON 159.560 53.220 159.565 53.220 159.565 53.210 ;
        RECT 159.565 53.210 160.045 53.220 ;
        POLYGON 159.565 53.210 159.590 53.210 159.590 53.175 ;
        RECT 159.590 53.175 160.045 53.210 ;
        RECT 150.735 53.150 158.760 53.175 ;
        POLYGON 150.695 53.150 150.695 53.130 150.680 53.130 ;
        RECT 150.695 53.145 158.760 53.150 ;
        POLYGON 158.760 53.175 158.790 53.145 158.760 53.145 ;
        POLYGON 159.590 53.175 159.615 53.175 159.615 53.145 ;
        RECT 159.615 53.145 160.045 53.175 ;
        POLYGON 160.045 53.295 160.155 53.145 160.045 53.145 ;
        POLYGON 160.545 53.295 160.555 53.295 160.555 53.280 ;
        RECT 160.555 53.280 161.080 53.295 ;
        POLYGON 161.080 53.475 161.190 53.280 161.080 53.280 ;
        POLYGON 161.755 53.475 161.770 53.475 161.770 53.455 ;
        RECT 161.770 53.450 162.585 53.475 ;
        POLYGON 161.770 53.450 161.805 53.450 161.805 53.390 ;
        RECT 161.805 53.390 162.585 53.450 ;
        POLYGON 161.805 53.390 161.850 53.390 161.850 53.305 ;
        RECT 161.850 53.305 162.585 53.390 ;
        POLYGON 161.850 53.305 161.860 53.305 161.860 53.285 ;
        RECT 161.860 53.280 162.585 53.305 ;
        POLYGON 160.555 53.280 160.580 53.280 160.580 53.245 ;
        RECT 160.580 53.245 161.190 53.280 ;
        POLYGON 160.580 53.245 160.585 53.245 160.585 53.240 ;
        RECT 160.585 53.240 161.190 53.245 ;
        POLYGON 160.585 53.240 160.610 53.240 160.610 53.200 ;
        RECT 160.610 53.215 161.190 53.240 ;
        POLYGON 161.190 53.280 161.225 53.215 161.190 53.215 ;
        POLYGON 161.860 53.280 161.885 53.280 161.885 53.235 ;
        RECT 161.885 53.235 162.585 53.280 ;
        POLYGON 161.885 53.235 161.895 53.235 161.895 53.215 ;
        RECT 161.895 53.215 162.585 53.235 ;
        RECT 160.610 53.200 161.225 53.215 ;
        POLYGON 160.610 53.200 160.630 53.200 160.630 53.165 ;
        RECT 160.630 53.165 161.225 53.200 ;
        POLYGON 160.630 53.165 160.640 53.165 160.640 53.150 ;
        RECT 160.640 53.145 161.225 53.165 ;
        RECT 150.695 53.130 158.790 53.145 ;
        RECT 149.185 53.115 149.690 53.125 ;
        POLYGON 149.170 53.115 149.170 53.065 149.145 53.065 ;
        RECT 149.170 53.100 149.690 53.115 ;
        POLYGON 149.690 53.125 149.705 53.125 149.690 53.100 ;
        POLYGON 150.680 53.125 150.680 53.100 150.660 53.100 ;
        RECT 150.680 53.115 158.790 53.130 ;
        POLYGON 158.790 53.145 158.815 53.115 158.790 53.115 ;
        POLYGON 159.615 53.145 159.625 53.145 159.625 53.135 ;
        RECT 159.625 53.130 160.155 53.145 ;
        POLYGON 160.155 53.145 160.165 53.130 160.155 53.130 ;
        POLYGON 160.640 53.145 160.650 53.145 160.650 53.135 ;
        RECT 160.650 53.130 161.225 53.145 ;
        POLYGON 159.625 53.130 159.640 53.130 159.640 53.115 ;
        RECT 159.640 53.115 160.165 53.130 ;
        RECT 150.680 53.100 158.815 53.115 ;
        RECT 149.170 53.065 149.670 53.100 ;
        RECT 147.865 53.035 148.540 53.065 ;
        POLYGON 148.540 53.065 148.550 53.065 148.540 53.035 ;
        POLYGON 149.145 53.065 149.145 53.035 149.130 53.035 ;
        RECT 149.145 53.060 149.670 53.065 ;
        POLYGON 149.670 53.100 149.690 53.100 149.670 53.060 ;
        POLYGON 150.660 53.100 150.660 53.060 150.630 53.060 ;
        RECT 150.660 53.065 158.815 53.100 ;
        POLYGON 158.815 53.115 158.855 53.065 158.815 53.065 ;
        POLYGON 159.640 53.115 159.670 53.115 159.670 53.070 ;
        RECT 159.670 53.080 160.165 53.115 ;
        POLYGON 160.165 53.130 160.205 53.080 160.165 53.080 ;
        POLYGON 160.650 53.130 160.660 53.130 160.660 53.120 ;
        RECT 160.660 53.120 161.225 53.130 ;
        POLYGON 160.660 53.120 160.675 53.120 160.675 53.095 ;
        RECT 160.675 53.095 161.225 53.120 ;
        POLYGON 160.675 53.095 160.680 53.095 160.680 53.085 ;
        RECT 160.680 53.080 161.225 53.095 ;
        RECT 159.670 53.065 160.205 53.080 ;
        RECT 150.660 53.060 158.855 53.065 ;
        RECT 149.145 53.035 149.590 53.060 ;
        RECT 147.865 53.025 148.515 53.035 ;
        RECT 117.235 52.945 147.360 53.025 ;
        POLYGON 147.360 53.025 147.385 52.945 147.360 52.945 ;
        POLYGON 147.830 53.025 147.830 52.945 147.800 52.945 ;
        RECT 147.830 52.975 148.515 53.025 ;
        POLYGON 148.515 53.035 148.540 53.035 148.515 52.975 ;
        POLYGON 149.130 53.035 149.130 52.975 149.100 52.975 ;
        RECT 149.130 52.975 149.590 53.035 ;
        RECT 147.830 52.945 148.485 52.975 ;
        RECT 117.235 52.930 147.385 52.945 ;
        RECT 117.225 52.900 147.385 52.930 ;
        POLYGON 147.385 52.945 147.400 52.900 147.385 52.900 ;
        POLYGON 147.800 52.945 147.800 52.920 147.790 52.920 ;
        RECT 147.800 52.920 148.485 52.945 ;
        RECT 117.225 52.835 147.400 52.900 ;
        POLYGON 147.790 52.915 147.790 52.895 147.780 52.895 ;
        RECT 147.790 52.905 148.485 52.920 ;
        POLYGON 148.485 52.975 148.515 52.975 148.485 52.905 ;
        POLYGON 149.100 52.975 149.100 52.905 149.065 52.905 ;
        RECT 149.100 52.905 149.590 52.975 ;
        RECT 147.790 52.895 148.460 52.905 ;
        POLYGON 147.400 52.895 147.420 52.835 147.400 52.835 ;
        RECT 53.295 51.455 111.460 52.805 ;
        POLYGON 111.460 52.805 111.645 51.455 111.460 51.455 ;
        POLYGON 117.225 52.805 117.225 51.865 117.205 51.865 ;
        RECT 117.225 52.695 147.420 52.835 ;
        POLYGON 147.780 52.895 147.780 52.830 147.760 52.830 ;
        RECT 147.780 52.845 148.460 52.895 ;
        POLYGON 148.460 52.905 148.485 52.905 148.460 52.845 ;
        POLYGON 149.065 52.900 149.065 52.850 149.040 52.850 ;
        RECT 149.065 52.890 149.590 52.905 ;
        POLYGON 149.590 53.060 149.670 53.060 149.590 52.890 ;
        POLYGON 150.630 53.055 150.630 53.035 150.615 53.035 ;
        RECT 150.630 53.035 158.855 53.060 ;
        POLYGON 150.615 53.035 150.615 53.025 150.605 53.025 ;
        RECT 150.615 53.025 158.855 53.035 ;
        POLYGON 150.605 53.025 150.605 52.925 150.540 52.925 ;
        RECT 150.605 52.925 158.855 53.025 ;
        POLYGON 150.540 52.925 150.540 52.890 150.515 52.890 ;
        RECT 150.540 52.905 158.855 52.925 ;
        POLYGON 158.855 53.065 158.995 52.905 158.855 52.905 ;
        POLYGON 159.670 53.065 159.680 53.065 159.680 53.055 ;
        RECT 159.680 53.055 160.205 53.065 ;
        POLYGON 159.680 53.055 159.705 53.055 159.705 53.025 ;
        RECT 159.705 53.025 160.205 53.055 ;
        POLYGON 159.705 53.025 159.735 53.025 159.735 52.975 ;
        RECT 159.735 52.975 160.205 53.025 ;
        POLYGON 159.735 52.975 159.760 52.975 159.760 52.940 ;
        RECT 159.760 52.970 160.205 52.975 ;
        POLYGON 160.205 53.080 160.280 52.970 160.205 52.970 ;
        POLYGON 160.680 53.080 160.705 53.080 160.705 53.045 ;
        RECT 160.705 53.045 161.225 53.080 ;
        POLYGON 160.705 53.045 160.720 53.045 160.720 53.020 ;
        RECT 160.720 53.020 161.225 53.045 ;
        POLYGON 160.720 53.020 160.745 53.020 160.745 52.970 ;
        RECT 160.745 52.970 161.225 53.020 ;
        RECT 159.760 52.950 160.280 52.970 ;
        POLYGON 160.280 52.970 160.295 52.950 160.280 52.950 ;
        POLYGON 160.745 52.970 160.760 52.970 160.760 52.950 ;
        RECT 160.760 52.950 161.225 52.970 ;
        RECT 159.760 52.940 160.295 52.950 ;
        POLYGON 159.760 52.940 159.780 52.940 159.780 52.905 ;
        RECT 159.780 52.905 160.295 52.940 ;
        RECT 150.540 52.890 158.995 52.905 ;
        RECT 149.065 52.860 149.580 52.890 ;
        POLYGON 149.580 52.890 149.590 52.890 149.580 52.860 ;
        POLYGON 150.515 52.890 150.515 52.860 150.495 52.860 ;
        RECT 150.515 52.860 158.995 52.890 ;
        RECT 149.065 52.850 149.565 52.860 ;
        RECT 147.780 52.830 148.445 52.845 ;
        POLYGON 147.420 52.830 147.465 52.695 147.420 52.695 ;
        POLYGON 147.760 52.830 147.760 52.695 147.715 52.695 ;
        RECT 147.760 52.815 148.445 52.830 ;
        POLYGON 148.445 52.845 148.460 52.845 148.445 52.815 ;
        POLYGON 149.040 52.845 149.040 52.820 149.025 52.820 ;
        RECT 149.040 52.825 149.565 52.850 ;
        POLYGON 149.565 52.860 149.580 52.860 149.565 52.825 ;
        POLYGON 150.495 52.860 150.495 52.830 150.475 52.830 ;
        RECT 150.495 52.830 158.995 52.860 ;
        RECT 150.475 52.825 158.995 52.830 ;
        POLYGON 158.995 52.905 159.060 52.825 158.995 52.825 ;
        POLYGON 159.780 52.905 159.785 52.905 159.785 52.900 ;
        RECT 159.785 52.900 160.295 52.905 ;
        POLYGON 159.785 52.900 159.795 52.900 159.795 52.885 ;
        RECT 159.795 52.885 160.295 52.900 ;
        POLYGON 159.795 52.885 159.810 52.885 159.810 52.865 ;
        RECT 159.810 52.875 160.295 52.885 ;
        POLYGON 160.295 52.950 160.340 52.875 160.295 52.875 ;
        POLYGON 160.760 52.950 160.795 52.950 160.795 52.885 ;
        RECT 160.795 52.945 161.225 52.950 ;
        POLYGON 161.225 53.215 161.360 52.945 161.225 52.945 ;
        POLYGON 161.895 53.215 161.920 53.215 161.920 53.170 ;
        RECT 161.920 53.170 162.585 53.215 ;
        POLYGON 161.920 53.170 161.960 53.170 161.960 53.090 ;
        RECT 161.960 53.095 162.585 53.170 ;
        POLYGON 162.585 53.495 162.785 53.095 162.585 53.095 ;
        POLYGON 163.605 53.495 163.610 53.495 163.610 53.485 ;
        RECT 163.610 53.485 164.855 53.495 ;
        POLYGON 163.610 53.485 163.665 53.485 163.665 53.350 ;
        RECT 163.665 53.440 164.855 53.485 ;
        POLYGON 164.855 53.560 164.895 53.440 164.855 53.440 ;
        POLYGON 166.315 53.560 166.355 53.560 166.355 53.445 ;
        RECT 166.355 53.520 168.325 53.560 ;
        POLYGON 168.325 53.770 168.405 53.520 168.325 53.520 ;
        POLYGON 171.025 53.770 171.100 53.770 171.100 53.520 ;
        RECT 171.100 53.730 175.315 53.770 ;
        POLYGON 175.315 53.900 175.360 53.730 175.315 53.730 ;
        POLYGON 182.175 53.900 182.215 53.900 182.215 53.740 ;
        RECT 182.215 53.730 196.470 53.900 ;
        RECT 171.100 53.645 175.360 53.730 ;
        POLYGON 175.360 53.730 175.385 53.645 175.360 53.645 ;
        POLYGON 182.215 53.730 182.235 53.730 182.235 53.655 ;
        RECT 182.235 53.710 196.470 53.730 ;
        POLYGON 196.470 54.130 196.575 53.710 196.470 53.710 ;
        POLYGON 206.375 54.130 206.415 54.130 206.415 53.750 ;
        RECT 206.415 53.710 222.225 54.130 ;
        RECT 182.235 53.695 196.575 53.710 ;
        POLYGON 196.575 53.710 196.580 53.695 196.575 53.695 ;
        POLYGON 206.415 53.710 206.420 53.710 206.420 53.705 ;
        RECT 206.420 53.695 222.225 53.710 ;
        RECT 182.235 53.645 196.580 53.695 ;
        RECT 171.100 53.575 175.385 53.645 ;
        POLYGON 175.385 53.645 175.400 53.575 175.385 53.575 ;
        POLYGON 182.235 53.645 182.250 53.645 182.250 53.590 ;
        RECT 182.250 53.575 196.580 53.645 ;
        RECT 171.100 53.520 175.400 53.575 ;
        RECT 166.355 53.440 168.405 53.520 ;
        RECT 163.665 53.350 164.895 53.440 ;
        POLYGON 163.665 53.350 163.735 53.350 163.735 53.180 ;
        RECT 163.735 53.285 164.895 53.350 ;
        POLYGON 164.895 53.440 164.955 53.285 164.895 53.285 ;
        POLYGON 166.355 53.440 166.390 53.440 166.390 53.340 ;
        RECT 166.390 53.340 168.405 53.440 ;
        POLYGON 166.390 53.340 166.405 53.340 166.405 53.290 ;
        RECT 166.405 53.285 168.405 53.340 ;
        RECT 163.735 53.200 164.955 53.285 ;
        POLYGON 164.955 53.285 164.980 53.200 164.955 53.200 ;
        POLYGON 166.405 53.285 166.425 53.285 166.425 53.225 ;
        RECT 166.425 53.225 168.405 53.285 ;
        POLYGON 166.425 53.225 166.430 53.225 166.430 53.205 ;
        RECT 166.430 53.200 168.405 53.225 ;
        RECT 163.735 53.180 164.980 53.200 ;
        POLYGON 163.735 53.180 163.765 53.180 163.765 53.100 ;
        RECT 163.765 53.095 164.980 53.180 ;
        RECT 161.960 53.090 162.785 53.095 ;
        POLYGON 161.960 53.090 161.985 53.090 161.985 53.035 ;
        RECT 161.985 53.035 162.785 53.090 ;
        POLYGON 161.985 53.035 162.015 53.035 162.015 52.970 ;
        RECT 162.015 53.005 162.785 53.035 ;
        POLYGON 162.785 53.095 162.825 53.005 162.785 53.005 ;
        POLYGON 163.765 53.095 163.775 53.095 163.775 53.075 ;
        RECT 163.775 53.075 164.980 53.095 ;
        RECT 162.015 52.970 162.825 53.005 ;
        POLYGON 163.775 53.075 163.800 53.075 163.800 53.000 ;
        RECT 163.800 52.995 164.980 53.075 ;
        POLYGON 162.015 52.970 162.020 52.970 162.020 52.955 ;
        RECT 162.020 52.945 162.825 52.970 ;
        RECT 160.795 52.885 161.360 52.945 ;
        POLYGON 160.795 52.885 160.800 52.885 160.800 52.875 ;
        RECT 160.800 52.875 161.360 52.885 ;
        RECT 159.810 52.865 160.340 52.875 ;
        POLYGON 159.810 52.865 159.830 52.865 159.830 52.835 ;
        RECT 159.830 52.835 160.340 52.865 ;
        POLYGON 159.830 52.835 159.835 52.835 159.835 52.825 ;
        RECT 159.835 52.825 160.340 52.835 ;
        RECT 149.040 52.820 149.475 52.825 ;
        RECT 147.760 52.795 148.440 52.815 ;
        POLYGON 148.440 52.815 148.445 52.815 148.440 52.795 ;
        POLYGON 149.025 52.815 149.025 52.795 149.015 52.795 ;
        RECT 149.025 52.795 149.475 52.820 ;
        RECT 147.760 52.765 148.425 52.795 ;
        POLYGON 148.425 52.795 148.440 52.795 148.425 52.765 ;
        POLYGON 149.015 52.795 149.015 52.765 149.000 52.765 ;
        RECT 149.015 52.765 149.475 52.795 ;
        RECT 147.760 52.745 148.420 52.765 ;
        POLYGON 148.420 52.765 148.425 52.765 148.420 52.750 ;
        POLYGON 149.000 52.765 149.000 52.750 148.990 52.750 ;
        RECT 149.000 52.750 149.475 52.765 ;
        RECT 147.760 52.715 148.405 52.745 ;
        POLYGON 148.405 52.745 148.420 52.745 148.405 52.715 ;
        POLYGON 148.990 52.745 148.990 52.715 148.975 52.715 ;
        RECT 148.990 52.715 149.475 52.750 ;
        RECT 147.760 52.695 148.360 52.715 ;
        RECT 117.225 52.595 147.465 52.695 ;
        POLYGON 147.465 52.695 147.495 52.595 147.465 52.595 ;
        POLYGON 147.715 52.695 147.715 52.645 147.695 52.645 ;
        RECT 147.715 52.645 148.360 52.695 ;
        RECT 117.225 52.580 147.495 52.595 ;
        POLYGON 147.695 52.645 147.695 52.590 147.675 52.590 ;
        RECT 147.695 52.590 148.360 52.645 ;
        POLYGON 148.360 52.715 148.405 52.715 148.360 52.590 ;
        POLYGON 148.975 52.710 148.975 52.685 148.965 52.685 ;
        RECT 148.975 52.685 149.475 52.715 ;
        POLYGON 148.965 52.685 148.965 52.605 148.930 52.605 ;
        RECT 148.965 52.615 149.475 52.685 ;
        POLYGON 149.475 52.825 149.560 52.825 149.475 52.615 ;
        POLYGON 150.475 52.825 150.475 52.660 150.370 52.660 ;
        RECT 150.475 52.815 159.060 52.825 ;
        POLYGON 159.060 52.825 159.070 52.815 159.060 52.815 ;
        POLYGON 159.835 52.825 159.840 52.825 159.840 52.815 ;
        RECT 159.840 52.820 160.340 52.825 ;
        POLYGON 160.340 52.875 160.380 52.820 160.340 52.820 ;
        POLYGON 160.800 52.875 160.820 52.875 160.820 52.845 ;
        RECT 160.820 52.840 161.360 52.875 ;
        POLYGON 160.820 52.840 160.830 52.840 160.830 52.820 ;
        RECT 160.830 52.820 161.360 52.840 ;
        RECT 159.840 52.815 160.380 52.820 ;
        RECT 150.475 52.765 159.070 52.815 ;
        POLYGON 159.070 52.815 159.105 52.765 159.070 52.765 ;
        POLYGON 159.840 52.815 159.870 52.815 159.870 52.770 ;
        RECT 159.870 52.810 160.380 52.815 ;
        POLYGON 160.380 52.820 160.385 52.810 160.380 52.810 ;
        POLYGON 160.830 52.820 160.835 52.820 160.835 52.810 ;
        RECT 160.835 52.810 161.360 52.820 ;
        RECT 159.870 52.785 160.385 52.810 ;
        POLYGON 160.385 52.810 160.400 52.785 160.385 52.785 ;
        POLYGON 160.835 52.810 160.845 52.810 160.845 52.790 ;
        RECT 160.845 52.785 161.360 52.810 ;
        RECT 159.870 52.765 160.400 52.785 ;
        RECT 150.475 52.660 159.105 52.765 ;
        POLYGON 150.370 52.660 150.370 52.625 150.350 52.625 ;
        RECT 150.370 52.625 159.105 52.660 ;
        POLYGON 159.105 52.765 159.210 52.625 159.105 52.625 ;
        POLYGON 159.870 52.765 159.880 52.765 159.880 52.750 ;
        RECT 159.880 52.750 160.400 52.765 ;
        POLYGON 159.880 52.750 159.895 52.750 159.895 52.730 ;
        RECT 159.895 52.730 160.400 52.750 ;
        POLYGON 159.895 52.730 159.900 52.730 159.900 52.715 ;
        RECT 159.900 52.715 160.400 52.730 ;
        POLYGON 159.900 52.715 159.930 52.715 159.930 52.665 ;
        RECT 159.930 52.690 160.400 52.715 ;
        POLYGON 160.400 52.785 160.455 52.690 160.400 52.690 ;
        POLYGON 160.845 52.785 160.860 52.785 160.860 52.765 ;
        RECT 160.860 52.765 161.360 52.785 ;
        POLYGON 161.360 52.945 161.445 52.765 161.360 52.765 ;
        POLYGON 162.020 52.945 162.030 52.945 162.030 52.930 ;
        RECT 162.030 52.930 162.825 52.945 ;
        POLYGON 162.030 52.930 162.055 52.930 162.055 52.885 ;
        RECT 162.055 52.880 162.825 52.930 ;
        POLYGON 162.055 52.880 162.065 52.880 162.065 52.850 ;
        RECT 162.065 52.850 162.825 52.880 ;
        POLYGON 162.065 52.850 162.085 52.850 162.085 52.815 ;
        RECT 162.085 52.815 162.825 52.850 ;
        POLYGON 162.085 52.815 162.090 52.815 162.090 52.795 ;
        RECT 162.090 52.795 162.825 52.815 ;
        POLYGON 162.090 52.795 162.100 52.795 162.100 52.780 ;
        RECT 162.100 52.765 162.825 52.795 ;
        POLYGON 160.860 52.765 160.875 52.765 160.875 52.730 ;
        RECT 160.875 52.740 161.445 52.765 ;
        POLYGON 161.445 52.765 161.455 52.740 161.445 52.740 ;
        POLYGON 162.100 52.765 162.110 52.765 162.110 52.745 ;
        RECT 162.110 52.740 162.825 52.765 ;
        RECT 160.875 52.730 161.455 52.740 ;
        POLYGON 160.875 52.730 160.895 52.730 160.895 52.690 ;
        RECT 160.895 52.690 161.455 52.730 ;
        RECT 159.930 52.665 160.455 52.690 ;
        POLYGON 159.930 52.665 159.950 52.665 159.950 52.625 ;
        RECT 159.950 52.650 160.455 52.665 ;
        POLYGON 160.455 52.690 160.475 52.650 160.455 52.650 ;
        POLYGON 160.895 52.690 160.910 52.690 160.910 52.665 ;
        RECT 160.910 52.665 161.455 52.690 ;
        POLYGON 161.455 52.740 161.490 52.665 161.455 52.665 ;
        POLYGON 162.110 52.740 162.115 52.740 162.115 52.735 ;
        RECT 162.115 52.735 162.825 52.740 ;
        POLYGON 162.115 52.735 162.140 52.735 162.140 52.675 ;
        RECT 162.140 52.685 162.825 52.735 ;
        POLYGON 162.825 52.995 162.960 52.685 162.825 52.685 ;
        POLYGON 163.800 52.995 163.905 52.995 163.905 52.695 ;
        RECT 163.905 52.950 164.980 52.995 ;
        POLYGON 164.980 53.200 165.055 52.950 164.980 52.950 ;
        POLYGON 166.430 53.200 166.495 53.200 166.495 52.960 ;
        RECT 166.495 53.185 168.405 53.200 ;
        POLYGON 168.405 53.520 168.510 53.185 168.405 53.185 ;
        POLYGON 171.100 53.520 171.180 53.520 171.180 53.240 ;
        RECT 171.180 53.335 175.400 53.520 ;
        POLYGON 175.400 53.575 175.450 53.335 175.400 53.335 ;
        POLYGON 182.250 53.575 182.305 53.575 182.305 53.350 ;
        RECT 182.305 53.335 196.580 53.575 ;
        RECT 171.180 53.240 175.450 53.335 ;
        POLYGON 171.180 53.240 171.190 53.240 171.190 53.195 ;
        RECT 171.190 53.235 175.450 53.240 ;
        POLYGON 175.450 53.335 175.470 53.235 175.450 53.235 ;
        POLYGON 182.305 53.335 182.330 53.335 182.330 53.240 ;
        RECT 182.330 53.235 196.580 53.335 ;
        RECT 171.190 53.185 175.470 53.235 ;
        RECT 166.495 53.030 168.510 53.185 ;
        POLYGON 168.510 53.185 168.555 53.030 168.510 53.030 ;
        POLYGON 171.190 53.185 171.225 53.185 171.225 53.045 ;
        RECT 171.225 53.030 175.470 53.185 ;
        RECT 166.495 52.950 168.555 53.030 ;
        RECT 163.905 52.875 165.055 52.950 ;
        POLYGON 165.055 52.950 165.080 52.875 165.055 52.875 ;
        POLYGON 166.495 52.950 166.515 52.950 166.515 52.890 ;
        RECT 166.515 52.875 168.555 52.950 ;
        RECT 163.905 52.805 165.080 52.875 ;
        POLYGON 165.080 52.875 165.100 52.805 165.080 52.805 ;
        POLYGON 166.515 52.875 166.535 52.875 166.535 52.825 ;
        RECT 166.535 52.805 168.555 52.875 ;
        RECT 163.905 52.695 165.100 52.805 ;
        POLYGON 165.100 52.805 165.125 52.695 165.100 52.695 ;
        POLYGON 166.535 52.805 166.565 52.805 166.565 52.700 ;
        RECT 166.565 52.715 168.555 52.805 ;
        POLYGON 168.555 53.030 168.640 52.715 168.555 52.715 ;
        POLYGON 171.225 53.030 171.260 53.030 171.260 52.900 ;
        RECT 171.260 53.015 175.470 53.030 ;
        POLYGON 175.470 53.235 175.510 53.015 175.470 53.015 ;
        POLYGON 182.330 53.235 182.375 53.235 182.375 53.045 ;
        RECT 182.375 53.045 196.580 53.235 ;
        POLYGON 182.375 53.045 182.380 53.045 182.380 53.015 ;
        RECT 182.380 53.015 196.580 53.045 ;
        RECT 171.260 52.900 175.510 53.015 ;
        POLYGON 171.260 52.900 171.300 52.900 171.300 52.730 ;
        RECT 171.300 52.880 175.510 52.900 ;
        POLYGON 175.510 53.015 175.530 52.880 175.510 52.880 ;
        POLYGON 182.380 53.015 182.400 53.015 182.400 52.900 ;
        RECT 182.400 52.880 196.580 53.015 ;
        RECT 171.300 52.715 175.530 52.880 ;
        RECT 166.565 52.695 168.640 52.715 ;
        RECT 163.905 52.685 165.125 52.695 ;
        RECT 162.140 52.665 162.960 52.685 ;
        POLYGON 160.910 52.665 160.915 52.665 160.915 52.655 ;
        RECT 160.915 52.650 161.490 52.665 ;
        RECT 159.950 52.625 160.475 52.650 ;
        POLYGON 150.350 52.625 150.350 52.620 150.345 52.620 ;
        RECT 150.350 52.620 159.210 52.625 ;
        RECT 148.965 52.605 149.465 52.615 ;
        POLYGON 148.930 52.605 148.930 52.595 148.925 52.595 ;
        RECT 148.930 52.595 149.465 52.605 ;
        RECT 148.925 52.590 149.465 52.595 ;
        POLYGON 149.465 52.615 149.475 52.615 149.465 52.590 ;
        POLYGON 150.345 52.615 150.345 52.610 150.340 52.610 ;
        RECT 150.345 52.610 159.210 52.620 ;
        POLYGON 150.340 52.610 150.340 52.590 150.330 52.590 ;
        RECT 150.340 52.590 159.210 52.610 ;
        POLYGON 147.495 52.590 147.500 52.580 147.495 52.580 ;
        POLYGON 147.675 52.590 147.675 52.580 147.670 52.580 ;
        RECT 147.675 52.580 148.340 52.590 ;
        RECT 117.225 52.390 147.500 52.580 ;
        POLYGON 147.500 52.580 147.560 52.390 147.500 52.390 ;
        RECT 117.225 52.375 147.560 52.390 ;
        POLYGON 147.670 52.575 147.670 52.380 147.615 52.380 ;
        RECT 147.670 52.535 148.340 52.580 ;
        POLYGON 148.340 52.590 148.360 52.590 148.340 52.535 ;
        POLYGON 148.925 52.590 148.925 52.535 148.900 52.535 ;
        RECT 148.925 52.535 149.430 52.590 ;
        RECT 147.670 52.380 148.285 52.535 ;
        POLYGON 147.560 52.380 147.565 52.375 147.560 52.375 ;
        RECT 117.225 52.330 147.565 52.375 ;
        POLYGON 147.615 52.380 147.615 52.365 147.610 52.365 ;
        RECT 147.615 52.365 148.285 52.380 ;
        POLYGON 148.285 52.535 148.340 52.535 148.285 52.365 ;
        POLYGON 148.900 52.530 148.900 52.435 148.860 52.435 ;
        RECT 148.900 52.495 149.430 52.535 ;
        POLYGON 149.430 52.590 149.465 52.590 149.430 52.495 ;
        POLYGON 150.330 52.590 150.330 52.580 150.325 52.580 ;
        RECT 150.330 52.580 159.210 52.590 ;
        POLYGON 150.325 52.580 150.325 52.495 150.275 52.495 ;
        RECT 150.325 52.565 159.210 52.580 ;
        POLYGON 159.210 52.625 159.250 52.565 159.210 52.565 ;
        POLYGON 159.950 52.625 159.955 52.625 159.955 52.620 ;
        RECT 159.955 52.620 160.475 52.625 ;
        POLYGON 159.955 52.620 159.975 52.620 159.975 52.585 ;
        RECT 159.975 52.585 160.475 52.620 ;
        POLYGON 159.975 52.585 159.980 52.585 159.980 52.575 ;
        RECT 159.980 52.580 160.475 52.585 ;
        POLYGON 160.475 52.650 160.515 52.580 160.475 52.580 ;
        POLYGON 160.915 52.650 160.925 52.650 160.925 52.640 ;
        RECT 160.925 52.640 161.490 52.650 ;
        POLYGON 160.925 52.640 160.945 52.640 160.945 52.595 ;
        RECT 160.945 52.595 161.490 52.640 ;
        POLYGON 160.945 52.595 160.955 52.595 160.955 52.580 ;
        RECT 159.980 52.565 160.515 52.580 ;
        RECT 150.325 52.495 159.250 52.565 ;
        RECT 148.900 52.435 149.370 52.495 ;
        POLYGON 148.860 52.435 148.860 52.365 148.830 52.365 ;
        RECT 148.860 52.365 149.370 52.435 ;
        POLYGON 147.565 52.365 147.580 52.330 147.565 52.330 ;
        RECT 117.225 52.295 147.580 52.330 ;
        POLYGON 147.610 52.365 147.610 52.330 147.600 52.330 ;
        RECT 147.610 52.330 148.265 52.365 ;
        POLYGON 147.580 52.325 147.590 52.295 147.580 52.295 ;
        POLYGON 147.600 52.325 147.600 52.295 147.590 52.295 ;
        RECT 147.600 52.310 148.265 52.330 ;
        POLYGON 148.265 52.365 148.285 52.365 148.265 52.310 ;
        POLYGON 148.830 52.360 148.830 52.315 148.815 52.315 ;
        RECT 148.830 52.330 149.370 52.365 ;
        POLYGON 149.370 52.495 149.430 52.495 149.370 52.330 ;
        POLYGON 150.275 52.495 150.275 52.475 150.265 52.475 ;
        RECT 150.275 52.485 159.250 52.495 ;
        POLYGON 159.250 52.565 159.305 52.485 159.250 52.485 ;
        POLYGON 159.980 52.565 159.995 52.565 159.995 52.550 ;
        RECT 159.995 52.560 160.515 52.565 ;
        POLYGON 160.515 52.580 160.525 52.560 160.515 52.560 ;
        RECT 160.955 52.575 161.490 52.595 ;
        POLYGON 160.955 52.575 160.960 52.575 160.960 52.565 ;
        RECT 160.960 52.560 161.490 52.575 ;
        RECT 159.995 52.545 160.525 52.560 ;
        POLYGON 159.995 52.545 160.010 52.545 160.010 52.520 ;
        RECT 160.010 52.515 160.525 52.545 ;
        POLYGON 160.010 52.515 160.025 52.515 160.025 52.485 ;
        RECT 160.025 52.495 160.525 52.515 ;
        POLYGON 160.525 52.560 160.555 52.495 160.525 52.495 ;
        POLYGON 160.960 52.560 160.970 52.560 160.970 52.550 ;
        RECT 160.970 52.550 161.490 52.560 ;
        POLYGON 160.970 52.550 160.975 52.550 160.975 52.540 ;
        RECT 160.975 52.530 161.490 52.550 ;
        POLYGON 160.975 52.530 160.990 52.530 160.990 52.495 ;
        RECT 160.990 52.500 161.490 52.530 ;
        POLYGON 161.490 52.665 161.555 52.500 161.490 52.500 ;
        POLYGON 162.140 52.665 162.175 52.665 162.175 52.595 ;
        RECT 162.175 52.625 162.960 52.665 ;
        POLYGON 162.960 52.685 162.985 52.625 162.960 52.625 ;
        POLYGON 163.905 52.685 163.915 52.685 163.915 52.670 ;
        RECT 163.915 52.670 165.125 52.685 ;
        POLYGON 163.915 52.670 163.920 52.670 163.920 52.655 ;
        RECT 163.920 52.655 165.125 52.670 ;
        POLYGON 163.920 52.655 163.925 52.655 163.925 52.635 ;
        RECT 163.925 52.630 165.125 52.655 ;
        POLYGON 165.125 52.695 165.140 52.630 165.125 52.630 ;
        POLYGON 166.565 52.695 166.580 52.695 166.580 52.640 ;
        RECT 166.580 52.630 168.640 52.695 ;
        RECT 163.925 52.625 165.140 52.630 ;
        RECT 162.175 52.595 162.985 52.625 ;
        POLYGON 162.985 52.625 162.995 52.595 162.985 52.595 ;
        POLYGON 163.925 52.625 163.935 52.625 163.935 52.605 ;
        RECT 163.935 52.595 165.140 52.625 ;
        POLYGON 162.175 52.595 162.210 52.595 162.210 52.500 ;
        RECT 162.210 52.500 162.995 52.595 ;
        RECT 160.990 52.495 161.555 52.500 ;
        RECT 150.275 52.480 159.305 52.485 ;
        POLYGON 159.305 52.485 159.310 52.480 159.305 52.480 ;
        RECT 160.025 52.480 160.555 52.495 ;
        RECT 150.275 52.475 159.310 52.480 ;
        POLYGON 150.265 52.475 150.265 52.330 150.190 52.330 ;
        RECT 150.265 52.465 159.310 52.475 ;
        POLYGON 159.310 52.480 159.320 52.465 159.310 52.465 ;
        POLYGON 160.025 52.480 160.035 52.480 160.035 52.465 ;
        RECT 160.035 52.465 160.555 52.480 ;
        RECT 150.265 52.440 159.320 52.465 ;
        POLYGON 159.320 52.465 159.335 52.440 159.320 52.440 ;
        POLYGON 160.035 52.465 160.045 52.465 160.045 52.450 ;
        RECT 160.045 52.450 160.555 52.465 ;
        POLYGON 160.045 52.450 160.050 52.450 160.050 52.440 ;
        RECT 160.050 52.445 160.555 52.450 ;
        POLYGON 160.555 52.495 160.580 52.445 160.555 52.445 ;
        POLYGON 160.990 52.495 161.015 52.495 161.015 52.445 ;
        RECT 161.015 52.460 161.555 52.495 ;
        POLYGON 161.555 52.500 161.570 52.460 161.555 52.460 ;
        POLYGON 162.210 52.500 162.225 52.500 162.225 52.460 ;
        RECT 162.225 52.460 162.995 52.500 ;
        RECT 160.050 52.440 160.580 52.445 ;
        POLYGON 160.580 52.445 160.585 52.440 160.580 52.440 ;
        RECT 161.015 52.440 161.570 52.460 ;
        RECT 150.265 52.335 159.335 52.440 ;
        POLYGON 159.335 52.440 159.400 52.335 159.335 52.335 ;
        POLYGON 160.050 52.440 160.100 52.440 160.100 52.340 ;
        RECT 160.100 52.375 160.585 52.440 ;
        POLYGON 160.585 52.440 160.610 52.375 160.585 52.375 ;
        POLYGON 161.015 52.440 161.040 52.440 161.040 52.395 ;
        RECT 161.040 52.395 161.570 52.440 ;
        POLYGON 161.040 52.395 161.045 52.395 161.045 52.380 ;
        RECT 161.045 52.380 161.570 52.395 ;
        POLYGON 161.570 52.460 161.605 52.380 161.570 52.380 ;
        POLYGON 162.225 52.460 162.255 52.460 162.255 52.380 ;
        RECT 162.255 52.380 162.995 52.460 ;
        RECT 161.045 52.375 161.605 52.380 ;
        RECT 160.100 52.335 160.610 52.375 ;
        RECT 150.265 52.330 159.400 52.335 ;
        RECT 148.830 52.315 149.365 52.330 ;
        RECT 148.815 52.310 149.365 52.315 ;
        POLYGON 149.365 52.330 149.370 52.330 149.365 52.310 ;
        POLYGON 150.190 52.330 150.190 52.310 150.180 52.310 ;
        RECT 150.190 52.310 159.400 52.330 ;
        POLYGON 159.400 52.335 159.415 52.310 159.400 52.310 ;
        POLYGON 160.100 52.335 160.115 52.335 160.115 52.310 ;
        RECT 160.115 52.310 160.610 52.335 ;
        RECT 147.600 52.295 148.260 52.310 ;
        RECT 117.225 52.290 148.260 52.295 ;
        POLYGON 148.260 52.310 148.265 52.310 148.260 52.290 ;
        POLYGON 148.815 52.310 148.815 52.290 148.805 52.290 ;
        RECT 148.815 52.290 149.350 52.310 ;
        RECT 117.225 52.140 148.215 52.290 ;
        POLYGON 148.215 52.290 148.260 52.290 148.215 52.140 ;
        POLYGON 148.805 52.285 148.805 52.185 148.770 52.185 ;
        RECT 148.805 52.260 149.350 52.290 ;
        POLYGON 149.350 52.310 149.365 52.310 149.350 52.260 ;
        POLYGON 150.180 52.310 150.180 52.300 150.175 52.300 ;
        RECT 150.180 52.300 159.415 52.310 ;
        POLYGON 150.175 52.300 150.175 52.285 150.165 52.285 ;
        RECT 150.175 52.285 159.415 52.300 ;
        POLYGON 150.165 52.285 150.165 52.265 150.155 52.265 ;
        RECT 150.165 52.265 159.415 52.285 ;
        RECT 148.805 52.185 149.305 52.260 ;
        POLYGON 148.770 52.185 148.770 52.140 148.755 52.140 ;
        RECT 148.770 52.140 149.305 52.185 ;
        RECT 117.225 52.095 148.205 52.140 ;
        POLYGON 148.205 52.140 148.215 52.140 148.205 52.095 ;
        POLYGON 148.755 52.140 148.755 52.095 148.740 52.095 ;
        RECT 148.755 52.115 149.305 52.140 ;
        POLYGON 149.305 52.260 149.350 52.260 149.305 52.115 ;
        POLYGON 150.155 52.260 150.155 52.115 150.085 52.115 ;
        RECT 150.155 52.185 159.415 52.265 ;
        POLYGON 159.415 52.310 159.485 52.185 159.415 52.185 ;
        POLYGON 160.115 52.310 160.165 52.310 160.165 52.200 ;
        RECT 160.165 52.250 160.610 52.310 ;
        POLYGON 160.610 52.375 160.660 52.250 160.610 52.250 ;
        POLYGON 161.045 52.375 161.075 52.375 161.075 52.315 ;
        RECT 161.075 52.355 161.605 52.375 ;
        POLYGON 161.605 52.380 161.615 52.355 161.605 52.355 ;
        POLYGON 162.255 52.380 162.260 52.380 162.260 52.365 ;
        RECT 162.260 52.355 162.995 52.380 ;
        RECT 161.075 52.315 161.615 52.355 ;
        POLYGON 161.075 52.315 161.080 52.315 161.080 52.310 ;
        RECT 161.080 52.310 161.615 52.315 ;
        POLYGON 161.080 52.310 161.100 52.310 161.100 52.255 ;
        RECT 161.100 52.250 161.615 52.310 ;
        RECT 160.165 52.205 160.660 52.250 ;
        POLYGON 160.660 52.250 160.675 52.205 160.660 52.205 ;
        POLYGON 161.100 52.250 161.120 52.250 161.120 52.205 ;
        RECT 160.165 52.200 160.675 52.205 ;
        RECT 161.120 52.200 161.615 52.250 ;
        POLYGON 160.165 52.200 160.170 52.200 160.170 52.185 ;
        RECT 150.155 52.180 159.485 52.185 ;
        POLYGON 159.485 52.185 159.490 52.180 159.485 52.180 ;
        RECT 160.170 52.180 160.675 52.200 ;
        RECT 150.155 52.115 159.490 52.180 ;
        RECT 148.755 52.095 149.280 52.115 ;
        RECT 117.225 52.080 148.200 52.095 ;
        POLYGON 148.200 52.095 148.205 52.095 148.200 52.080 ;
        POLYGON 148.740 52.095 148.740 52.080 148.735 52.080 ;
        RECT 148.740 52.080 149.280 52.095 ;
        RECT 117.225 52.000 148.175 52.080 ;
        POLYGON 148.175 52.080 148.200 52.080 148.175 52.000 ;
        POLYGON 148.735 52.080 148.735 52.000 148.705 52.000 ;
        RECT 148.735 52.040 149.280 52.080 ;
        POLYGON 149.280 52.115 149.305 52.115 149.280 52.040 ;
        POLYGON 150.085 52.115 150.085 52.095 150.075 52.095 ;
        RECT 150.085 52.095 159.490 52.115 ;
        POLYGON 150.075 52.095 150.075 52.040 150.050 52.040 ;
        RECT 150.075 52.050 159.490 52.095 ;
        POLYGON 159.490 52.180 159.560 52.050 159.490 52.050 ;
        POLYGON 160.170 52.180 160.205 52.180 160.205 52.110 ;
        RECT 160.205 52.115 160.675 52.180 ;
        POLYGON 160.675 52.200 160.705 52.115 160.675 52.115 ;
        POLYGON 161.120 52.200 161.155 52.200 161.155 52.120 ;
        RECT 161.155 52.180 161.615 52.200 ;
        POLYGON 161.615 52.355 161.675 52.180 161.615 52.180 ;
        POLYGON 162.260 52.355 162.285 52.355 162.285 52.300 ;
        RECT 162.285 52.300 162.995 52.355 ;
        POLYGON 162.285 52.300 162.325 52.300 162.325 52.180 ;
        RECT 162.325 52.275 162.995 52.300 ;
        POLYGON 162.995 52.595 163.115 52.275 162.995 52.275 ;
        POLYGON 163.935 52.595 164.010 52.595 164.010 52.370 ;
        RECT 164.010 52.430 165.140 52.595 ;
        POLYGON 165.140 52.630 165.190 52.430 165.140 52.430 ;
        POLYGON 166.580 52.630 166.630 52.630 166.630 52.440 ;
        RECT 166.630 52.530 168.640 52.630 ;
        POLYGON 168.640 52.715 168.685 52.530 168.640 52.530 ;
        POLYGON 171.300 52.715 171.345 52.715 171.345 52.545 ;
        RECT 171.345 52.675 175.530 52.715 ;
        POLYGON 175.530 52.880 175.555 52.675 175.530 52.675 ;
        POLYGON 182.400 52.880 182.435 52.880 182.435 52.695 ;
        RECT 182.435 52.675 196.580 52.880 ;
        RECT 171.345 52.530 175.555 52.675 ;
        RECT 166.630 52.430 168.685 52.530 ;
        RECT 164.010 52.370 165.190 52.430 ;
        POLYGON 164.010 52.370 164.035 52.370 164.035 52.285 ;
        RECT 164.035 52.295 165.190 52.370 ;
        POLYGON 165.190 52.430 165.220 52.295 165.190 52.295 ;
        POLYGON 166.630 52.430 166.635 52.430 166.635 52.420 ;
        RECT 166.635 52.420 168.685 52.430 ;
        POLYGON 166.635 52.420 166.655 52.420 166.655 52.310 ;
        RECT 166.655 52.295 168.685 52.420 ;
        RECT 164.035 52.275 165.220 52.295 ;
        RECT 162.325 52.265 163.115 52.275 ;
        POLYGON 163.115 52.275 163.120 52.265 163.115 52.265 ;
        POLYGON 164.035 52.275 164.040 52.275 164.040 52.265 ;
        RECT 164.040 52.265 165.220 52.275 ;
        RECT 162.325 52.180 163.120 52.265 ;
        POLYGON 163.120 52.265 163.145 52.180 163.120 52.180 ;
        POLYGON 164.040 52.265 164.050 52.265 164.050 52.235 ;
        RECT 164.050 52.235 165.220 52.265 ;
        POLYGON 164.050 52.235 164.060 52.235 164.060 52.190 ;
        RECT 164.060 52.180 165.220 52.235 ;
        RECT 161.155 52.115 161.675 52.180 ;
        RECT 160.205 52.110 160.705 52.115 ;
        POLYGON 160.205 52.110 160.215 52.110 160.215 52.100 ;
        RECT 160.215 52.100 160.705 52.110 ;
        POLYGON 160.215 52.100 160.230 52.100 160.230 52.060 ;
        RECT 160.230 52.060 160.705 52.100 ;
        POLYGON 160.705 52.115 160.720 52.060 160.705 52.060 ;
        POLYGON 161.155 52.115 161.175 52.115 161.175 52.070 ;
        RECT 161.175 52.085 161.675 52.115 ;
        POLYGON 161.675 52.180 161.710 52.085 161.675 52.085 ;
        POLYGON 162.325 52.180 162.355 52.180 162.355 52.090 ;
        RECT 162.355 52.085 163.145 52.180 ;
        RECT 161.175 52.060 161.710 52.085 ;
        RECT 160.230 52.050 160.720 52.060 ;
        RECT 150.075 52.040 159.560 52.050 ;
        RECT 148.735 52.000 149.185 52.040 ;
        RECT 117.225 51.910 148.150 52.000 ;
        POLYGON 148.150 52.000 148.175 52.000 148.150 51.910 ;
        POLYGON 148.705 51.995 148.705 51.980 148.700 51.980 ;
        RECT 148.705 51.980 149.185 52.000 ;
        POLYGON 148.700 51.980 148.700 51.910 148.680 51.910 ;
        RECT 148.700 51.910 149.185 51.980 ;
        RECT 117.225 51.865 148.140 51.910 ;
        RECT 117.205 51.855 148.140 51.865 ;
        POLYGON 148.140 51.910 148.150 51.910 148.140 51.855 ;
        POLYGON 148.680 51.905 148.680 51.865 148.670 51.865 ;
        RECT 148.680 51.865 149.185 51.910 ;
        POLYGON 117.205 51.785 117.205 51.455 117.195 51.455 ;
        RECT 117.205 51.750 148.115 51.855 ;
        POLYGON 148.115 51.855 148.140 51.855 148.115 51.750 ;
        POLYGON 148.670 51.855 148.670 51.825 148.660 51.825 ;
        RECT 148.670 51.825 149.185 51.865 ;
        POLYGON 148.660 51.825 148.660 51.750 148.640 51.750 ;
        RECT 148.660 51.750 149.185 51.825 ;
        RECT 117.205 51.685 148.100 51.750 ;
        POLYGON 148.100 51.750 148.115 51.750 148.100 51.685 ;
        POLYGON 148.640 51.750 148.640 51.685 148.620 51.685 ;
        RECT 148.640 51.685 149.185 51.750 ;
        RECT 117.205 51.625 148.085 51.685 ;
        POLYGON 148.085 51.685 148.100 51.685 148.085 51.625 ;
        POLYGON 148.620 51.680 148.620 51.630 148.605 51.630 ;
        RECT 148.620 51.660 149.185 51.685 ;
        POLYGON 149.185 52.040 149.280 52.040 149.185 51.660 ;
        POLYGON 150.050 52.035 150.050 51.945 150.010 51.945 ;
        RECT 150.050 51.945 159.560 52.040 ;
        POLYGON 150.010 51.940 150.010 51.900 149.995 51.900 ;
        RECT 150.010 51.920 159.560 51.945 ;
        POLYGON 159.560 52.050 159.625 51.920 159.560 51.920 ;
        POLYGON 160.230 52.050 160.280 52.050 160.280 51.935 ;
        RECT 160.280 51.965 160.720 52.050 ;
        POLYGON 160.720 52.060 160.745 51.965 160.720 51.965 ;
        POLYGON 161.175 52.060 161.185 52.060 161.185 52.045 ;
        RECT 161.185 52.045 161.710 52.060 ;
        POLYGON 161.185 52.045 161.190 52.045 161.190 52.035 ;
        RECT 161.190 52.035 161.710 52.045 ;
        POLYGON 161.190 52.035 161.210 52.035 161.210 51.975 ;
        RECT 161.210 51.965 161.710 52.035 ;
        RECT 160.280 51.935 160.745 51.965 ;
        POLYGON 160.280 51.935 160.285 51.935 160.285 51.920 ;
        RECT 150.010 51.900 159.625 51.920 ;
        RECT 160.285 51.915 160.745 51.935 ;
        POLYGON 160.745 51.965 160.760 51.915 160.745 51.915 ;
        POLYGON 161.210 51.965 161.225 51.965 161.225 51.930 ;
        RECT 161.225 51.930 161.710 51.965 ;
        POLYGON 161.225 51.930 161.230 51.930 161.230 51.915 ;
        RECT 161.230 51.915 161.710 51.930 ;
        POLYGON 149.995 51.900 149.995 51.705 149.920 51.705 ;
        RECT 149.995 51.890 159.625 51.900 ;
        POLYGON 159.625 51.915 159.640 51.890 159.625 51.890 ;
        POLYGON 160.285 51.915 160.295 51.915 160.295 51.895 ;
        RECT 160.295 51.890 160.760 51.915 ;
        RECT 149.995 51.785 159.640 51.890 ;
        POLYGON 159.640 51.890 159.680 51.785 159.640 51.785 ;
        POLYGON 160.295 51.890 160.300 51.890 160.300 51.885 ;
        RECT 160.300 51.885 160.760 51.890 ;
        POLYGON 160.300 51.885 160.335 51.885 160.335 51.790 ;
        RECT 160.335 51.785 160.760 51.885 ;
        RECT 149.995 51.740 159.680 51.785 ;
        POLYGON 159.680 51.785 159.705 51.740 159.680 51.740 ;
        POLYGON 160.335 51.785 160.350 51.785 160.350 51.750 ;
        RECT 160.350 51.770 160.760 51.785 ;
        POLYGON 160.760 51.915 160.795 51.770 160.760 51.770 ;
        POLYGON 161.230 51.915 161.280 51.915 161.280 51.775 ;
        RECT 161.280 51.890 161.710 51.915 ;
        POLYGON 161.710 52.085 161.770 51.890 161.710 51.890 ;
        POLYGON 162.355 52.085 162.365 52.085 162.365 52.060 ;
        RECT 162.365 52.060 163.145 52.085 ;
        POLYGON 162.365 52.060 162.380 52.060 162.380 52.000 ;
        RECT 162.380 52.000 163.145 52.060 ;
        POLYGON 162.380 52.000 162.410 52.000 162.410 51.895 ;
        RECT 162.410 51.960 163.145 52.000 ;
        POLYGON 163.145 52.180 163.215 51.960 163.145 51.960 ;
        POLYGON 164.060 52.180 164.115 52.180 164.115 51.965 ;
        RECT 164.115 51.960 165.220 52.180 ;
        RECT 161.280 51.785 161.770 51.890 ;
        RECT 162.410 51.885 163.215 51.960 ;
        POLYGON 161.770 51.885 161.805 51.785 161.770 51.785 ;
        POLYGON 162.410 51.885 162.440 51.885 162.440 51.785 ;
        RECT 162.440 51.860 163.215 51.885 ;
        POLYGON 163.215 51.960 163.245 51.860 163.215 51.860 ;
        POLYGON 164.115 51.960 164.140 51.960 164.140 51.865 ;
        RECT 164.140 51.935 165.220 51.960 ;
        POLYGON 165.220 52.295 165.290 51.935 165.220 51.935 ;
        POLYGON 166.655 52.295 166.665 52.295 166.665 52.260 ;
        RECT 166.665 52.260 168.685 52.295 ;
        POLYGON 166.665 52.260 166.720 52.260 166.720 52.005 ;
        RECT 166.720 52.245 168.685 52.260 ;
        POLYGON 168.685 52.530 168.755 52.245 168.685 52.245 ;
        POLYGON 171.345 52.530 171.350 52.530 171.350 52.525 ;
        RECT 171.350 52.525 175.555 52.530 ;
        RECT 166.720 52.035 168.755 52.245 ;
        POLYGON 171.350 52.525 171.405 52.525 171.405 52.230 ;
        RECT 171.405 52.390 175.555 52.525 ;
        POLYGON 175.555 52.675 175.575 52.390 175.555 52.390 ;
        POLYGON 182.435 52.675 182.485 52.675 182.485 52.410 ;
        RECT 182.485 52.590 196.580 52.675 ;
        POLYGON 196.580 53.695 196.860 52.590 196.580 52.590 ;
        POLYGON 206.420 53.695 206.440 53.695 206.440 53.515 ;
        RECT 206.440 53.515 222.225 53.695 ;
        POLYGON 206.440 53.515 206.510 53.515 206.510 52.800 ;
        RECT 206.510 52.800 222.225 53.515 ;
        POLYGON 222.225 55.655 222.255 55.655 222.225 53.075 ;
        POLYGON 229.525 55.650 229.525 55.445 229.485 55.445 ;
        RECT 229.525 55.615 233.815 55.655 ;
        POLYGON 233.815 56.245 234.010 56.245 233.815 55.625 ;
        POLYGON 237.100 56.240 237.100 56.075 237.025 56.075 ;
        RECT 237.100 56.175 239.340 56.245 ;
        POLYGON 239.340 56.385 239.450 56.385 239.340 56.175 ;
        POLYGON 241.245 56.385 241.245 56.175 241.115 56.175 ;
        RECT 241.245 56.215 242.685 56.385 ;
        POLYGON 242.685 56.400 242.840 56.400 242.685 56.215 ;
        POLYGON 244.180 56.400 244.180 56.320 244.100 56.320 ;
        RECT 244.180 56.380 245.250 56.400 ;
        POLYGON 245.250 56.445 245.335 56.445 245.250 56.380 ;
        POLYGON 246.705 56.445 246.705 56.415 246.655 56.415 ;
        RECT 246.705 56.415 247.945 56.445 ;
        POLYGON 246.655 56.415 246.655 56.380 246.595 56.380 ;
        RECT 246.655 56.380 247.945 56.415 ;
        RECT 244.180 56.320 245.115 56.380 ;
        POLYGON 244.100 56.320 244.100 56.235 244.020 56.235 ;
        RECT 244.100 56.265 245.115 56.320 ;
        POLYGON 245.115 56.380 245.250 56.380 245.115 56.265 ;
        POLYGON 246.595 56.380 246.595 56.350 246.540 56.350 ;
        RECT 246.595 56.360 247.945 56.380 ;
        POLYGON 247.945 56.445 248.200 56.445 247.945 56.360 ;
        POLYGON 252.450 56.445 252.500 56.445 252.500 56.430 ;
        RECT 252.500 56.430 253.800 56.445 ;
        POLYGON 252.500 56.430 252.510 56.430 252.510 56.425 ;
        RECT 252.510 56.425 253.800 56.430 ;
        POLYGON 252.510 56.425 252.540 56.425 252.540 56.415 ;
        RECT 252.540 56.415 253.800 56.425 ;
        POLYGON 252.545 56.415 252.680 56.415 252.680 56.360 ;
        RECT 252.680 56.400 253.800 56.415 ;
        POLYGON 253.800 56.450 253.880 56.400 253.800 56.400 ;
        POLYGON 255.060 56.450 255.070 56.450 255.070 56.445 ;
        RECT 255.070 56.445 256.275 56.450 ;
        POLYGON 255.070 56.445 255.125 56.445 255.125 56.400 ;
        RECT 255.125 56.400 256.275 56.445 ;
        POLYGON 256.275 56.615 256.515 56.400 256.275 56.400 ;
        POLYGON 257.870 56.615 257.935 56.615 257.935 56.545 ;
        RECT 257.935 56.545 259.655 56.615 ;
        POLYGON 257.935 56.545 257.975 56.545 257.975 56.500 ;
        RECT 257.975 56.505 259.655 56.545 ;
        POLYGON 259.655 56.720 259.815 56.505 259.655 56.505 ;
        POLYGON 261.910 56.720 261.930 56.720 261.930 56.685 ;
        RECT 261.930 56.685 264.755 56.720 ;
        POLYGON 261.930 56.685 261.955 56.685 261.955 56.645 ;
        RECT 261.955 56.645 264.755 56.685 ;
        POLYGON 261.955 56.645 261.960 56.645 261.960 56.640 ;
        RECT 261.960 56.640 264.755 56.645 ;
        POLYGON 261.960 56.640 262.045 56.640 262.045 56.505 ;
        RECT 257.975 56.500 259.815 56.505 ;
        POLYGON 259.815 56.505 259.820 56.500 259.815 56.500 ;
        RECT 262.045 56.500 264.755 56.640 ;
        POLYGON 257.975 56.500 257.990 56.500 257.990 56.485 ;
        RECT 257.990 56.485 259.820 56.500 ;
        POLYGON 257.990 56.485 258.060 56.485 258.060 56.400 ;
        RECT 258.060 56.455 259.820 56.485 ;
        POLYGON 259.820 56.500 259.855 56.455 259.820 56.455 ;
        POLYGON 262.045 56.500 262.075 56.500 262.075 56.455 ;
        RECT 262.075 56.455 264.755 56.500 ;
        RECT 258.060 56.400 259.855 56.455 ;
        RECT 252.680 56.360 253.880 56.400 ;
        RECT 246.595 56.350 247.830 56.360 ;
        POLYGON 246.540 56.350 246.540 56.345 246.530 56.345 ;
        RECT 246.540 56.345 247.830 56.350 ;
        POLYGON 246.530 56.345 246.530 56.330 246.505 56.330 ;
        RECT 246.530 56.330 247.830 56.345 ;
        POLYGON 246.505 56.330 246.505 56.265 246.400 56.265 ;
        RECT 246.505 56.315 247.830 56.330 ;
        POLYGON 247.830 56.360 247.945 56.360 247.830 56.315 ;
        POLYGON 252.690 56.360 252.760 56.360 252.760 56.330 ;
        RECT 252.760 56.330 253.880 56.360 ;
        POLYGON 253.880 56.400 253.995 56.330 253.880 56.330 ;
        POLYGON 255.125 56.400 255.165 56.400 255.165 56.370 ;
        RECT 255.165 56.370 256.515 56.400 ;
        POLYGON 255.165 56.370 255.170 56.370 255.170 56.365 ;
        RECT 255.170 56.365 256.515 56.370 ;
        POLYGON 255.175 56.365 255.215 56.365 255.215 56.330 ;
        RECT 255.215 56.345 256.515 56.365 ;
        POLYGON 256.515 56.400 256.570 56.345 256.515 56.345 ;
        POLYGON 258.060 56.400 258.110 56.400 258.110 56.345 ;
        RECT 258.110 56.345 259.855 56.400 ;
        RECT 255.215 56.330 256.570 56.345 ;
        POLYGON 252.760 56.330 252.790 56.330 252.790 56.315 ;
        RECT 252.790 56.325 253.995 56.330 ;
        POLYGON 253.995 56.330 254.000 56.325 253.995 56.325 ;
        POLYGON 255.215 56.330 255.220 56.330 255.220 56.325 ;
        RECT 255.220 56.325 256.570 56.330 ;
        RECT 252.790 56.320 254.005 56.325 ;
        POLYGON 254.005 56.325 254.015 56.320 254.005 56.320 ;
        POLYGON 255.220 56.325 255.225 56.325 255.225 56.320 ;
        RECT 255.225 56.320 256.570 56.325 ;
        RECT 252.790 56.315 254.015 56.320 ;
        RECT 246.505 56.295 247.785 56.315 ;
        POLYGON 247.785 56.315 247.830 56.315 247.785 56.295 ;
        POLYGON 252.790 56.315 252.830 56.315 252.830 56.300 ;
        RECT 252.830 56.300 254.015 56.315 ;
        POLYGON 252.830 56.300 252.840 56.300 252.840 56.295 ;
        RECT 252.840 56.295 254.015 56.300 ;
        RECT 246.505 56.265 247.695 56.295 ;
        RECT 244.100 56.260 245.110 56.265 ;
        POLYGON 245.110 56.265 245.115 56.265 245.110 56.260 ;
        POLYGON 246.400 56.265 246.400 56.260 246.395 56.260 ;
        RECT 246.400 56.260 247.695 56.265 ;
        POLYGON 247.695 56.295 247.785 56.295 247.695 56.260 ;
        POLYGON 252.840 56.295 252.930 56.295 252.930 56.260 ;
        RECT 252.930 56.260 254.015 56.295 ;
        RECT 244.100 56.235 245.065 56.260 ;
        POLYGON 244.020 56.235 244.020 56.215 244.000 56.215 ;
        RECT 244.020 56.225 245.065 56.235 ;
        POLYGON 245.065 56.260 245.110 56.260 245.065 56.225 ;
        POLYGON 246.395 56.260 246.395 56.225 246.335 56.225 ;
        RECT 246.395 56.225 247.555 56.260 ;
        RECT 244.020 56.215 244.905 56.225 ;
        RECT 241.245 56.175 242.585 56.215 ;
        RECT 237.100 56.075 239.205 56.175 ;
        POLYGON 237.025 56.075 237.025 56.035 237.005 56.035 ;
        RECT 237.025 56.035 239.205 56.075 ;
        POLYGON 237.005 56.035 237.005 55.675 236.875 55.675 ;
        RECT 237.005 55.905 239.205 56.035 ;
        POLYGON 239.205 56.175 239.340 56.175 239.205 55.905 ;
        POLYGON 241.115 56.175 241.115 56.135 241.090 56.135 ;
        RECT 241.115 56.135 242.585 56.175 ;
        POLYGON 241.090 56.135 241.090 56.005 241.015 56.005 ;
        RECT 241.090 56.095 242.585 56.135 ;
        POLYGON 242.585 56.215 242.685 56.215 242.585 56.095 ;
        POLYGON 244.000 56.215 244.000 56.165 243.955 56.165 ;
        RECT 244.000 56.165 244.905 56.215 ;
        POLYGON 243.955 56.165 243.955 56.095 243.890 56.095 ;
        RECT 243.955 56.095 244.905 56.165 ;
        RECT 241.090 56.015 242.525 56.095 ;
        POLYGON 242.525 56.095 242.585 56.095 242.525 56.020 ;
        POLYGON 243.890 56.090 243.890 56.070 243.870 56.070 ;
        RECT 243.890 56.075 244.905 56.095 ;
        POLYGON 244.905 56.225 245.065 56.225 244.905 56.075 ;
        POLYGON 246.335 56.225 246.335 56.190 246.280 56.190 ;
        RECT 246.335 56.200 247.555 56.225 ;
        POLYGON 247.555 56.260 247.690 56.260 247.555 56.200 ;
        POLYGON 252.930 56.260 252.940 56.260 252.940 56.255 ;
        RECT 252.940 56.255 254.015 56.260 ;
        POLYGON 250.180 56.255 250.180 56.250 250.055 56.250 ;
        RECT 250.180 56.250 250.220 56.255 ;
        POLYGON 250.220 56.255 250.255 56.250 250.220 56.250 ;
        POLYGON 252.940 56.255 252.950 56.255 252.950 56.250 ;
        RECT 252.950 56.250 254.015 56.255 ;
        POLYGON 250.040 56.250 250.040 56.245 249.930 56.245 ;
        RECT 250.040 56.245 250.445 56.250 ;
        POLYGON 250.445 56.250 250.565 56.245 250.445 56.245 ;
        POLYGON 252.950 56.250 252.960 56.250 252.960 56.245 ;
        RECT 252.960 56.245 254.015 56.250 ;
        POLYGON 254.015 56.320 254.130 56.245 254.015 56.245 ;
        POLYGON 255.225 56.320 255.240 56.320 255.240 56.310 ;
        RECT 255.240 56.310 256.570 56.320 ;
        POLYGON 255.240 56.310 255.285 56.310 255.285 56.270 ;
        RECT 255.285 56.270 256.570 56.310 ;
        POLYGON 255.290 56.270 255.320 56.270 255.320 56.245 ;
        RECT 255.320 56.245 256.570 56.270 ;
        POLYGON 249.845 56.245 249.845 56.240 249.780 56.240 ;
        RECT 249.845 56.240 250.595 56.245 ;
        POLYGON 250.595 56.245 250.695 56.240 250.595 56.240 ;
        POLYGON 252.960 56.245 252.970 56.245 252.970 56.240 ;
        RECT 252.970 56.240 254.135 56.245 ;
        POLYGON 249.770 56.240 249.770 56.235 249.655 56.235 ;
        RECT 249.770 56.235 250.705 56.240 ;
        POLYGON 249.650 56.235 249.650 56.225 249.515 56.225 ;
        RECT 249.650 56.230 250.705 56.235 ;
        POLYGON 250.705 56.240 250.860 56.230 250.705 56.230 ;
        POLYGON 252.975 56.240 252.995 56.240 252.995 56.230 ;
        RECT 252.995 56.230 254.135 56.240 ;
        RECT 249.650 56.225 250.865 56.230 ;
        POLYGON 250.865 56.230 250.930 56.225 250.865 56.225 ;
        POLYGON 252.995 56.230 253.010 56.230 253.010 56.225 ;
        RECT 253.010 56.225 254.135 56.230 ;
        POLYGON 249.505 56.225 249.505 56.220 249.500 56.220 ;
        RECT 249.505 56.220 250.930 56.225 ;
        POLYGON 250.930 56.225 250.965 56.220 250.930 56.220 ;
        POLYGON 253.010 56.225 253.020 56.225 253.020 56.220 ;
        RECT 253.020 56.220 254.135 56.225 ;
        POLYGON 249.495 56.220 249.495 56.210 249.390 56.210 ;
        RECT 249.495 56.210 250.965 56.220 ;
        POLYGON 249.385 56.210 249.385 56.200 249.290 56.200 ;
        RECT 249.385 56.205 250.965 56.210 ;
        POLYGON 250.965 56.220 251.125 56.205 250.965 56.205 ;
        POLYGON 253.020 56.220 253.050 56.220 253.050 56.205 ;
        RECT 253.050 56.205 254.135 56.220 ;
        RECT 249.385 56.200 251.135 56.205 ;
        RECT 246.335 56.190 247.515 56.200 ;
        POLYGON 246.275 56.190 246.275 56.165 246.240 56.165 ;
        RECT 246.275 56.180 247.515 56.190 ;
        POLYGON 247.515 56.200 247.555 56.200 247.515 56.180 ;
        POLYGON 249.290 56.200 249.290 56.195 249.240 56.195 ;
        RECT 249.290 56.195 251.135 56.200 ;
        POLYGON 251.135 56.205 251.220 56.195 251.135 56.195 ;
        POLYGON 253.050 56.205 253.070 56.205 253.070 56.195 ;
        RECT 253.070 56.195 254.135 56.205 ;
        POLYGON 249.235 56.195 249.235 56.190 249.225 56.190 ;
        RECT 249.235 56.190 251.225 56.195 ;
        POLYGON 249.190 56.190 249.190 56.180 249.145 56.180 ;
        RECT 249.190 56.185 251.225 56.190 ;
        POLYGON 251.225 56.195 251.275 56.185 251.225 56.185 ;
        POLYGON 253.070 56.195 253.090 56.195 253.090 56.185 ;
        RECT 253.090 56.185 254.135 56.195 ;
        POLYGON 254.135 56.245 254.220 56.185 254.135 56.185 ;
        POLYGON 255.320 56.245 255.390 56.245 255.390 56.185 ;
        RECT 255.390 56.185 256.570 56.245 ;
        RECT 249.190 56.180 251.275 56.185 ;
        RECT 246.275 56.165 247.455 56.180 ;
        POLYGON 246.235 56.165 246.235 56.075 246.100 56.075 ;
        RECT 246.235 56.155 247.455 56.165 ;
        POLYGON 247.455 56.180 247.515 56.180 247.455 56.155 ;
        POLYGON 249.145 56.180 249.145 56.175 249.120 56.175 ;
        RECT 249.145 56.175 251.275 56.180 ;
        POLYGON 249.120 56.175 249.120 56.155 248.975 56.155 ;
        RECT 249.120 56.170 251.275 56.175 ;
        POLYGON 251.275 56.185 251.400 56.170 251.275 56.170 ;
        POLYGON 253.090 56.185 253.115 56.185 253.115 56.175 ;
        RECT 253.115 56.175 254.220 56.185 ;
        POLYGON 254.220 56.185 254.235 56.175 254.220 56.175 ;
        POLYGON 255.390 56.185 255.405 56.185 255.405 56.175 ;
        RECT 255.405 56.175 256.570 56.185 ;
        POLYGON 253.115 56.175 253.125 56.175 253.125 56.170 ;
        RECT 253.125 56.170 254.235 56.175 ;
        RECT 249.120 56.165 251.400 56.170 ;
        POLYGON 251.400 56.170 251.405 56.165 251.400 56.165 ;
        POLYGON 253.125 56.170 253.135 56.170 253.135 56.165 ;
        RECT 253.135 56.165 254.235 56.170 ;
        RECT 249.120 56.155 251.405 56.165 ;
        POLYGON 251.405 56.165 251.485 56.155 251.405 56.155 ;
        POLYGON 253.135 56.165 253.155 56.165 253.155 56.155 ;
        RECT 253.155 56.155 254.235 56.165 ;
        RECT 246.235 56.135 247.415 56.155 ;
        POLYGON 247.415 56.155 247.455 56.155 247.415 56.135 ;
        POLYGON 248.975 56.155 248.975 56.150 248.945 56.150 ;
        RECT 248.975 56.150 251.485 56.155 ;
        POLYGON 248.945 56.150 248.945 56.140 248.875 56.140 ;
        RECT 248.945 56.140 251.485 56.150 ;
        POLYGON 248.875 56.140 248.875 56.135 248.850 56.135 ;
        RECT 248.875 56.135 251.485 56.140 ;
        POLYGON 251.485 56.155 251.610 56.135 251.485 56.135 ;
        POLYGON 253.155 56.155 253.170 56.155 253.170 56.150 ;
        RECT 253.170 56.150 254.235 56.155 ;
        POLYGON 253.170 56.150 253.200 56.150 253.200 56.135 ;
        RECT 253.200 56.135 254.235 56.150 ;
        RECT 246.235 56.075 247.275 56.135 ;
        RECT 243.890 56.070 244.890 56.075 ;
        POLYGON 243.870 56.070 243.870 56.020 243.825 56.020 ;
        RECT 243.870 56.065 244.890 56.070 ;
        POLYGON 244.890 56.075 244.905 56.075 244.890 56.065 ;
        POLYGON 246.100 56.075 246.100 56.065 246.085 56.065 ;
        RECT 246.100 56.070 247.275 56.075 ;
        POLYGON 247.275 56.135 247.415 56.135 247.275 56.070 ;
        POLYGON 248.850 56.135 248.850 56.105 248.710 56.105 ;
        RECT 248.850 56.125 251.610 56.135 ;
        POLYGON 251.610 56.135 251.660 56.125 251.610 56.125 ;
        POLYGON 253.200 56.135 253.220 56.135 253.220 56.125 ;
        RECT 253.220 56.125 254.235 56.135 ;
        RECT 248.850 56.120 251.660 56.125 ;
        POLYGON 251.660 56.125 251.680 56.120 251.660 56.120 ;
        POLYGON 253.220 56.125 253.230 56.125 253.230 56.120 ;
        RECT 253.230 56.120 254.235 56.125 ;
        POLYGON 254.235 56.175 254.315 56.120 254.235 56.120 ;
        POLYGON 255.405 56.175 255.460 56.175 255.460 56.130 ;
        RECT 255.460 56.165 256.570 56.175 ;
        POLYGON 256.570 56.345 256.755 56.165 256.570 56.165 ;
        POLYGON 258.110 56.345 258.120 56.345 258.120 56.335 ;
        RECT 258.120 56.335 259.855 56.345 ;
        POLYGON 258.120 56.335 258.140 56.335 258.140 56.310 ;
        RECT 258.140 56.310 259.855 56.335 ;
        POLYGON 258.140 56.310 258.155 56.310 258.155 56.295 ;
        RECT 258.155 56.295 259.855 56.310 ;
        POLYGON 258.155 56.295 258.245 56.295 258.245 56.180 ;
        RECT 258.245 56.180 259.855 56.295 ;
        POLYGON 258.245 56.180 258.255 56.180 258.255 56.165 ;
        RECT 258.255 56.165 259.855 56.180 ;
        RECT 255.460 56.150 256.755 56.165 ;
        POLYGON 256.755 56.165 256.765 56.150 256.755 56.150 ;
        POLYGON 258.255 56.165 258.270 56.165 258.270 56.150 ;
        RECT 258.270 56.150 259.855 56.165 ;
        RECT 255.460 56.130 256.765 56.150 ;
        POLYGON 255.460 56.130 255.470 56.130 255.470 56.120 ;
        RECT 255.470 56.120 256.765 56.130 ;
        RECT 248.850 56.105 251.680 56.120 ;
        POLYGON 251.680 56.120 251.745 56.105 251.680 56.105 ;
        POLYGON 253.230 56.120 253.260 56.120 253.260 56.105 ;
        RECT 253.260 56.105 254.315 56.120 ;
        POLYGON 248.710 56.105 248.710 56.095 248.665 56.095 ;
        RECT 248.710 56.095 251.745 56.105 ;
        POLYGON 248.665 56.095 248.665 56.080 248.585 56.080 ;
        RECT 248.665 56.080 251.745 56.095 ;
        POLYGON 248.585 56.080 248.585 56.070 248.545 56.070 ;
        RECT 248.585 56.070 251.745 56.080 ;
        POLYGON 251.745 56.105 251.920 56.070 251.745 56.070 ;
        POLYGON 253.260 56.105 253.305 56.105 253.305 56.080 ;
        RECT 253.305 56.080 254.315 56.105 ;
        POLYGON 253.305 56.080 253.325 56.080 253.325 56.070 ;
        RECT 253.325 56.075 254.315 56.080 ;
        POLYGON 254.315 56.120 254.380 56.075 254.315 56.075 ;
        POLYGON 255.470 56.120 255.515 56.120 255.515 56.075 ;
        RECT 255.515 56.075 256.765 56.120 ;
        RECT 253.325 56.070 254.380 56.075 ;
        RECT 246.100 56.065 247.250 56.070 ;
        RECT 243.870 56.020 244.845 56.065 ;
        RECT 241.090 56.005 242.370 56.015 ;
        POLYGON 241.015 56.005 241.015 56.000 241.010 56.000 ;
        RECT 241.015 56.000 242.370 56.005 ;
        POLYGON 241.010 56.000 241.010 55.905 240.955 55.905 ;
        RECT 241.010 55.905 242.370 56.000 ;
        RECT 237.005 55.780 239.145 55.905 ;
        POLYGON 239.145 55.905 239.205 55.905 239.145 55.780 ;
        POLYGON 240.955 55.905 240.955 55.840 240.915 55.840 ;
        RECT 240.955 55.840 242.370 55.905 ;
        POLYGON 240.915 55.840 240.915 55.780 240.880 55.780 ;
        RECT 240.915 55.815 242.370 55.840 ;
        POLYGON 242.370 56.015 242.525 56.015 242.370 55.815 ;
        POLYGON 243.825 56.020 243.825 55.960 243.775 55.960 ;
        RECT 243.825 56.015 244.845 56.020 ;
        POLYGON 244.845 56.065 244.890 56.065 244.845 56.015 ;
        POLYGON 246.085 56.065 246.085 56.045 246.055 56.045 ;
        RECT 246.085 56.055 247.250 56.065 ;
        POLYGON 247.250 56.070 247.275 56.070 247.250 56.055 ;
        POLYGON 248.545 56.070 248.545 56.055 248.490 56.055 ;
        RECT 248.545 56.065 251.920 56.070 ;
        POLYGON 251.920 56.070 251.935 56.065 251.920 56.065 ;
        POLYGON 253.325 56.070 253.335 56.070 253.335 56.065 ;
        RECT 253.335 56.065 254.380 56.070 ;
        RECT 248.545 56.060 251.935 56.065 ;
        POLYGON 251.935 56.065 251.955 56.060 251.935 56.060 ;
        POLYGON 253.335 56.065 253.345 56.065 253.345 56.060 ;
        RECT 253.345 56.060 254.380 56.065 ;
        RECT 248.545 56.055 251.955 56.060 ;
        RECT 246.085 56.045 247.215 56.055 ;
        POLYGON 246.055 56.045 246.055 56.025 246.030 56.025 ;
        RECT 246.055 56.040 247.215 56.045 ;
        POLYGON 247.215 56.055 247.250 56.055 247.215 56.040 ;
        POLYGON 248.490 56.055 248.490 56.045 248.455 56.045 ;
        RECT 248.490 56.050 251.955 56.055 ;
        POLYGON 251.955 56.060 252.000 56.050 251.955 56.050 ;
        POLYGON 253.345 56.060 253.365 56.060 253.365 56.050 ;
        RECT 253.365 56.050 254.380 56.060 ;
        RECT 248.490 56.045 252.000 56.050 ;
        POLYGON 248.455 56.045 248.455 56.040 248.435 56.040 ;
        RECT 248.455 56.040 252.000 56.045 ;
        RECT 246.055 56.025 247.150 56.040 ;
        POLYGON 246.030 56.025 246.030 56.015 246.015 56.015 ;
        RECT 246.030 56.015 247.150 56.025 ;
        RECT 243.825 55.960 244.725 56.015 ;
        POLYGON 243.775 55.960 243.775 55.830 243.660 55.830 ;
        RECT 243.775 55.900 244.725 55.960 ;
        POLYGON 244.725 56.015 244.845 56.015 244.725 55.900 ;
        POLYGON 246.015 56.015 246.015 55.965 245.945 55.965 ;
        RECT 246.015 56.005 247.150 56.015 ;
        POLYGON 247.150 56.040 247.215 56.040 247.150 56.005 ;
        POLYGON 248.435 56.040 248.435 56.030 248.390 56.030 ;
        RECT 248.435 56.030 252.000 56.040 ;
        POLYGON 248.385 56.030 248.385 56.010 248.320 56.010 ;
        RECT 248.385 56.010 252.000 56.030 ;
        POLYGON 248.320 56.010 248.320 56.005 248.295 56.005 ;
        RECT 248.320 56.005 252.000 56.010 ;
        RECT 246.015 55.965 247.000 56.005 ;
        POLYGON 245.945 55.965 245.945 55.900 245.860 55.900 ;
        RECT 245.945 55.925 247.000 55.965 ;
        POLYGON 247.000 56.005 247.150 56.005 247.000 55.925 ;
        POLYGON 248.295 56.005 248.295 56.000 248.265 56.000 ;
        RECT 248.295 56.000 252.000 56.005 ;
        POLYGON 252.000 56.050 252.175 56.000 252.000 56.000 ;
        POLYGON 253.365 56.050 253.390 56.050 253.390 56.040 ;
        RECT 253.390 56.040 254.380 56.050 ;
        POLYGON 253.390 56.040 253.410 56.040 253.410 56.030 ;
        RECT 253.410 56.030 254.380 56.040 ;
        POLYGON 253.410 56.030 253.460 56.030 253.460 56.000 ;
        RECT 253.460 56.010 254.380 56.030 ;
        POLYGON 254.380 56.075 254.475 56.010 254.380 56.010 ;
        POLYGON 255.515 56.075 255.545 56.075 255.545 56.050 ;
        RECT 255.545 56.050 256.765 56.075 ;
        POLYGON 255.545 56.050 255.585 56.050 255.585 56.010 ;
        RECT 255.585 56.020 256.765 56.050 ;
        POLYGON 256.765 56.150 256.890 56.020 256.765 56.020 ;
        POLYGON 258.270 56.150 258.295 56.150 258.295 56.120 ;
        RECT 258.295 56.125 259.855 56.150 ;
        POLYGON 259.855 56.455 260.080 56.125 259.855 56.125 ;
        POLYGON 262.075 56.455 262.080 56.455 262.080 56.450 ;
        RECT 262.080 56.450 264.755 56.455 ;
        POLYGON 264.755 56.920 264.995 56.450 264.755 56.450 ;
        POLYGON 269.125 56.920 269.350 56.920 269.350 56.450 ;
        RECT 269.350 56.680 276.115 56.920 ;
        POLYGON 276.115 57.275 276.330 56.680 276.115 56.680 ;
        RECT 269.350 56.450 276.330 56.680 ;
        POLYGON 262.080 56.450 262.265 56.450 262.265 56.125 ;
        RECT 262.265 56.390 264.995 56.450 ;
        POLYGON 264.995 56.450 265.025 56.390 264.995 56.390 ;
        POLYGON 269.350 56.450 269.370 56.450 269.370 56.410 ;
        RECT 269.370 56.410 276.330 56.450 ;
        POLYGON 269.370 56.410 269.375 56.410 269.375 56.395 ;
        RECT 269.375 56.390 276.330 56.410 ;
        RECT 262.265 56.125 265.025 56.390 ;
        RECT 258.295 56.120 260.080 56.125 ;
        POLYGON 258.295 56.120 258.310 56.120 258.310 56.105 ;
        RECT 258.310 56.105 260.080 56.120 ;
        POLYGON 258.310 56.105 258.375 56.105 258.375 56.025 ;
        RECT 258.375 56.045 260.080 56.105 ;
        POLYGON 260.080 56.125 260.130 56.045 260.080 56.045 ;
        POLYGON 262.265 56.125 262.310 56.125 262.310 56.050 ;
        RECT 262.310 56.045 265.025 56.125 ;
        RECT 258.375 56.020 260.130 56.045 ;
        RECT 255.585 56.010 256.890 56.020 ;
        RECT 253.460 56.000 254.475 56.010 ;
        POLYGON 248.265 56.000 248.265 55.975 248.200 55.975 ;
        RECT 248.265 55.985 252.180 56.000 ;
        POLYGON 252.180 56.000 252.225 55.985 252.180 55.985 ;
        POLYGON 253.460 56.000 253.485 56.000 253.485 55.985 ;
        RECT 253.485 55.985 254.475 56.000 ;
        RECT 248.265 55.980 252.225 55.985 ;
        POLYGON 252.225 55.985 252.245 55.980 252.225 55.980 ;
        POLYGON 253.485 55.985 253.495 55.985 253.495 55.980 ;
        RECT 253.495 55.980 254.475 55.985 ;
        RECT 248.265 55.975 252.245 55.980 ;
        POLYGON 252.245 55.980 252.255 55.975 252.245 55.975 ;
        POLYGON 253.495 55.980 253.505 55.980 253.505 55.975 ;
        RECT 253.505 55.975 254.475 55.980 ;
        POLYGON 248.200 55.975 248.200 55.950 248.110 55.950 ;
        RECT 248.200 55.950 252.255 55.975 ;
        POLYGON 248.110 55.950 248.110 55.930 248.050 55.930 ;
        RECT 248.110 55.930 252.255 55.950 ;
        POLYGON 252.255 55.975 252.395 55.930 252.255 55.930 ;
        POLYGON 253.505 55.975 253.570 55.975 253.570 55.940 ;
        RECT 253.570 55.940 254.475 55.975 ;
        POLYGON 253.570 55.940 253.585 55.940 253.585 55.930 ;
        RECT 253.585 55.930 254.475 55.940 ;
        POLYGON 248.050 55.930 248.050 55.925 248.030 55.925 ;
        RECT 248.050 55.925 252.395 55.930 ;
        RECT 245.945 55.915 246.985 55.925 ;
        POLYGON 246.985 55.925 247.000 55.925 246.985 55.915 ;
        POLYGON 248.030 55.925 248.030 55.915 247.995 55.915 ;
        RECT 248.030 55.915 252.395 55.925 ;
        POLYGON 252.395 55.930 252.435 55.915 252.395 55.915 ;
        POLYGON 253.585 55.930 253.610 55.930 253.610 55.915 ;
        RECT 253.610 55.915 254.475 55.930 ;
        RECT 245.945 55.900 246.890 55.915 ;
        RECT 243.775 55.875 244.700 55.900 ;
        POLYGON 244.700 55.900 244.725 55.900 244.700 55.880 ;
        POLYGON 245.860 55.900 245.860 55.890 245.845 55.890 ;
        RECT 245.860 55.890 246.890 55.900 ;
        POLYGON 245.840 55.890 245.840 55.880 245.830 55.880 ;
        RECT 245.840 55.880 246.890 55.890 ;
        RECT 243.775 55.830 244.590 55.875 ;
        POLYGON 243.660 55.830 243.660 55.815 243.650 55.815 ;
        RECT 243.660 55.815 244.590 55.830 ;
        RECT 240.915 55.780 242.340 55.815 ;
        RECT 237.005 55.740 239.130 55.780 ;
        POLYGON 239.130 55.780 239.145 55.780 239.130 55.740 ;
        RECT 240.880 55.775 242.340 55.780 ;
        POLYGON 242.340 55.815 242.370 55.815 242.340 55.775 ;
        POLYGON 243.650 55.815 243.650 55.790 243.630 55.790 ;
        RECT 243.650 55.790 244.590 55.815 ;
        POLYGON 243.630 55.790 243.630 55.775 243.620 55.775 ;
        RECT 243.630 55.775 244.590 55.790 ;
        POLYGON 240.880 55.775 240.880 55.740 240.860 55.740 ;
        RECT 240.880 55.740 242.300 55.775 ;
        RECT 237.005 55.735 239.125 55.740 ;
        POLYGON 239.125 55.740 239.130 55.740 239.125 55.735 ;
        POLYGON 240.860 55.740 240.860 55.735 240.855 55.735 ;
        RECT 240.860 55.735 242.300 55.740 ;
        RECT 237.005 55.675 238.980 55.735 ;
        POLYGON 236.875 55.675 236.875 55.625 236.855 55.625 ;
        RECT 236.875 55.625 238.980 55.675 ;
        RECT 229.525 55.445 233.620 55.615 ;
        POLYGON 229.485 55.445 229.485 54.090 229.305 54.090 ;
        RECT 229.485 54.845 233.620 55.445 ;
        POLYGON 233.620 55.615 233.815 55.615 233.620 54.845 ;
        POLYGON 236.855 55.620 236.855 55.275 236.725 55.275 ;
        RECT 236.855 55.410 238.980 55.625 ;
        POLYGON 238.980 55.735 239.125 55.735 238.980 55.410 ;
        POLYGON 240.855 55.730 240.855 55.685 240.830 55.685 ;
        RECT 240.855 55.725 242.300 55.735 ;
        POLYGON 242.300 55.775 242.340 55.775 242.300 55.725 ;
        POLYGON 243.620 55.775 243.620 55.725 243.580 55.725 ;
        RECT 243.620 55.760 244.590 55.775 ;
        POLYGON 244.590 55.875 244.700 55.875 244.590 55.760 ;
        POLYGON 245.830 55.880 245.830 55.850 245.790 55.850 ;
        RECT 245.830 55.865 246.890 55.880 ;
        POLYGON 246.890 55.915 246.975 55.915 246.890 55.865 ;
        POLYGON 247.995 55.915 247.995 55.910 247.975 55.910 ;
        RECT 247.995 55.910 252.435 55.915 ;
        POLYGON 247.975 55.910 247.975 55.900 247.945 55.900 ;
        RECT 247.975 55.900 252.435 55.910 ;
        POLYGON 247.945 55.900 247.945 55.865 247.855 55.865 ;
        RECT 247.945 55.895 252.435 55.900 ;
        POLYGON 252.435 55.915 252.500 55.895 252.435 55.895 ;
        POLYGON 253.610 55.915 253.650 55.915 253.650 55.895 ;
        RECT 253.650 55.900 254.475 55.915 ;
        POLYGON 254.475 56.010 254.615 55.900 254.475 55.900 ;
        POLYGON 255.585 56.010 255.695 56.010 255.695 55.915 ;
        RECT 255.695 55.925 256.890 56.010 ;
        POLYGON 256.890 56.020 256.985 55.925 256.890 55.925 ;
        POLYGON 258.375 56.020 258.400 56.020 258.400 55.995 ;
        RECT 258.400 56.015 260.130 56.020 ;
        POLYGON 260.130 56.045 260.150 56.015 260.130 56.015 ;
        POLYGON 262.310 56.045 262.330 56.045 262.330 56.015 ;
        RECT 262.330 56.015 265.025 56.045 ;
        RECT 258.400 55.995 260.150 56.015 ;
        POLYGON 258.400 55.995 258.445 55.995 258.445 55.940 ;
        RECT 258.445 55.940 260.150 55.995 ;
        POLYGON 258.445 55.940 258.455 55.940 258.455 55.925 ;
        RECT 258.455 55.925 260.150 55.940 ;
        RECT 255.695 55.915 256.985 55.925 ;
        POLYGON 255.695 55.915 255.710 55.915 255.710 55.900 ;
        RECT 255.710 55.910 256.985 55.915 ;
        POLYGON 256.985 55.925 256.995 55.910 256.985 55.910 ;
        POLYGON 258.455 55.925 258.460 55.925 258.460 55.920 ;
        RECT 258.460 55.920 260.150 55.925 ;
        POLYGON 258.460 55.920 258.465 55.920 258.465 55.910 ;
        RECT 258.465 55.910 260.150 55.920 ;
        RECT 255.710 55.900 256.995 55.910 ;
        RECT 253.650 55.895 254.615 55.900 ;
        POLYGON 254.615 55.900 254.630 55.895 254.615 55.895 ;
        POLYGON 255.710 55.900 255.715 55.900 255.715 55.895 ;
        RECT 255.715 55.895 256.995 55.900 ;
        RECT 247.945 55.890 252.500 55.895 ;
        POLYGON 252.500 55.895 252.510 55.890 252.500 55.890 ;
        POLYGON 253.650 55.895 253.660 55.895 253.660 55.890 ;
        RECT 253.660 55.890 254.630 55.895 ;
        RECT 247.945 55.875 252.510 55.890 ;
        POLYGON 252.510 55.890 252.545 55.875 252.510 55.875 ;
        POLYGON 253.660 55.890 253.680 55.890 253.680 55.875 ;
        RECT 253.680 55.875 254.630 55.890 ;
        RECT 247.945 55.865 252.545 55.875 ;
        RECT 245.830 55.850 246.745 55.865 ;
        POLYGON 245.790 55.850 245.790 55.760 245.675 55.760 ;
        RECT 245.790 55.780 246.745 55.850 ;
        POLYGON 246.745 55.865 246.890 55.865 246.745 55.780 ;
        POLYGON 247.855 55.865 247.855 55.855 247.830 55.855 ;
        RECT 247.855 55.855 252.545 55.865 ;
        POLYGON 247.830 55.855 247.830 55.840 247.785 55.840 ;
        RECT 247.830 55.840 252.545 55.855 ;
        POLYGON 247.785 55.840 247.785 55.810 247.700 55.810 ;
        RECT 247.785 55.820 252.545 55.840 ;
        POLYGON 252.545 55.875 252.680 55.820 252.545 55.820 ;
        POLYGON 253.680 55.875 253.750 55.875 253.750 55.835 ;
        RECT 253.750 55.835 254.630 55.875 ;
        POLYGON 254.630 55.895 254.710 55.835 254.630 55.835 ;
        POLYGON 255.715 55.895 255.740 55.895 255.740 55.875 ;
        RECT 255.740 55.875 256.995 55.895 ;
        POLYGON 255.740 55.875 255.780 55.875 255.780 55.835 ;
        RECT 255.780 55.835 256.995 55.875 ;
        POLYGON 253.750 55.835 253.775 55.835 253.775 55.820 ;
        RECT 253.775 55.820 254.710 55.835 ;
        RECT 247.785 55.810 252.690 55.820 ;
        POLYGON 247.695 55.810 247.695 55.805 247.690 55.805 ;
        RECT 247.695 55.805 252.690 55.810 ;
        POLYGON 247.690 55.805 247.690 55.780 247.630 55.780 ;
        RECT 247.690 55.785 252.690 55.805 ;
        POLYGON 252.690 55.820 252.760 55.785 252.690 55.785 ;
        POLYGON 253.775 55.820 253.835 55.820 253.835 55.785 ;
        RECT 253.835 55.785 254.710 55.820 ;
        RECT 247.690 55.780 252.770 55.785 ;
        RECT 245.790 55.775 246.740 55.780 ;
        POLYGON 246.740 55.780 246.745 55.780 246.740 55.775 ;
        POLYGON 247.630 55.780 247.630 55.775 247.615 55.775 ;
        RECT 247.630 55.775 252.770 55.780 ;
        RECT 245.790 55.765 246.725 55.775 ;
        POLYGON 246.725 55.775 246.740 55.775 246.725 55.765 ;
        POLYGON 247.615 55.775 247.615 55.765 247.590 55.765 ;
        RECT 247.615 55.765 252.770 55.775 ;
        RECT 245.790 55.760 246.645 55.765 ;
        RECT 243.620 55.725 244.505 55.760 ;
        RECT 240.855 55.685 242.235 55.725 ;
        POLYGON 240.830 55.685 240.830 55.540 240.755 55.540 ;
        RECT 240.830 55.625 242.235 55.685 ;
        POLYGON 242.235 55.725 242.300 55.725 242.235 55.625 ;
        POLYGON 243.580 55.725 243.580 55.625 243.500 55.625 ;
        RECT 243.580 55.675 244.505 55.725 ;
        POLYGON 244.505 55.760 244.590 55.760 244.505 55.675 ;
        POLYGON 245.675 55.760 245.675 55.750 245.660 55.750 ;
        RECT 245.675 55.750 246.645 55.760 ;
        POLYGON 245.660 55.750 245.660 55.735 245.640 55.735 ;
        RECT 245.660 55.735 246.645 55.750 ;
        POLYGON 245.640 55.735 245.640 55.675 245.565 55.675 ;
        RECT 245.640 55.715 246.645 55.735 ;
        POLYGON 246.645 55.765 246.725 55.765 246.645 55.715 ;
        POLYGON 247.590 55.765 247.590 55.750 247.555 55.750 ;
        RECT 247.590 55.755 252.770 55.765 ;
        POLYGON 252.770 55.785 252.830 55.755 252.770 55.755 ;
        POLYGON 253.835 55.785 253.870 55.785 253.870 55.760 ;
        RECT 253.870 55.760 254.710 55.785 ;
        POLYGON 253.870 55.760 253.875 55.760 253.875 55.755 ;
        RECT 253.875 55.755 254.710 55.760 ;
        RECT 247.590 55.750 250.650 55.755 ;
        POLYGON 250.650 55.755 250.815 55.755 250.650 55.750 ;
        POLYGON 250.980 55.755 251.025 55.755 251.025 55.750 ;
        RECT 251.025 55.750 252.830 55.755 ;
        POLYGON 247.555 55.750 247.555 55.730 247.515 55.730 ;
        RECT 247.555 55.745 250.585 55.750 ;
        POLYGON 250.585 55.750 250.645 55.750 250.585 55.745 ;
        POLYGON 251.095 55.750 251.140 55.750 251.140 55.745 ;
        RECT 251.140 55.745 252.830 55.750 ;
        RECT 247.555 55.740 250.485 55.745 ;
        POLYGON 250.485 55.745 250.565 55.745 250.485 55.740 ;
        POLYGON 251.140 55.745 251.220 55.745 251.220 55.740 ;
        RECT 251.220 55.740 252.830 55.745 ;
        RECT 247.555 55.735 250.455 55.740 ;
        POLYGON 250.455 55.740 250.470 55.740 250.455 55.735 ;
        POLYGON 251.235 55.740 251.270 55.740 251.270 55.735 ;
        RECT 251.270 55.735 252.830 55.740 ;
        RECT 247.555 55.730 250.380 55.735 ;
        POLYGON 250.380 55.735 250.455 55.735 250.380 55.730 ;
        POLYGON 251.300 55.735 251.330 55.735 251.330 55.730 ;
        RECT 251.330 55.730 252.830 55.735 ;
        POLYGON 247.515 55.730 247.515 55.715 247.480 55.715 ;
        RECT 247.515 55.720 250.290 55.730 ;
        POLYGON 250.290 55.730 250.375 55.730 250.290 55.720 ;
        POLYGON 251.330 55.730 251.365 55.730 251.365 55.725 ;
        RECT 251.365 55.725 252.830 55.730 ;
        POLYGON 251.375 55.725 251.410 55.725 251.410 55.720 ;
        RECT 251.410 55.720 252.830 55.725 ;
        RECT 247.515 55.715 250.210 55.720 ;
        RECT 245.640 55.675 246.520 55.715 ;
        RECT 243.580 55.625 244.410 55.675 ;
        RECT 240.830 55.560 242.185 55.625 ;
        POLYGON 242.185 55.625 242.235 55.625 242.185 55.560 ;
        POLYGON 243.500 55.625 243.500 55.570 243.455 55.570 ;
        RECT 243.500 55.570 244.410 55.625 ;
        POLYGON 244.410 55.675 244.505 55.675 244.410 55.570 ;
        POLYGON 245.565 55.675 245.565 55.670 245.560 55.670 ;
        RECT 245.565 55.670 246.520 55.675 ;
        POLYGON 245.560 55.670 245.560 55.575 245.445 55.575 ;
        RECT 245.560 55.640 246.520 55.670 ;
        POLYGON 246.520 55.715 246.640 55.715 246.520 55.640 ;
        POLYGON 247.480 55.715 247.480 55.705 247.455 55.705 ;
        RECT 247.480 55.710 250.210 55.715 ;
        POLYGON 250.210 55.720 250.255 55.720 250.210 55.710 ;
        POLYGON 251.410 55.720 251.450 55.720 251.450 55.715 ;
        RECT 251.450 55.715 252.830 55.720 ;
        POLYGON 251.450 55.715 251.480 55.715 251.480 55.710 ;
        RECT 251.480 55.710 252.830 55.715 ;
        POLYGON 252.830 55.755 252.930 55.710 252.830 55.710 ;
        POLYGON 253.875 55.755 253.925 55.755 253.925 55.725 ;
        RECT 253.925 55.725 254.710 55.755 ;
        POLYGON 253.925 55.725 253.945 55.725 253.945 55.710 ;
        RECT 253.945 55.720 254.710 55.725 ;
        POLYGON 254.710 55.835 254.850 55.720 254.710 55.720 ;
        POLYGON 255.780 55.835 255.880 55.835 255.880 55.745 ;
        RECT 255.880 55.745 256.995 55.835 ;
        POLYGON 255.880 55.745 255.905 55.745 255.905 55.720 ;
        RECT 255.905 55.720 256.995 55.745 ;
        RECT 253.945 55.710 254.850 55.720 ;
        POLYGON 254.850 55.720 254.860 55.710 254.850 55.710 ;
        POLYGON 255.905 55.720 255.915 55.720 255.915 55.710 ;
        RECT 255.915 55.710 256.995 55.720 ;
        RECT 247.480 55.705 250.185 55.710 ;
        POLYGON 250.185 55.710 250.205 55.710 250.185 55.705 ;
        POLYGON 251.480 55.710 251.515 55.710 251.515 55.705 ;
        RECT 251.515 55.705 252.930 55.710 ;
        POLYGON 247.455 55.705 247.455 55.690 247.415 55.690 ;
        RECT 247.455 55.700 250.135 55.705 ;
        POLYGON 250.135 55.705 250.180 55.705 250.135 55.700 ;
        POLYGON 251.515 55.705 251.540 55.705 251.540 55.700 ;
        RECT 251.540 55.700 252.930 55.705 ;
        RECT 247.455 55.690 250.070 55.700 ;
        POLYGON 250.070 55.700 250.135 55.700 250.070 55.690 ;
        POLYGON 251.540 55.700 251.590 55.700 251.590 55.690 ;
        RECT 251.590 55.690 252.930 55.700 ;
        POLYGON 252.930 55.710 252.975 55.690 252.930 55.690 ;
        POLYGON 253.945 55.710 253.975 55.710 253.975 55.690 ;
        RECT 253.975 55.690 254.860 55.710 ;
        POLYGON 247.415 55.690 247.415 55.640 247.305 55.640 ;
        RECT 247.415 55.685 250.020 55.690 ;
        POLYGON 250.020 55.690 250.055 55.690 250.020 55.685 ;
        POLYGON 251.610 55.690 251.630 55.690 251.630 55.685 ;
        RECT 251.630 55.685 252.975 55.690 ;
        RECT 247.415 55.680 249.975 55.685 ;
        POLYGON 249.975 55.685 250.020 55.685 249.975 55.680 ;
        POLYGON 251.630 55.685 251.655 55.685 251.655 55.680 ;
        RECT 251.655 55.680 252.975 55.685 ;
        RECT 247.415 55.675 249.935 55.680 ;
        POLYGON 249.935 55.680 249.975 55.680 249.935 55.675 ;
        POLYGON 251.660 55.680 251.680 55.680 251.680 55.675 ;
        RECT 251.680 55.675 252.975 55.680 ;
        RECT 247.415 55.670 249.920 55.675 ;
        POLYGON 249.920 55.675 249.935 55.675 249.920 55.670 ;
        POLYGON 251.680 55.675 251.700 55.675 251.700 55.670 ;
        RECT 251.700 55.670 252.975 55.675 ;
        POLYGON 252.975 55.690 253.010 55.670 252.975 55.670 ;
        POLYGON 253.975 55.690 253.995 55.690 253.995 55.680 ;
        RECT 253.995 55.680 254.860 55.690 ;
        POLYGON 253.995 55.680 254.010 55.680 254.010 55.670 ;
        RECT 254.010 55.670 254.860 55.680 ;
        RECT 247.415 55.665 249.890 55.670 ;
        POLYGON 249.890 55.670 249.905 55.670 249.890 55.665 ;
        POLYGON 251.700 55.670 251.720 55.670 251.720 55.665 ;
        RECT 251.720 55.665 253.010 55.670 ;
        RECT 247.415 55.660 249.850 55.665 ;
        POLYGON 249.850 55.665 249.875 55.665 249.850 55.660 ;
        POLYGON 251.720 55.665 251.735 55.665 251.735 55.660 ;
        RECT 251.735 55.660 253.010 55.665 ;
        RECT 247.415 55.655 249.845 55.660 ;
        POLYGON 249.845 55.660 249.850 55.660 249.845 55.655 ;
        POLYGON 251.735 55.660 251.750 55.660 251.750 55.655 ;
        RECT 251.750 55.655 253.010 55.660 ;
        POLYGON 253.010 55.670 253.040 55.655 253.010 55.655 ;
        POLYGON 254.010 55.670 254.030 55.670 254.030 55.655 ;
        RECT 254.030 55.655 254.860 55.670 ;
        RECT 247.415 55.640 249.725 55.655 ;
        RECT 245.560 55.630 246.505 55.640 ;
        POLYGON 246.505 55.640 246.520 55.640 246.505 55.630 ;
        POLYGON 247.305 55.640 247.305 55.630 247.285 55.630 ;
        RECT 247.305 55.635 249.725 55.640 ;
        POLYGON 249.725 55.655 249.845 55.655 249.725 55.635 ;
        POLYGON 251.750 55.655 251.770 55.655 251.770 55.650 ;
        RECT 251.770 55.650 253.040 55.655 ;
        POLYGON 251.770 55.650 251.800 55.650 251.800 55.645 ;
        RECT 251.800 55.645 253.040 55.650 ;
        POLYGON 251.805 55.645 251.835 55.645 251.835 55.635 ;
        RECT 251.835 55.635 253.040 55.645 ;
        RECT 247.305 55.630 249.690 55.635 ;
        POLYGON 249.690 55.635 249.725 55.635 249.690 55.630 ;
        POLYGON 251.835 55.635 251.850 55.635 251.850 55.630 ;
        RECT 251.850 55.630 253.040 55.635 ;
        RECT 245.560 55.615 246.490 55.630 ;
        POLYGON 246.490 55.630 246.505 55.630 246.490 55.615 ;
        POLYGON 247.285 55.630 247.285 55.625 247.275 55.625 ;
        RECT 247.285 55.625 249.670 55.630 ;
        POLYGON 249.670 55.630 249.690 55.630 249.670 55.625 ;
        POLYGON 251.850 55.630 251.865 55.630 251.865 55.625 ;
        RECT 251.865 55.625 253.040 55.630 ;
        POLYGON 247.275 55.625 247.275 55.615 247.260 55.615 ;
        RECT 247.275 55.615 249.515 55.625 ;
        RECT 245.560 55.575 246.405 55.615 ;
        POLYGON 245.445 55.575 245.445 55.570 245.440 55.570 ;
        RECT 245.445 55.570 246.405 55.575 ;
        POLYGON 243.455 55.570 243.455 55.560 243.445 55.560 ;
        RECT 243.455 55.560 244.350 55.570 ;
        RECT 240.830 55.540 242.105 55.560 ;
        POLYGON 240.755 55.540 240.755 55.515 240.745 55.515 ;
        RECT 240.755 55.515 242.105 55.540 ;
        POLYGON 240.745 55.515 240.745 55.410 240.690 55.410 ;
        RECT 240.745 55.440 242.105 55.515 ;
        POLYGON 242.105 55.560 242.185 55.560 242.105 55.445 ;
        POLYGON 243.445 55.560 243.445 55.550 243.435 55.550 ;
        RECT 243.445 55.550 244.350 55.560 ;
        POLYGON 243.435 55.550 243.435 55.470 243.375 55.470 ;
        RECT 243.435 55.500 244.350 55.550 ;
        POLYGON 244.350 55.570 244.410 55.570 244.350 55.500 ;
        POLYGON 245.440 55.570 245.440 55.520 245.380 55.520 ;
        RECT 245.440 55.560 246.405 55.570 ;
        POLYGON 246.405 55.615 246.490 55.615 246.405 55.560 ;
        POLYGON 247.260 55.615 247.260 55.610 247.250 55.610 ;
        RECT 247.260 55.610 249.515 55.615 ;
        POLYGON 247.250 55.610 247.250 55.595 247.215 55.595 ;
        RECT 247.250 55.595 249.515 55.610 ;
        POLYGON 249.515 55.625 249.665 55.625 249.515 55.595 ;
        POLYGON 251.865 55.625 251.930 55.625 251.930 55.605 ;
        RECT 251.930 55.615 253.040 55.625 ;
        POLYGON 253.040 55.655 253.115 55.615 253.040 55.615 ;
        POLYGON 254.030 55.655 254.095 55.655 254.095 55.615 ;
        RECT 254.095 55.650 254.860 55.655 ;
        POLYGON 254.860 55.710 254.935 55.650 254.860 55.650 ;
        POLYGON 255.915 55.710 255.975 55.710 255.975 55.650 ;
        RECT 255.975 55.680 256.995 55.710 ;
        POLYGON 256.995 55.910 257.200 55.680 256.995 55.680 ;
        POLYGON 258.465 55.910 258.545 55.910 258.545 55.805 ;
        RECT 258.545 55.805 260.150 55.910 ;
        POLYGON 258.545 55.805 258.580 55.805 258.580 55.760 ;
        RECT 258.580 55.795 260.150 55.805 ;
        POLYGON 260.150 56.015 260.290 55.795 260.150 55.795 ;
        POLYGON 262.330 56.015 262.345 56.015 262.345 55.990 ;
        RECT 262.345 55.990 265.025 56.015 ;
        POLYGON 262.345 55.990 262.440 55.990 262.440 55.800 ;
        RECT 262.440 55.910 265.025 55.990 ;
        POLYGON 265.025 56.390 265.255 55.910 265.025 55.910 ;
        POLYGON 269.375 56.390 269.575 56.390 269.575 55.910 ;
        RECT 269.575 56.355 276.330 56.390 ;
        POLYGON 276.330 56.680 276.450 56.355 276.330 56.355 ;
        RECT 269.575 56.095 276.450 56.355 ;
        POLYGON 276.450 56.355 276.535 56.095 276.450 56.095 ;
        RECT 269.575 55.910 276.535 56.095 ;
        RECT 262.440 55.845 265.255 55.910 ;
        POLYGON 265.255 55.910 265.280 55.845 265.255 55.845 ;
        POLYGON 269.575 55.910 269.600 55.910 269.600 55.850 ;
        RECT 269.600 55.845 276.535 55.910 ;
        RECT 262.440 55.795 265.280 55.845 ;
        RECT 258.580 55.760 260.290 55.795 ;
        POLYGON 258.580 55.760 258.595 55.760 258.595 55.740 ;
        RECT 258.595 55.740 260.290 55.760 ;
        POLYGON 258.595 55.740 258.635 55.740 258.635 55.685 ;
        RECT 258.635 55.680 260.290 55.740 ;
        RECT 255.975 55.660 257.200 55.680 ;
        POLYGON 257.200 55.680 257.215 55.660 257.200 55.660 ;
        POLYGON 258.635 55.680 258.650 55.680 258.650 55.665 ;
        RECT 258.650 55.660 260.290 55.680 ;
        RECT 255.975 55.650 257.215 55.660 ;
        RECT 254.095 55.645 254.935 55.650 ;
        POLYGON 254.935 55.650 254.940 55.645 254.935 55.645 ;
        POLYGON 255.975 55.650 255.980 55.650 255.980 55.645 ;
        RECT 255.980 55.645 257.215 55.650 ;
        RECT 254.095 55.615 254.940 55.645 ;
        RECT 251.930 55.605 253.115 55.615 ;
        POLYGON 251.935 55.605 251.965 55.605 251.965 55.595 ;
        RECT 251.965 55.595 253.115 55.605 ;
        POLYGON 247.215 55.595 247.215 55.560 247.150 55.560 ;
        RECT 247.215 55.590 249.510 55.595 ;
        POLYGON 249.510 55.595 249.515 55.595 249.510 55.590 ;
        POLYGON 251.965 55.595 251.985 55.595 251.985 55.590 ;
        RECT 251.985 55.590 253.115 55.595 ;
        RECT 247.215 55.585 249.490 55.590 ;
        POLYGON 249.490 55.590 249.505 55.590 249.490 55.585 ;
        POLYGON 251.985 55.590 251.995 55.590 251.995 55.585 ;
        RECT 251.995 55.585 253.115 55.590 ;
        POLYGON 253.115 55.615 253.170 55.585 253.115 55.585 ;
        POLYGON 254.095 55.615 254.135 55.615 254.135 55.585 ;
        RECT 254.135 55.585 254.940 55.615 ;
        RECT 247.215 55.565 249.400 55.585 ;
        POLYGON 249.400 55.585 249.485 55.585 249.400 55.565 ;
        POLYGON 251.995 55.585 252.055 55.585 252.055 55.565 ;
        RECT 252.055 55.565 253.170 55.585 ;
        RECT 247.215 55.560 249.305 55.565 ;
        RECT 245.440 55.520 246.300 55.560 ;
        POLYGON 245.380 55.520 245.380 55.500 245.360 55.500 ;
        RECT 245.380 55.500 246.300 55.520 ;
        RECT 243.435 55.490 244.340 55.500 ;
        POLYGON 244.340 55.500 244.350 55.500 244.340 55.490 ;
        POLYGON 245.360 55.500 245.360 55.490 245.350 55.490 ;
        RECT 245.360 55.490 246.300 55.500 ;
        POLYGON 246.300 55.560 246.405 55.560 246.300 55.490 ;
        POLYGON 247.150 55.560 247.150 55.490 247.020 55.490 ;
        RECT 247.150 55.545 249.305 55.560 ;
        POLYGON 249.305 55.565 249.400 55.565 249.305 55.545 ;
        POLYGON 252.055 55.565 252.100 55.565 252.100 55.550 ;
        RECT 252.100 55.550 253.170 55.565 ;
        POLYGON 252.100 55.550 252.105 55.550 252.105 55.545 ;
        RECT 252.105 55.545 253.170 55.550 ;
        RECT 247.150 55.515 249.195 55.545 ;
        POLYGON 249.195 55.545 249.305 55.545 249.195 55.515 ;
        POLYGON 252.105 55.545 252.115 55.545 252.115 55.540 ;
        RECT 252.115 55.540 253.170 55.545 ;
        POLYGON 253.170 55.585 253.250 55.540 253.170 55.540 ;
        POLYGON 254.135 55.585 254.185 55.585 254.185 55.550 ;
        RECT 254.185 55.550 254.940 55.585 ;
        POLYGON 254.185 55.550 254.195 55.550 254.195 55.540 ;
        RECT 254.195 55.540 254.940 55.550 ;
        POLYGON 252.125 55.540 252.180 55.540 252.180 55.515 ;
        RECT 252.180 55.535 253.250 55.540 ;
        POLYGON 253.250 55.540 253.260 55.535 253.250 55.535 ;
        POLYGON 254.195 55.540 254.205 55.540 254.205 55.535 ;
        RECT 254.205 55.535 254.940 55.540 ;
        POLYGON 254.940 55.645 255.070 55.535 254.940 55.535 ;
        POLYGON 255.980 55.645 256.035 55.645 256.035 55.590 ;
        RECT 256.035 55.590 257.215 55.645 ;
        POLYGON 257.215 55.660 257.275 55.590 257.215 55.590 ;
        POLYGON 258.650 55.660 258.665 55.660 258.665 55.645 ;
        RECT 258.665 55.645 260.290 55.660 ;
        POLYGON 258.665 55.645 258.705 55.645 258.705 55.590 ;
        RECT 258.705 55.635 260.290 55.645 ;
        POLYGON 260.290 55.795 260.385 55.635 260.290 55.635 ;
        POLYGON 262.440 55.795 262.525 55.795 262.525 55.640 ;
        RECT 262.525 55.635 265.280 55.795 ;
        RECT 258.705 55.590 260.385 55.635 ;
        POLYGON 256.035 55.590 256.070 55.590 256.070 55.550 ;
        RECT 256.070 55.550 257.275 55.590 ;
        POLYGON 256.070 55.550 256.085 55.550 256.085 55.535 ;
        RECT 256.085 55.535 257.275 55.550 ;
        RECT 252.180 55.515 253.260 55.535 ;
        RECT 247.150 55.505 249.150 55.515 ;
        POLYGON 249.150 55.515 249.185 55.515 249.150 55.505 ;
        POLYGON 252.180 55.515 252.205 55.515 252.205 55.505 ;
        RECT 252.205 55.510 253.260 55.515 ;
        POLYGON 253.260 55.535 253.305 55.510 253.260 55.510 ;
        POLYGON 254.205 55.535 254.235 55.535 254.235 55.515 ;
        RECT 254.235 55.515 255.070 55.535 ;
        POLYGON 254.235 55.515 254.240 55.515 254.240 55.510 ;
        RECT 254.240 55.510 255.070 55.515 ;
        RECT 252.205 55.505 253.305 55.510 ;
        RECT 247.150 55.500 249.125 55.505 ;
        POLYGON 249.125 55.505 249.150 55.505 249.125 55.500 ;
        POLYGON 252.205 55.505 252.215 55.505 252.215 55.500 ;
        RECT 252.215 55.500 253.305 55.505 ;
        RECT 247.150 55.490 249.085 55.500 ;
        RECT 243.435 55.470 244.265 55.490 ;
        POLYGON 243.375 55.470 243.375 55.445 243.355 55.445 ;
        RECT 243.375 55.445 244.265 55.470 ;
        RECT 240.745 55.410 242.050 55.440 ;
        RECT 236.855 55.370 238.965 55.410 ;
        POLYGON 238.965 55.410 238.980 55.410 238.965 55.370 ;
        POLYGON 240.690 55.405 240.690 55.370 240.670 55.370 ;
        RECT 240.690 55.370 242.050 55.410 ;
        POLYGON 242.050 55.440 242.105 55.440 242.050 55.370 ;
        POLYGON 243.355 55.445 243.355 55.370 243.300 55.370 ;
        RECT 243.355 55.400 244.265 55.445 ;
        POLYGON 244.265 55.490 244.340 55.490 244.265 55.400 ;
        POLYGON 245.350 55.490 245.350 55.475 245.335 55.475 ;
        RECT 245.350 55.475 246.275 55.490 ;
        POLYGON 246.275 55.490 246.300 55.490 246.275 55.475 ;
        POLYGON 247.020 55.490 247.020 55.480 247.000 55.480 ;
        RECT 247.020 55.485 249.085 55.490 ;
        POLYGON 249.085 55.500 249.125 55.500 249.085 55.485 ;
        POLYGON 250.560 55.500 250.560 55.495 250.475 55.495 ;
        RECT 250.560 55.495 250.815 55.500 ;
        POLYGON 250.815 55.500 250.830 55.495 250.815 55.495 ;
        POLYGON 252.215 55.500 252.225 55.500 252.225 55.495 ;
        RECT 252.225 55.495 253.305 55.500 ;
        POLYGON 250.450 55.495 250.450 55.485 250.375 55.485 ;
        RECT 250.450 55.490 250.845 55.495 ;
        POLYGON 250.845 55.495 250.925 55.490 250.845 55.490 ;
        POLYGON 252.225 55.495 252.240 55.495 252.240 55.490 ;
        RECT 252.240 55.490 253.305 55.495 ;
        RECT 250.450 55.485 250.930 55.490 ;
        POLYGON 250.930 55.490 250.950 55.485 250.930 55.485 ;
        POLYGON 252.245 55.490 252.255 55.490 252.255 55.485 ;
        RECT 252.255 55.485 253.305 55.490 ;
        RECT 247.020 55.480 248.950 55.485 ;
        POLYGON 247.000 55.480 247.000 55.475 246.995 55.475 ;
        RECT 247.000 55.475 248.950 55.480 ;
        POLYGON 245.335 55.475 245.335 55.400 245.250 55.400 ;
        RECT 245.335 55.460 246.260 55.475 ;
        POLYGON 246.260 55.475 246.275 55.475 246.260 55.460 ;
        POLYGON 246.995 55.475 246.995 55.470 246.985 55.470 ;
        RECT 246.995 55.470 248.950 55.475 ;
        POLYGON 246.975 55.470 246.975 55.460 246.960 55.460 ;
        RECT 246.975 55.460 248.950 55.470 ;
        RECT 245.335 55.400 246.175 55.460 ;
        POLYGON 246.175 55.460 246.260 55.460 246.175 55.400 ;
        POLYGON 246.960 55.460 246.960 55.400 246.855 55.400 ;
        RECT 246.960 55.445 248.950 55.460 ;
        POLYGON 248.950 55.485 249.080 55.485 248.950 55.445 ;
        POLYGON 250.375 55.485 250.375 55.475 250.285 55.475 ;
        RECT 250.375 55.475 250.980 55.485 ;
        POLYGON 250.980 55.485 251.035 55.475 250.980 55.475 ;
        POLYGON 252.255 55.485 252.275 55.485 252.275 55.475 ;
        RECT 252.275 55.475 253.305 55.485 ;
        POLYGON 250.285 55.475 250.285 55.470 250.255 55.470 ;
        RECT 250.285 55.470 251.035 55.475 ;
        POLYGON 250.255 55.470 250.255 55.465 250.205 55.465 ;
        RECT 250.255 55.465 251.035 55.470 ;
        POLYGON 251.035 55.475 251.095 55.465 251.035 55.465 ;
        POLYGON 252.275 55.475 252.290 55.475 252.290 55.470 ;
        RECT 252.290 55.470 253.305 55.475 ;
        POLYGON 252.290 55.470 252.300 55.470 252.300 55.465 ;
        RECT 252.300 55.465 253.305 55.470 ;
        POLYGON 250.205 55.465 250.205 55.460 250.185 55.460 ;
        RECT 250.205 55.460 251.095 55.465 ;
        POLYGON 251.095 55.465 251.140 55.460 251.095 55.460 ;
        POLYGON 252.300 55.465 252.310 55.465 252.310 55.460 ;
        RECT 252.310 55.460 253.305 55.465 ;
        POLYGON 253.305 55.510 253.390 55.460 253.305 55.460 ;
        POLYGON 254.240 55.510 254.300 55.510 254.300 55.460 ;
        RECT 254.300 55.460 255.070 55.510 ;
        POLYGON 250.180 55.460 250.180 55.450 250.135 55.450 ;
        RECT 250.180 55.450 251.140 55.460 ;
        POLYGON 250.135 55.450 250.135 55.445 250.120 55.445 ;
        RECT 250.135 55.445 251.140 55.450 ;
        POLYGON 251.140 55.460 251.225 55.445 251.140 55.445 ;
        POLYGON 252.310 55.460 252.345 55.460 252.345 55.445 ;
        RECT 252.345 55.445 253.390 55.460 ;
        POLYGON 253.390 55.460 253.410 55.445 253.390 55.445 ;
        POLYGON 254.300 55.460 254.310 55.460 254.310 55.455 ;
        RECT 254.310 55.455 255.070 55.460 ;
        POLYGON 255.070 55.535 255.165 55.455 255.070 55.455 ;
        POLYGON 256.085 55.535 256.165 55.535 256.165 55.455 ;
        RECT 256.165 55.455 257.275 55.535 ;
        POLYGON 254.310 55.455 254.325 55.455 254.325 55.445 ;
        RECT 254.325 55.450 255.165 55.455 ;
        POLYGON 255.165 55.455 255.175 55.450 255.165 55.450 ;
        POLYGON 256.165 55.455 256.170 55.455 256.170 55.450 ;
        RECT 256.170 55.450 257.275 55.455 ;
        RECT 254.325 55.445 255.175 55.450 ;
        RECT 246.960 55.425 248.875 55.445 ;
        POLYGON 248.875 55.445 248.950 55.445 248.875 55.425 ;
        POLYGON 250.120 55.445 250.120 55.430 250.070 55.430 ;
        RECT 250.120 55.440 251.225 55.445 ;
        POLYGON 251.225 55.445 251.235 55.440 251.225 55.440 ;
        POLYGON 252.345 55.445 252.355 55.445 252.355 55.440 ;
        RECT 252.355 55.440 253.410 55.445 ;
        RECT 250.120 55.430 251.235 55.440 ;
        POLYGON 251.235 55.440 251.275 55.430 251.235 55.430 ;
        POLYGON 252.355 55.440 252.375 55.440 252.375 55.430 ;
        RECT 252.375 55.430 253.410 55.440 ;
        POLYGON 250.070 55.430 250.070 55.425 250.055 55.425 ;
        RECT 250.070 55.425 251.275 55.430 ;
        RECT 246.960 55.400 248.770 55.425 ;
        RECT 243.355 55.370 244.135 55.400 ;
        RECT 236.855 55.275 238.795 55.370 ;
        POLYGON 236.725 55.275 236.725 54.845 236.590 54.845 ;
        RECT 236.725 54.955 238.795 55.275 ;
        POLYGON 238.795 55.370 238.965 55.370 238.795 54.955 ;
        POLYGON 240.670 55.370 240.670 55.230 240.600 55.230 ;
        RECT 240.670 55.270 241.990 55.370 ;
        POLYGON 241.990 55.370 242.050 55.370 241.990 55.270 ;
        POLYGON 243.300 55.370 243.300 55.295 243.245 55.295 ;
        RECT 243.300 55.295 244.135 55.370 ;
        POLYGON 243.245 55.295 243.245 55.275 243.235 55.275 ;
        RECT 243.245 55.275 244.135 55.295 ;
        POLYGON 243.235 55.275 243.235 55.270 243.230 55.270 ;
        RECT 243.235 55.270 244.135 55.275 ;
        RECT 240.670 55.230 241.885 55.270 ;
        POLYGON 240.600 55.230 240.600 54.960 240.480 54.960 ;
        RECT 240.600 55.105 241.885 55.230 ;
        POLYGON 241.885 55.270 241.990 55.270 241.885 55.105 ;
        POLYGON 243.230 55.270 243.230 55.145 243.145 55.145 ;
        RECT 243.230 55.245 244.135 55.270 ;
        POLYGON 244.135 55.400 244.265 55.400 244.135 55.245 ;
        POLYGON 245.250 55.400 245.250 55.275 245.115 55.275 ;
        RECT 245.250 55.335 246.085 55.400 ;
        POLYGON 246.085 55.400 246.175 55.400 246.085 55.335 ;
        POLYGON 246.855 55.400 246.855 55.335 246.745 55.335 ;
        RECT 246.855 55.395 248.770 55.400 ;
        POLYGON 248.770 55.425 248.870 55.425 248.770 55.395 ;
        POLYGON 250.055 55.425 250.055 55.415 250.020 55.415 ;
        RECT 250.055 55.415 251.275 55.425 ;
        POLYGON 250.020 55.415 250.020 55.395 249.985 55.395 ;
        RECT 250.020 55.410 251.275 55.415 ;
        POLYGON 251.275 55.430 251.375 55.410 251.275 55.410 ;
        POLYGON 252.375 55.430 252.390 55.430 252.390 55.425 ;
        RECT 252.390 55.425 253.410 55.430 ;
        POLYGON 252.395 55.425 252.425 55.425 252.425 55.410 ;
        RECT 252.425 55.410 253.410 55.425 ;
        RECT 250.020 55.395 251.375 55.410 ;
        RECT 246.855 55.390 248.750 55.395 ;
        POLYGON 248.750 55.395 248.770 55.395 248.750 55.390 ;
        POLYGON 249.985 55.395 249.985 55.390 249.975 55.390 ;
        RECT 249.985 55.390 251.375 55.395 ;
        POLYGON 251.375 55.410 251.445 55.390 251.375 55.390 ;
        POLYGON 252.425 55.410 252.460 55.410 252.460 55.395 ;
        RECT 252.460 55.395 253.410 55.410 ;
        POLYGON 252.460 55.395 252.470 55.395 252.470 55.390 ;
        RECT 252.470 55.390 253.410 55.395 ;
        RECT 246.855 55.335 248.595 55.390 ;
        POLYGON 248.595 55.390 248.750 55.390 248.595 55.335 ;
        POLYGON 249.975 55.390 249.975 55.370 249.935 55.370 ;
        RECT 249.975 55.370 251.450 55.390 ;
        POLYGON 251.450 55.390 251.515 55.370 251.450 55.370 ;
        POLYGON 252.470 55.390 252.510 55.390 252.510 55.370 ;
        RECT 252.510 55.380 253.410 55.390 ;
        POLYGON 253.410 55.445 253.505 55.380 253.410 55.380 ;
        POLYGON 254.325 55.445 254.350 55.445 254.350 55.430 ;
        RECT 254.350 55.430 255.175 55.445 ;
        POLYGON 254.350 55.430 254.410 55.430 254.410 55.380 ;
        RECT 254.410 55.385 255.175 55.430 ;
        POLYGON 255.175 55.450 255.240 55.385 255.175 55.385 ;
        POLYGON 256.170 55.450 256.195 55.450 256.195 55.430 ;
        RECT 256.195 55.430 257.275 55.450 ;
        POLYGON 256.195 55.430 256.230 55.430 256.230 55.385 ;
        RECT 256.230 55.425 257.275 55.430 ;
        POLYGON 257.275 55.590 257.410 55.425 257.275 55.425 ;
        POLYGON 258.705 55.590 258.720 55.590 258.720 55.570 ;
        RECT 258.720 55.570 260.385 55.590 ;
        POLYGON 260.385 55.635 260.420 55.570 260.385 55.570 ;
        POLYGON 262.525 55.635 262.560 55.635 262.560 55.575 ;
        RECT 262.560 55.570 265.280 55.635 ;
        POLYGON 258.720 55.570 258.820 55.570 258.820 55.430 ;
        RECT 258.820 55.475 260.420 55.570 ;
        POLYGON 260.420 55.570 260.475 55.475 260.420 55.475 ;
        POLYGON 262.560 55.570 262.590 55.570 262.590 55.520 ;
        RECT 262.590 55.520 265.280 55.570 ;
        POLYGON 262.590 55.520 262.610 55.520 262.610 55.475 ;
        RECT 262.610 55.475 265.280 55.520 ;
        RECT 258.820 55.450 260.475 55.475 ;
        POLYGON 260.475 55.475 260.490 55.450 260.475 55.450 ;
        POLYGON 262.610 55.475 262.620 55.475 262.620 55.455 ;
        RECT 262.620 55.450 265.280 55.475 ;
        RECT 258.820 55.425 260.490 55.450 ;
        RECT 256.230 55.410 257.410 55.425 ;
        POLYGON 257.410 55.425 257.425 55.410 257.410 55.410 ;
        POLYGON 258.820 55.425 258.830 55.425 258.830 55.410 ;
        RECT 258.830 55.410 260.490 55.425 ;
        RECT 256.230 55.385 257.425 55.410 ;
        RECT 254.410 55.380 255.240 55.385 ;
        RECT 252.510 55.370 253.505 55.380 ;
        POLYGON 249.935 55.370 249.935 55.335 249.900 55.335 ;
        RECT 249.935 55.345 251.515 55.370 ;
        POLYGON 251.515 55.370 251.590 55.345 251.515 55.345 ;
        POLYGON 252.510 55.370 252.545 55.370 252.545 55.355 ;
        RECT 252.545 55.355 253.505 55.370 ;
        POLYGON 252.545 55.355 252.565 55.355 252.565 55.345 ;
        RECT 252.565 55.345 253.505 55.355 ;
        RECT 249.935 55.340 251.595 55.345 ;
        POLYGON 251.595 55.345 251.610 55.340 251.595 55.340 ;
        POLYGON 252.565 55.345 252.575 55.345 252.575 55.340 ;
        RECT 252.575 55.340 253.505 55.345 ;
        RECT 249.935 55.335 251.610 55.340 ;
        RECT 245.250 55.310 246.055 55.335 ;
        POLYGON 246.055 55.335 246.085 55.335 246.055 55.310 ;
        POLYGON 246.745 55.335 246.745 55.330 246.740 55.330 ;
        RECT 246.745 55.330 248.565 55.335 ;
        POLYGON 246.740 55.330 246.740 55.310 246.710 55.310 ;
        RECT 246.740 55.325 248.565 55.330 ;
        POLYGON 248.565 55.335 248.595 55.335 248.565 55.325 ;
        POLYGON 249.900 55.335 249.900 55.325 249.895 55.325 ;
        RECT 249.900 55.325 251.610 55.335 ;
        POLYGON 251.610 55.340 251.660 55.325 251.610 55.325 ;
        POLYGON 252.575 55.340 252.605 55.340 252.605 55.325 ;
        RECT 252.605 55.335 253.505 55.340 ;
        POLYGON 253.505 55.380 253.570 55.335 253.505 55.335 ;
        POLYGON 254.410 55.380 254.445 55.380 254.445 55.355 ;
        RECT 254.445 55.355 255.240 55.380 ;
        POLYGON 254.445 55.355 254.475 55.355 254.475 55.335 ;
        RECT 254.475 55.345 255.240 55.355 ;
        POLYGON 255.240 55.385 255.290 55.345 255.240 55.345 ;
        POLYGON 256.230 55.385 256.270 55.385 256.270 55.345 ;
        RECT 256.270 55.345 257.425 55.385 ;
        RECT 254.475 55.335 255.290 55.345 ;
        RECT 252.605 55.325 253.570 55.335 ;
        RECT 246.740 55.320 248.545 55.325 ;
        POLYGON 248.545 55.325 248.565 55.325 248.545 55.320 ;
        POLYGON 249.895 55.325 249.895 55.320 249.890 55.320 ;
        RECT 249.895 55.320 251.660 55.325 ;
        RECT 246.740 55.310 248.470 55.320 ;
        RECT 245.250 55.295 246.035 55.310 ;
        POLYGON 246.035 55.310 246.055 55.310 246.035 55.295 ;
        POLYGON 246.710 55.310 246.710 55.295 246.685 55.295 ;
        RECT 246.710 55.295 248.470 55.310 ;
        RECT 245.250 55.275 245.955 55.295 ;
        POLYGON 245.115 55.275 245.115 55.265 245.110 55.265 ;
        RECT 245.115 55.265 245.955 55.275 ;
        POLYGON 245.110 55.265 245.110 55.245 245.085 55.245 ;
        RECT 245.110 55.245 245.955 55.265 ;
        RECT 243.230 55.235 244.130 55.245 ;
        POLYGON 244.130 55.245 244.135 55.245 244.130 55.235 ;
        POLYGON 245.085 55.245 245.085 55.235 245.070 55.235 ;
        RECT 245.085 55.235 245.955 55.245 ;
        RECT 243.230 55.200 244.100 55.235 ;
        POLYGON 244.100 55.235 244.130 55.235 244.100 55.200 ;
        POLYGON 245.070 55.235 245.070 55.200 245.035 55.200 ;
        RECT 245.070 55.230 245.955 55.235 ;
        POLYGON 245.955 55.295 246.035 55.295 245.955 55.230 ;
        POLYGON 246.685 55.295 246.685 55.270 246.645 55.270 ;
        RECT 246.685 55.290 248.470 55.295 ;
        POLYGON 248.470 55.320 248.545 55.320 248.470 55.290 ;
        POLYGON 249.890 55.320 249.890 55.305 249.880 55.305 ;
        RECT 249.890 55.305 251.660 55.320 ;
        RECT 249.880 55.300 251.660 55.305 ;
        POLYGON 251.660 55.325 251.720 55.300 251.660 55.300 ;
        POLYGON 252.605 55.325 252.625 55.325 252.625 55.315 ;
        RECT 252.625 55.315 253.570 55.325 ;
        POLYGON 252.625 55.315 252.650 55.315 252.650 55.300 ;
        RECT 252.650 55.300 253.570 55.315 ;
        POLYGON 249.880 55.300 249.880 55.290 249.875 55.290 ;
        RECT 249.880 55.290 251.720 55.300 ;
        RECT 246.685 55.275 248.425 55.290 ;
        POLYGON 248.425 55.290 248.470 55.290 248.425 55.275 ;
        RECT 249.875 55.285 251.720 55.290 ;
        POLYGON 251.720 55.300 251.770 55.285 251.720 55.285 ;
        POLYGON 252.650 55.300 252.680 55.300 252.680 55.285 ;
        RECT 252.680 55.290 253.570 55.300 ;
        POLYGON 253.570 55.335 253.640 55.290 253.570 55.290 ;
        POLYGON 254.475 55.335 254.525 55.335 254.525 55.295 ;
        RECT 254.525 55.295 255.290 55.335 ;
        POLYGON 254.525 55.295 254.530 55.295 254.530 55.290 ;
        RECT 254.530 55.290 255.290 55.295 ;
        RECT 252.680 55.285 253.640 55.290 ;
        RECT 246.685 55.270 248.340 55.275 ;
        POLYGON 246.640 55.270 246.640 55.230 246.585 55.230 ;
        RECT 246.640 55.240 248.340 55.270 ;
        POLYGON 248.340 55.275 248.425 55.275 248.340 55.240 ;
        RECT 249.875 55.270 251.775 55.285 ;
        POLYGON 251.775 55.285 251.805 55.270 251.775 55.270 ;
        POLYGON 252.680 55.285 252.690 55.285 252.690 55.280 ;
        RECT 252.690 55.280 253.640 55.285 ;
        POLYGON 253.640 55.290 253.660 55.280 253.640 55.280 ;
        POLYGON 254.530 55.290 254.540 55.290 254.540 55.280 ;
        RECT 254.540 55.280 255.290 55.290 ;
        POLYGON 252.695 55.280 252.710 55.280 252.710 55.270 ;
        RECT 252.710 55.270 253.660 55.280 ;
        RECT 249.875 55.255 251.805 55.270 ;
        POLYGON 251.805 55.270 251.850 55.255 251.805 55.255 ;
        POLYGON 252.710 55.270 252.735 55.270 252.735 55.255 ;
        RECT 252.735 55.255 253.660 55.270 ;
        RECT 249.875 55.240 251.850 55.255 ;
        RECT 246.640 55.230 248.265 55.240 ;
        RECT 245.070 55.200 245.880 55.230 ;
        RECT 243.230 55.145 244.015 55.200 ;
        POLYGON 243.145 55.145 243.145 55.105 243.115 55.105 ;
        RECT 243.145 55.105 244.015 55.145 ;
        RECT 240.600 55.100 241.880 55.105 ;
        POLYGON 241.880 55.105 241.885 55.105 241.880 55.100 ;
        POLYGON 243.115 55.105 243.115 55.100 243.110 55.100 ;
        RECT 243.115 55.100 244.015 55.105 ;
        RECT 240.600 55.075 241.865 55.100 ;
        POLYGON 241.865 55.100 241.880 55.100 241.865 55.075 ;
        POLYGON 243.110 55.100 243.110 55.085 243.100 55.085 ;
        RECT 243.110 55.090 244.015 55.100 ;
        POLYGON 244.015 55.200 244.100 55.200 244.015 55.090 ;
        POLYGON 245.035 55.200 245.035 55.090 244.935 55.090 ;
        RECT 245.035 55.170 245.880 55.200 ;
        POLYGON 245.880 55.230 245.955 55.230 245.880 55.170 ;
        POLYGON 246.585 55.230 246.585 55.185 246.520 55.185 ;
        RECT 246.585 55.210 248.265 55.230 ;
        POLYGON 248.265 55.240 248.340 55.240 248.265 55.210 ;
        POLYGON 249.875 55.240 249.880 55.240 249.880 55.235 ;
        RECT 249.880 55.230 251.850 55.240 ;
        POLYGON 249.880 55.230 249.890 55.230 249.890 55.210 ;
        RECT 249.890 55.220 251.850 55.230 ;
        POLYGON 251.850 55.255 251.935 55.220 251.850 55.220 ;
        POLYGON 252.735 55.255 252.785 55.255 252.785 55.225 ;
        RECT 252.785 55.225 253.660 55.255 ;
        POLYGON 252.785 55.225 252.790 55.225 252.790 55.220 ;
        RECT 252.790 55.220 253.660 55.225 ;
        RECT 249.890 55.210 251.935 55.220 ;
        POLYGON 251.935 55.220 251.950 55.210 251.935 55.210 ;
        POLYGON 252.790 55.220 252.810 55.220 252.810 55.210 ;
        RECT 252.810 55.210 253.660 55.220 ;
        POLYGON 253.660 55.280 253.750 55.210 253.660 55.210 ;
        POLYGON 254.540 55.280 254.545 55.280 254.545 55.275 ;
        RECT 254.545 55.275 255.290 55.280 ;
        POLYGON 254.545 55.275 254.625 55.275 254.625 55.210 ;
        RECT 254.625 55.210 255.290 55.275 ;
        RECT 246.585 55.200 248.250 55.210 ;
        POLYGON 248.250 55.210 248.265 55.210 248.250 55.200 ;
        POLYGON 249.890 55.210 249.895 55.210 249.895 55.200 ;
        RECT 249.895 55.200 251.950 55.210 ;
        POLYGON 251.950 55.210 251.985 55.200 251.950 55.200 ;
        POLYGON 252.810 55.210 252.830 55.210 252.830 55.200 ;
        RECT 252.830 55.200 253.750 55.210 ;
        RECT 246.585 55.185 248.180 55.200 ;
        POLYGON 246.520 55.185 246.520 55.175 246.505 55.175 ;
        RECT 246.520 55.175 248.180 55.185 ;
        POLYGON 246.505 55.175 246.505 55.170 246.500 55.170 ;
        RECT 246.505 55.170 248.180 55.175 ;
        POLYGON 248.180 55.200 248.250 55.200 248.180 55.170 ;
        POLYGON 249.895 55.200 249.910 55.200 249.910 55.180 ;
        RECT 249.910 55.180 251.985 55.200 ;
        POLYGON 249.910 55.180 249.915 55.180 249.915 55.170 ;
        RECT 249.915 55.170 251.985 55.180 ;
        RECT 245.035 55.140 245.845 55.170 ;
        POLYGON 245.845 55.170 245.880 55.170 245.845 55.140 ;
        POLYGON 246.500 55.170 246.500 55.165 246.490 55.165 ;
        RECT 246.500 55.165 248.135 55.170 ;
        POLYGON 246.490 55.165 246.490 55.140 246.455 55.140 ;
        RECT 246.490 55.150 248.135 55.165 ;
        POLYGON 248.135 55.170 248.180 55.170 248.135 55.150 ;
        POLYGON 249.915 55.170 249.935 55.170 249.935 55.150 ;
        RECT 249.935 55.150 251.985 55.170 ;
        POLYGON 251.985 55.200 252.100 55.150 251.985 55.150 ;
        POLYGON 252.830 55.200 252.920 55.200 252.920 55.150 ;
        RECT 252.920 55.150 253.750 55.200 ;
        RECT 246.490 55.140 248.085 55.150 ;
        RECT 245.035 55.120 245.820 55.140 ;
        POLYGON 245.820 55.140 245.845 55.140 245.820 55.120 ;
        POLYGON 246.455 55.140 246.455 55.120 246.425 55.120 ;
        RECT 246.455 55.125 248.085 55.140 ;
        POLYGON 248.085 55.150 248.135 55.150 248.085 55.125 ;
        POLYGON 249.935 55.150 249.960 55.150 249.960 55.125 ;
        RECT 249.960 55.140 252.100 55.150 ;
        POLYGON 252.100 55.150 252.115 55.140 252.100 55.140 ;
        POLYGON 252.920 55.150 252.940 55.150 252.940 55.140 ;
        RECT 252.940 55.145 253.750 55.150 ;
        POLYGON 253.750 55.210 253.835 55.145 253.750 55.145 ;
        POLYGON 254.625 55.210 254.705 55.210 254.705 55.145 ;
        RECT 254.705 55.185 255.290 55.210 ;
        POLYGON 255.290 55.345 255.460 55.185 255.290 55.185 ;
        POLYGON 256.270 55.345 256.280 55.345 256.280 55.335 ;
        RECT 256.280 55.335 257.425 55.345 ;
        POLYGON 256.280 55.335 256.410 55.335 256.410 55.190 ;
        RECT 256.410 55.275 257.425 55.335 ;
        POLYGON 257.425 55.410 257.530 55.275 257.425 55.275 ;
        POLYGON 258.830 55.410 258.920 55.410 258.920 55.285 ;
        RECT 258.920 55.285 260.490 55.410 ;
        POLYGON 258.920 55.285 258.925 55.285 258.925 55.280 ;
        RECT 258.925 55.275 260.490 55.285 ;
        RECT 256.410 55.185 257.530 55.275 ;
        RECT 254.705 55.150 255.460 55.185 ;
        POLYGON 255.460 55.185 255.495 55.150 255.460 55.150 ;
        POLYGON 256.410 55.185 256.445 55.185 256.445 55.150 ;
        RECT 256.445 55.170 257.530 55.185 ;
        POLYGON 257.530 55.275 257.610 55.170 257.530 55.170 ;
        POLYGON 258.925 55.275 258.935 55.275 258.935 55.260 ;
        RECT 258.935 55.260 260.490 55.275 ;
        POLYGON 258.935 55.260 258.990 55.260 258.990 55.175 ;
        RECT 258.990 55.170 260.490 55.260 ;
        RECT 256.445 55.165 257.610 55.170 ;
        POLYGON 257.610 55.170 257.615 55.165 257.610 55.165 ;
        POLYGON 258.990 55.170 258.995 55.170 258.995 55.165 ;
        RECT 258.995 55.165 260.490 55.170 ;
        RECT 256.445 55.150 257.615 55.165 ;
        POLYGON 257.615 55.165 257.625 55.150 257.615 55.150 ;
        POLYGON 258.995 55.165 259.005 55.165 259.005 55.150 ;
        RECT 259.005 55.150 260.490 55.165 ;
        RECT 254.705 55.145 255.495 55.150 ;
        RECT 252.940 55.140 253.835 55.145 ;
        RECT 249.960 55.125 252.125 55.140 ;
        RECT 246.455 55.120 247.975 55.125 ;
        RECT 245.035 55.090 245.750 55.120 ;
        RECT 243.110 55.085 244.000 55.090 ;
        POLYGON 243.100 55.085 243.100 55.080 243.095 55.080 ;
        RECT 243.100 55.080 244.000 55.085 ;
        RECT 240.600 55.010 241.825 55.075 ;
        POLYGON 241.825 55.075 241.865 55.075 241.825 55.010 ;
        POLYGON 243.095 55.075 243.095 55.010 243.050 55.010 ;
        RECT 243.095 55.065 244.000 55.080 ;
        POLYGON 244.000 55.090 244.015 55.090 244.000 55.065 ;
        POLYGON 244.935 55.090 244.935 55.065 244.910 55.065 ;
        RECT 244.935 55.065 245.750 55.090 ;
        RECT 243.095 55.020 243.960 55.065 ;
        POLYGON 243.960 55.065 244.000 55.065 243.960 55.020 ;
        POLYGON 244.910 55.065 244.910 55.060 244.905 55.060 ;
        RECT 244.910 55.060 245.750 55.065 ;
        POLYGON 245.750 55.120 245.820 55.120 245.750 55.060 ;
        POLYGON 246.425 55.120 246.425 55.060 246.345 55.060 ;
        RECT 246.425 55.075 247.975 55.120 ;
        POLYGON 247.975 55.125 248.085 55.125 247.975 55.075 ;
        POLYGON 249.960 55.125 249.975 55.125 249.975 55.115 ;
        RECT 249.975 55.115 252.125 55.125 ;
        POLYGON 249.975 55.115 249.980 55.115 249.980 55.110 ;
        RECT 249.980 55.110 252.125 55.115 ;
        POLYGON 249.980 55.110 250.020 55.110 250.020 55.085 ;
        RECT 250.020 55.085 252.125 55.110 ;
        POLYGON 250.020 55.085 250.025 55.085 250.025 55.075 ;
        RECT 250.025 55.080 252.125 55.085 ;
        POLYGON 252.125 55.140 252.245 55.080 252.125 55.080 ;
        POLYGON 252.940 55.140 252.955 55.140 252.955 55.130 ;
        RECT 252.955 55.130 253.835 55.140 ;
        POLYGON 252.955 55.130 252.975 55.130 252.975 55.120 ;
        RECT 252.975 55.120 253.835 55.130 ;
        POLYGON 253.835 55.145 253.870 55.120 253.835 55.120 ;
        POLYGON 254.705 55.145 254.730 55.145 254.730 55.120 ;
        RECT 254.730 55.120 255.495 55.145 ;
        POLYGON 252.975 55.120 252.985 55.120 252.985 55.110 ;
        RECT 252.985 55.110 253.870 55.120 ;
        POLYGON 252.985 55.110 253.035 55.110 253.035 55.080 ;
        RECT 253.035 55.080 253.870 55.110 ;
        POLYGON 253.870 55.120 253.925 55.080 253.870 55.080 ;
        POLYGON 254.730 55.120 254.775 55.120 254.775 55.080 ;
        RECT 254.775 55.095 255.495 55.120 ;
        POLYGON 255.495 55.150 255.545 55.095 255.495 55.095 ;
        POLYGON 256.445 55.150 256.485 55.150 256.485 55.105 ;
        RECT 256.485 55.105 257.625 55.150 ;
        POLYGON 256.485 55.105 256.495 55.105 256.495 55.095 ;
        RECT 256.495 55.095 257.625 55.105 ;
        RECT 254.775 55.080 255.545 55.095 ;
        RECT 250.025 55.075 252.245 55.080 ;
        RECT 246.425 55.060 247.915 55.075 ;
        POLYGON 244.905 55.060 244.905 55.050 244.890 55.050 ;
        RECT 244.905 55.050 245.675 55.060 ;
        POLYGON 244.890 55.050 244.890 55.020 244.865 55.020 ;
        RECT 244.890 55.020 245.675 55.050 ;
        RECT 243.095 55.010 243.875 55.020 ;
        RECT 240.600 54.960 241.790 55.010 ;
        RECT 240.480 54.955 241.790 54.960 ;
        POLYGON 241.790 55.010 241.825 55.010 241.790 54.955 ;
        POLYGON 243.050 55.010 243.050 54.995 243.040 54.995 ;
        RECT 243.050 54.995 243.875 55.010 ;
        POLYGON 243.040 54.995 243.040 54.955 243.015 54.955 ;
        RECT 243.040 54.955 243.875 54.995 ;
        RECT 236.725 54.905 238.775 54.955 ;
        POLYGON 238.775 54.955 238.795 54.955 238.775 54.905 ;
        POLYGON 240.480 54.955 240.480 54.905 240.455 54.905 ;
        RECT 240.480 54.905 241.710 54.955 ;
        RECT 236.725 54.845 238.640 54.905 ;
        RECT 229.485 54.755 233.600 54.845 ;
        POLYGON 233.600 54.845 233.620 54.845 233.600 54.755 ;
        POLYGON 236.590 54.840 236.590 54.790 236.575 54.790 ;
        RECT 236.590 54.790 238.640 54.845 ;
        POLYGON 236.575 54.790 236.575 54.760 236.565 54.760 ;
        RECT 236.575 54.760 238.640 54.790 ;
        RECT 229.485 54.695 233.590 54.755 ;
        POLYGON 233.590 54.755 233.600 54.755 233.590 54.695 ;
        POLYGON 236.565 54.755 236.565 54.695 236.545 54.695 ;
        RECT 236.565 54.695 238.640 54.760 ;
        RECT 229.485 54.105 233.475 54.695 ;
        POLYGON 233.475 54.695 233.590 54.695 233.475 54.105 ;
        POLYGON 236.545 54.695 236.545 54.505 236.485 54.505 ;
        RECT 236.545 54.530 238.640 54.695 ;
        POLYGON 238.640 54.905 238.775 54.905 238.640 54.530 ;
        POLYGON 240.455 54.905 240.455 54.605 240.335 54.605 ;
        RECT 240.455 54.815 241.710 54.905 ;
        POLYGON 241.710 54.955 241.790 54.955 241.710 54.815 ;
        POLYGON 243.015 54.955 243.015 54.815 242.925 54.815 ;
        RECT 243.015 54.900 243.875 54.955 ;
        POLYGON 243.875 55.020 243.960 55.020 243.875 54.900 ;
        POLYGON 244.865 55.020 244.865 54.995 244.845 54.995 ;
        RECT 244.865 55.000 245.675 55.020 ;
        POLYGON 245.675 55.060 245.750 55.060 245.675 55.000 ;
        POLYGON 246.345 55.060 246.345 55.025 246.300 55.025 ;
        RECT 246.345 55.045 247.915 55.060 ;
        POLYGON 247.915 55.075 247.975 55.075 247.915 55.045 ;
        POLYGON 250.025 55.075 250.055 55.075 250.055 55.060 ;
        RECT 250.055 55.060 252.245 55.075 ;
        POLYGON 250.055 55.060 250.070 55.060 250.070 55.050 ;
        RECT 250.070 55.055 252.245 55.060 ;
        POLYGON 252.245 55.080 252.290 55.055 252.245 55.055 ;
        POLYGON 253.035 55.080 253.075 55.080 253.075 55.055 ;
        RECT 253.075 55.055 253.925 55.080 ;
        RECT 250.070 55.050 252.295 55.055 ;
        POLYGON 250.070 55.050 250.080 55.050 250.080 55.045 ;
        RECT 250.080 55.045 252.295 55.050 ;
        RECT 246.345 55.030 247.890 55.045 ;
        POLYGON 247.890 55.045 247.915 55.045 247.890 55.030 ;
        POLYGON 250.080 55.045 250.105 55.045 250.105 55.030 ;
        RECT 250.105 55.030 252.295 55.045 ;
        RECT 246.345 55.025 247.750 55.030 ;
        POLYGON 246.300 55.025 246.300 55.010 246.275 55.010 ;
        RECT 246.300 55.010 247.750 55.025 ;
        POLYGON 246.275 55.010 246.275 55.000 246.265 55.000 ;
        RECT 246.275 55.000 247.750 55.010 ;
        RECT 244.865 54.995 245.615 55.000 ;
        POLYGON 244.845 54.995 244.845 54.900 244.755 54.900 ;
        RECT 244.845 54.940 245.615 54.995 ;
        POLYGON 245.615 55.000 245.675 55.000 245.615 54.940 ;
        POLYGON 246.265 55.000 246.265 54.995 246.260 54.995 ;
        RECT 246.265 54.995 247.750 55.000 ;
        POLYGON 246.260 54.995 246.260 54.940 246.190 54.940 ;
        RECT 246.260 54.955 247.750 54.995 ;
        POLYGON 247.750 55.030 247.890 55.030 247.750 54.955 ;
        POLYGON 250.105 55.030 250.135 55.030 250.135 55.015 ;
        RECT 250.135 55.015 252.295 55.030 ;
        POLYGON 250.135 55.015 250.140 55.015 250.140 55.010 ;
        RECT 250.140 55.010 252.295 55.015 ;
        POLYGON 250.140 55.010 250.205 55.010 250.205 54.980 ;
        RECT 250.205 55.005 252.295 55.010 ;
        POLYGON 252.295 55.055 252.395 55.005 252.295 55.005 ;
        POLYGON 253.075 55.055 253.095 55.055 253.095 55.045 ;
        RECT 253.095 55.045 253.925 55.055 ;
        POLYGON 253.095 55.045 253.115 55.045 253.115 55.030 ;
        RECT 253.115 55.030 253.925 55.045 ;
        POLYGON 253.115 55.030 253.150 55.030 253.150 55.005 ;
        RECT 253.150 55.020 253.925 55.030 ;
        POLYGON 253.925 55.080 253.995 55.020 253.925 55.020 ;
        POLYGON 254.775 55.080 254.840 55.080 254.840 55.020 ;
        RECT 254.840 55.020 255.545 55.080 ;
        RECT 253.150 55.005 253.995 55.020 ;
        RECT 250.205 54.980 252.395 55.005 ;
        POLYGON 250.210 54.980 250.255 54.980 250.255 54.960 ;
        RECT 250.255 54.970 252.395 54.980 ;
        POLYGON 252.395 55.005 252.460 54.970 252.395 54.970 ;
        POLYGON 253.150 55.005 253.205 55.005 253.205 54.970 ;
        RECT 253.205 54.970 253.995 55.005 ;
        RECT 250.255 54.960 252.460 54.970 ;
        POLYGON 250.255 54.960 250.270 54.960 250.270 54.955 ;
        RECT 250.270 54.955 252.460 54.960 ;
        RECT 246.260 54.950 247.740 54.955 ;
        POLYGON 247.740 54.955 247.750 54.955 247.740 54.950 ;
        POLYGON 250.270 54.955 250.285 54.955 250.285 54.950 ;
        RECT 246.260 54.940 247.590 54.950 ;
        RECT 244.845 54.900 245.550 54.940 ;
        RECT 243.015 54.890 243.870 54.900 ;
        POLYGON 243.870 54.900 243.875 54.900 243.870 54.890 ;
        POLYGON 244.755 54.900 244.755 54.890 244.750 54.890 ;
        RECT 244.755 54.890 245.550 54.900 ;
        RECT 243.015 54.815 243.795 54.890 ;
        RECT 240.455 54.740 241.670 54.815 ;
        POLYGON 241.670 54.815 241.710 54.815 241.670 54.740 ;
        POLYGON 242.925 54.810 242.925 54.740 242.880 54.740 ;
        RECT 242.925 54.790 243.795 54.815 ;
        POLYGON 243.795 54.890 243.870 54.890 243.795 54.790 ;
        POLYGON 244.750 54.890 244.750 54.840 244.700 54.840 ;
        RECT 244.750 54.885 245.550 54.890 ;
        POLYGON 245.550 54.940 245.615 54.940 245.550 54.885 ;
        POLYGON 246.190 54.940 246.190 54.930 246.175 54.930 ;
        RECT 246.190 54.930 247.590 54.940 ;
        POLYGON 246.175 54.930 246.175 54.885 246.120 54.885 ;
        RECT 246.175 54.885 247.590 54.930 ;
        RECT 244.750 54.840 245.480 54.885 ;
        POLYGON 244.700 54.835 244.700 54.790 244.660 54.790 ;
        RECT 244.700 54.820 245.480 54.840 ;
        POLYGON 245.480 54.885 245.550 54.885 245.480 54.820 ;
        POLYGON 246.120 54.885 246.120 54.855 246.085 54.855 ;
        RECT 246.120 54.860 247.590 54.885 ;
        POLYGON 247.590 54.950 247.740 54.950 247.590 54.860 ;
        RECT 250.285 54.945 252.460 54.955 ;
        POLYGON 250.285 54.945 250.375 54.945 250.375 54.915 ;
        RECT 250.375 54.925 252.460 54.945 ;
        POLYGON 252.460 54.970 252.545 54.925 252.460 54.925 ;
        POLYGON 253.205 54.970 253.235 54.970 253.235 54.950 ;
        RECT 253.235 54.950 253.995 54.970 ;
        POLYGON 253.245 54.950 253.250 54.950 253.250 54.945 ;
        RECT 253.250 54.940 253.995 54.950 ;
        POLYGON 253.250 54.940 253.275 54.940 253.275 54.925 ;
        RECT 253.275 54.935 253.995 54.940 ;
        POLYGON 253.995 55.020 254.095 54.935 253.995 54.935 ;
        POLYGON 254.840 55.020 254.910 55.020 254.910 54.960 ;
        RECT 254.910 54.960 255.545 55.020 ;
        POLYGON 254.910 54.960 254.935 54.960 254.935 54.940 ;
        RECT 254.935 54.935 255.545 54.960 ;
        RECT 253.275 54.925 254.095 54.935 ;
        RECT 250.375 54.915 252.545 54.925 ;
        POLYGON 250.375 54.915 250.455 54.915 250.455 54.885 ;
        RECT 250.455 54.885 252.545 54.915 ;
        POLYGON 250.455 54.885 250.475 54.885 250.475 54.880 ;
        RECT 250.475 54.880 252.545 54.885 ;
        POLYGON 252.545 54.925 252.625 54.880 252.545 54.880 ;
        POLYGON 253.275 54.925 253.335 54.925 253.335 54.880 ;
        RECT 253.335 54.880 254.095 54.925 ;
        POLYGON 250.475 54.880 250.545 54.880 250.545 54.860 ;
        RECT 250.545 54.860 252.625 54.880 ;
        RECT 246.120 54.855 247.550 54.860 ;
        POLYGON 246.085 54.855 246.085 54.830 246.055 54.830 ;
        RECT 246.085 54.840 247.550 54.855 ;
        POLYGON 247.550 54.860 247.590 54.860 247.550 54.840 ;
        POLYGON 250.545 54.860 250.585 54.860 250.585 54.850 ;
        RECT 250.585 54.855 252.625 54.860 ;
        POLYGON 252.625 54.880 252.670 54.855 252.625 54.855 ;
        POLYGON 253.335 54.880 253.375 54.880 253.375 54.855 ;
        RECT 253.375 54.860 254.095 54.880 ;
        POLYGON 254.095 54.935 254.185 54.860 254.095 54.860 ;
        POLYGON 254.935 54.935 254.940 54.935 254.940 54.930 ;
        RECT 254.940 54.930 255.545 54.935 ;
        POLYGON 254.940 54.930 254.965 54.930 254.965 54.910 ;
        RECT 254.965 54.910 255.545 54.930 ;
        POLYGON 254.965 54.910 255.015 54.910 255.015 54.860 ;
        RECT 255.015 54.900 255.545 54.910 ;
        POLYGON 255.545 55.095 255.740 54.900 255.545 54.900 ;
        POLYGON 256.495 55.095 256.505 55.095 256.505 55.085 ;
        RECT 256.505 55.085 257.625 55.095 ;
        POLYGON 256.505 55.085 256.525 55.085 256.525 55.060 ;
        RECT 256.525 55.060 257.625 55.085 ;
        POLYGON 256.525 55.060 256.570 55.060 256.570 55.005 ;
        RECT 256.570 55.005 257.625 55.060 ;
        POLYGON 256.570 55.005 256.655 55.005 256.655 54.900 ;
        RECT 256.655 54.905 257.625 55.005 ;
        POLYGON 257.625 55.150 257.795 54.905 257.625 54.905 ;
        POLYGON 259.005 55.150 259.020 55.150 259.020 55.130 ;
        RECT 259.020 55.130 260.490 55.150 ;
        POLYGON 259.020 55.130 259.030 55.130 259.030 55.115 ;
        RECT 259.030 55.115 260.490 55.130 ;
        POLYGON 259.030 55.115 259.105 55.115 259.105 55.000 ;
        RECT 259.105 55.100 260.490 55.115 ;
        POLYGON 260.490 55.450 260.680 55.100 260.490 55.100 ;
        POLYGON 262.620 55.450 262.770 55.450 262.770 55.135 ;
        RECT 262.770 55.435 265.280 55.450 ;
        POLYGON 265.280 55.845 265.455 55.435 265.280 55.435 ;
        POLYGON 269.600 55.845 269.610 55.845 269.610 55.830 ;
        RECT 269.610 55.830 276.535 55.845 ;
        POLYGON 269.610 55.830 269.770 55.830 269.770 55.435 ;
        RECT 269.770 55.435 276.535 55.830 ;
        RECT 262.770 55.360 265.455 55.435 ;
        POLYGON 265.455 55.435 265.490 55.360 265.455 55.360 ;
        POLYGON 269.770 55.435 269.800 55.435 269.800 55.365 ;
        RECT 269.800 55.360 276.535 55.435 ;
        POLYGON 276.535 56.095 276.770 55.360 276.535 55.360 ;
        RECT 262.770 55.345 265.490 55.360 ;
        POLYGON 265.490 55.360 265.495 55.345 265.490 55.345 ;
        POLYGON 269.800 55.360 269.805 55.360 269.805 55.350 ;
        RECT 269.805 55.345 276.770 55.360 ;
        RECT 262.770 55.295 265.495 55.345 ;
        POLYGON 265.495 55.345 265.515 55.295 265.495 55.295 ;
        POLYGON 269.805 55.345 269.825 55.345 269.825 55.300 ;
        RECT 269.825 55.295 276.770 55.345 ;
        RECT 262.770 55.135 265.515 55.295 ;
        POLYGON 262.770 55.135 262.785 55.135 262.785 55.100 ;
        RECT 262.785 55.100 265.515 55.135 ;
        RECT 259.105 55.065 260.680 55.100 ;
        POLYGON 260.680 55.100 260.695 55.065 260.680 55.065 ;
        POLYGON 262.785 55.100 262.800 55.100 262.800 55.070 ;
        RECT 262.800 55.065 265.515 55.100 ;
        RECT 259.105 54.995 260.695 55.065 ;
        POLYGON 259.105 54.995 259.110 54.995 259.110 54.985 ;
        RECT 259.110 54.985 260.695 54.995 ;
        POLYGON 259.110 54.985 259.160 54.985 259.160 54.915 ;
        RECT 259.160 54.915 260.695 54.985 ;
        POLYGON 259.160 54.915 259.165 54.915 259.165 54.905 ;
        RECT 259.165 54.905 260.695 54.915 ;
        RECT 256.655 54.900 257.795 54.905 ;
        RECT 255.015 54.870 255.740 54.900 ;
        POLYGON 255.740 54.900 255.765 54.870 255.740 54.870 ;
        POLYGON 256.655 54.900 256.680 54.900 256.680 54.870 ;
        RECT 256.680 54.885 257.795 54.900 ;
        POLYGON 257.795 54.905 257.810 54.885 257.795 54.885 ;
        POLYGON 259.165 54.905 259.175 54.905 259.175 54.885 ;
        RECT 259.175 54.885 260.695 54.905 ;
        RECT 256.680 54.870 257.810 54.885 ;
        RECT 255.015 54.860 255.765 54.870 ;
        RECT 253.375 54.855 254.185 54.860 ;
        RECT 250.585 54.850 252.670 54.855 ;
        POLYGON 250.585 54.850 250.615 54.850 250.615 54.840 ;
        RECT 250.615 54.845 252.670 54.850 ;
        POLYGON 252.670 54.855 252.690 54.845 252.670 54.845 ;
        POLYGON 253.375 54.855 253.390 54.855 253.390 54.845 ;
        RECT 253.390 54.845 254.185 54.855 ;
        RECT 250.615 54.840 252.690 54.845 ;
        POLYGON 252.690 54.845 252.695 54.840 252.690 54.840 ;
        POLYGON 253.390 54.845 253.395 54.845 253.395 54.840 ;
        RECT 253.395 54.840 254.185 54.845 ;
        RECT 246.085 54.830 247.430 54.840 ;
        POLYGON 246.055 54.830 246.055 54.820 246.045 54.820 ;
        RECT 246.055 54.820 247.430 54.830 ;
        RECT 244.700 54.790 245.365 54.820 ;
        RECT 242.925 54.740 243.760 54.790 ;
        RECT 240.455 54.700 241.645 54.740 ;
        POLYGON 241.645 54.740 241.670 54.740 241.645 54.700 ;
        POLYGON 242.880 54.740 242.880 54.710 242.860 54.710 ;
        RECT 242.880 54.735 243.760 54.740 ;
        POLYGON 243.760 54.790 243.795 54.790 243.760 54.735 ;
        POLYGON 244.660 54.790 244.660 54.735 244.615 54.735 ;
        RECT 244.660 54.735 245.365 54.790 ;
        RECT 242.880 54.710 243.695 54.735 ;
        POLYGON 242.860 54.710 242.860 54.700 242.855 54.700 ;
        RECT 242.860 54.700 243.695 54.710 ;
        RECT 240.455 54.645 241.615 54.700 ;
        POLYGON 241.615 54.700 241.645 54.700 241.615 54.645 ;
        POLYGON 242.855 54.700 242.855 54.690 242.850 54.690 ;
        RECT 242.855 54.690 243.695 54.700 ;
        POLYGON 242.850 54.690 242.850 54.645 242.820 54.645 ;
        RECT 242.850 54.645 243.695 54.690 ;
        RECT 240.455 54.605 241.590 54.645 ;
        POLYGON 240.335 54.605 240.335 54.590 240.330 54.590 ;
        RECT 240.335 54.600 241.590 54.605 ;
        POLYGON 241.590 54.645 241.615 54.645 241.590 54.600 ;
        RECT 242.820 54.640 243.695 54.645 ;
        POLYGON 243.695 54.735 243.760 54.735 243.695 54.640 ;
        POLYGON 244.615 54.735 244.615 54.675 244.565 54.675 ;
        RECT 244.615 54.705 245.365 54.735 ;
        POLYGON 245.365 54.820 245.480 54.820 245.365 54.705 ;
        POLYGON 246.045 54.820 246.045 54.810 246.035 54.810 ;
        RECT 246.045 54.810 247.430 54.820 ;
        POLYGON 246.035 54.810 246.035 54.745 245.955 54.745 ;
        RECT 246.035 54.765 247.430 54.810 ;
        POLYGON 247.430 54.840 247.550 54.840 247.430 54.765 ;
        POLYGON 250.615 54.840 250.650 54.840 250.650 54.830 ;
        RECT 250.650 54.830 252.695 54.840 ;
        POLYGON 250.655 54.830 250.700 54.830 250.700 54.820 ;
        RECT 250.700 54.820 252.695 54.830 ;
        POLYGON 250.700 54.820 250.830 54.820 250.830 54.790 ;
        RECT 250.830 54.790 252.695 54.820 ;
        POLYGON 250.830 54.790 250.845 54.790 250.845 54.785 ;
        RECT 250.845 54.785 252.695 54.790 ;
        POLYGON 252.695 54.840 252.785 54.785 252.695 54.785 ;
        POLYGON 253.395 54.840 253.475 54.840 253.475 54.785 ;
        RECT 253.475 54.815 254.185 54.840 ;
        POLYGON 254.185 54.860 254.235 54.815 254.185 54.815 ;
        POLYGON 255.015 54.860 255.060 54.860 255.060 54.815 ;
        RECT 255.060 54.815 255.765 54.860 ;
        RECT 253.475 54.785 254.235 54.815 ;
        POLYGON 250.845 54.785 250.885 54.785 250.885 54.775 ;
        RECT 250.885 54.775 252.785 54.785 ;
        POLYGON 250.885 54.775 250.960 54.775 250.960 54.765 ;
        RECT 250.960 54.765 252.785 54.775 ;
        RECT 246.035 54.755 247.415 54.765 ;
        POLYGON 247.415 54.765 247.430 54.765 247.415 54.755 ;
        POLYGON 250.960 54.765 251.010 54.765 251.010 54.755 ;
        RECT 251.010 54.755 252.785 54.765 ;
        POLYGON 252.785 54.785 252.830 54.755 252.785 54.755 ;
        POLYGON 253.475 54.785 253.520 54.785 253.520 54.755 ;
        RECT 253.520 54.755 254.235 54.785 ;
        RECT 246.035 54.745 247.360 54.755 ;
        POLYGON 245.955 54.745 245.955 54.705 245.915 54.705 ;
        RECT 245.955 54.720 247.360 54.745 ;
        POLYGON 247.360 54.755 247.415 54.755 247.360 54.720 ;
        POLYGON 251.010 54.755 251.035 54.755 251.035 54.750 ;
        RECT 251.035 54.750 252.830 54.755 ;
        POLYGON 251.035 54.750 251.090 54.750 251.090 54.740 ;
        RECT 251.090 54.740 252.830 54.750 ;
        POLYGON 251.095 54.740 251.140 54.740 251.140 54.730 ;
        RECT 251.140 54.730 252.830 54.740 ;
        POLYGON 251.140 54.730 251.190 54.730 251.190 54.720 ;
        RECT 251.190 54.720 252.830 54.730 ;
        RECT 245.955 54.705 247.270 54.720 ;
        RECT 244.615 54.675 245.290 54.705 ;
        POLYGON 244.565 54.675 244.565 54.640 244.535 54.640 ;
        RECT 244.565 54.640 245.290 54.675 ;
        POLYGON 242.820 54.640 242.820 54.600 242.795 54.600 ;
        RECT 242.820 54.600 243.655 54.640 ;
        RECT 240.335 54.590 241.560 54.600 ;
        POLYGON 240.330 54.590 240.330 54.535 240.310 54.535 ;
        RECT 240.330 54.540 241.560 54.590 ;
        POLYGON 241.560 54.600 241.590 54.600 241.560 54.540 ;
        POLYGON 242.795 54.600 242.795 54.540 242.760 54.540 ;
        RECT 242.795 54.575 243.655 54.600 ;
        POLYGON 243.655 54.640 243.695 54.640 243.655 54.575 ;
        POLYGON 244.535 54.640 244.535 54.600 244.505 54.600 ;
        RECT 244.535 54.635 245.290 54.640 ;
        POLYGON 245.290 54.705 245.365 54.705 245.290 54.635 ;
        POLYGON 245.915 54.705 245.915 54.635 245.845 54.635 ;
        RECT 245.915 54.660 247.270 54.705 ;
        POLYGON 247.270 54.720 247.360 54.720 247.270 54.660 ;
        POLYGON 251.190 54.720 251.220 54.720 251.220 54.715 ;
        RECT 251.220 54.715 252.830 54.720 ;
        POLYGON 251.235 54.715 251.295 54.715 251.295 54.700 ;
        RECT 251.295 54.700 252.830 54.715 ;
        POLYGON 251.295 54.700 251.370 54.700 251.370 54.685 ;
        RECT 251.370 54.685 252.830 54.700 ;
        POLYGON 252.830 54.755 252.940 54.685 252.830 54.685 ;
        POLYGON 253.520 54.755 253.535 54.755 253.535 54.745 ;
        RECT 253.535 54.745 254.235 54.755 ;
        POLYGON 253.535 54.745 253.555 54.745 253.555 54.730 ;
        RECT 253.555 54.740 254.235 54.745 ;
        POLYGON 254.235 54.815 254.310 54.740 254.235 54.740 ;
        POLYGON 255.060 54.815 255.080 54.815 255.080 54.795 ;
        RECT 255.080 54.795 255.765 54.815 ;
        POLYGON 255.080 54.795 255.135 54.795 255.135 54.745 ;
        RECT 255.135 54.740 255.765 54.795 ;
        POLYGON 255.765 54.870 255.880 54.740 255.765 54.740 ;
        POLYGON 256.680 54.870 256.710 54.870 256.710 54.835 ;
        RECT 256.710 54.855 257.810 54.870 ;
        POLYGON 257.810 54.885 257.830 54.855 257.810 54.855 ;
        POLYGON 259.175 54.885 259.185 54.885 259.185 54.870 ;
        RECT 259.185 54.870 260.695 54.885 ;
        POLYGON 259.185 54.870 259.190 54.870 259.190 54.860 ;
        RECT 259.190 54.855 260.695 54.870 ;
        RECT 256.710 54.835 257.830 54.855 ;
        POLYGON 256.710 54.835 256.715 54.835 256.715 54.830 ;
        RECT 256.715 54.830 257.830 54.835 ;
        POLYGON 256.715 54.830 256.755 54.830 256.755 54.780 ;
        RECT 256.755 54.780 257.830 54.830 ;
        POLYGON 256.755 54.780 256.765 54.780 256.765 54.765 ;
        RECT 256.765 54.765 257.830 54.780 ;
        POLYGON 256.765 54.765 256.780 54.765 256.780 54.745 ;
        RECT 256.780 54.740 257.830 54.765 ;
        RECT 253.555 54.730 254.310 54.740 ;
        POLYGON 253.555 54.730 253.610 54.730 253.610 54.685 ;
        RECT 253.610 54.705 254.310 54.730 ;
        POLYGON 254.310 54.740 254.350 54.705 254.310 54.705 ;
        POLYGON 255.135 54.740 255.170 54.740 255.170 54.705 ;
        RECT 255.170 54.730 255.880 54.740 ;
        POLYGON 255.880 54.740 255.890 54.730 255.880 54.730 ;
        POLYGON 256.780 54.740 256.790 54.740 256.790 54.730 ;
        RECT 256.790 54.730 257.830 54.740 ;
        RECT 255.170 54.705 255.890 54.730 ;
        RECT 253.610 54.685 254.350 54.705 ;
        POLYGON 251.375 54.685 251.410 54.685 251.410 54.675 ;
        RECT 251.410 54.675 252.940 54.685 ;
        POLYGON 252.940 54.685 252.955 54.675 252.940 54.675 ;
        POLYGON 253.610 54.685 253.625 54.685 253.625 54.675 ;
        RECT 253.625 54.675 254.350 54.685 ;
        POLYGON 251.410 54.675 251.450 54.675 251.450 54.665 ;
        RECT 251.450 54.665 252.955 54.675 ;
        POLYGON 252.955 54.675 252.975 54.665 252.955 54.665 ;
        POLYGON 253.625 54.675 253.640 54.675 253.640 54.665 ;
        RECT 253.640 54.665 254.350 54.675 ;
        POLYGON 251.450 54.665 251.465 54.665 251.465 54.660 ;
        RECT 251.465 54.660 252.975 54.665 ;
        RECT 245.915 54.635 247.175 54.660 ;
        RECT 244.535 54.600 245.250 54.635 ;
        POLYGON 244.505 54.600 244.505 54.575 244.485 54.575 ;
        RECT 244.505 54.590 245.250 54.600 ;
        POLYGON 245.250 54.635 245.290 54.635 245.250 54.590 ;
        POLYGON 245.845 54.635 245.845 54.615 245.820 54.615 ;
        RECT 245.845 54.615 247.175 54.635 ;
        POLYGON 245.820 54.615 245.820 54.590 245.795 54.590 ;
        RECT 245.820 54.595 247.175 54.615 ;
        POLYGON 247.175 54.660 247.270 54.660 247.175 54.595 ;
        POLYGON 251.465 54.660 251.515 54.660 251.515 54.645 ;
        RECT 251.515 54.655 252.975 54.660 ;
        POLYGON 252.975 54.665 252.985 54.655 252.975 54.655 ;
        POLYGON 253.640 54.665 253.650 54.665 253.650 54.655 ;
        RECT 253.650 54.655 254.350 54.665 ;
        RECT 251.515 54.645 252.985 54.655 ;
        POLYGON 251.515 54.645 251.590 54.645 251.590 54.625 ;
        RECT 251.590 54.625 252.985 54.645 ;
        POLYGON 251.595 54.625 251.605 54.625 251.605 54.620 ;
        RECT 251.605 54.620 252.985 54.625 ;
        POLYGON 251.605 54.620 251.660 54.620 251.660 54.600 ;
        RECT 251.660 54.600 252.985 54.620 ;
        POLYGON 251.660 54.600 251.670 54.600 251.670 54.595 ;
        RECT 251.670 54.595 252.985 54.600 ;
        RECT 245.820 54.590 247.150 54.595 ;
        RECT 244.505 54.575 245.225 54.590 ;
        RECT 242.795 54.565 243.650 54.575 ;
        POLYGON 243.650 54.575 243.655 54.575 243.650 54.565 ;
        POLYGON 244.485 54.575 244.485 54.565 244.475 54.565 ;
        RECT 244.485 54.565 245.225 54.575 ;
        POLYGON 245.225 54.590 245.250 54.590 245.225 54.565 ;
        POLYGON 245.795 54.590 245.795 54.565 245.765 54.565 ;
        RECT 245.795 54.575 247.150 54.590 ;
        POLYGON 247.150 54.595 247.175 54.595 247.150 54.575 ;
        POLYGON 251.670 54.595 251.730 54.595 251.730 54.575 ;
        RECT 251.730 54.580 252.985 54.595 ;
        POLYGON 252.985 54.655 253.095 54.580 252.985 54.580 ;
        POLYGON 253.650 54.655 253.660 54.655 253.660 54.650 ;
        RECT 253.660 54.650 254.350 54.655 ;
        POLYGON 253.660 54.650 253.670 54.650 253.670 54.640 ;
        RECT 253.670 54.640 254.350 54.650 ;
        POLYGON 253.670 54.640 253.745 54.640 253.745 54.580 ;
        RECT 253.745 54.620 254.350 54.640 ;
        POLYGON 254.350 54.705 254.445 54.620 254.350 54.620 ;
        POLYGON 255.170 54.705 255.175 54.705 255.175 54.700 ;
        RECT 255.175 54.700 255.890 54.705 ;
        POLYGON 255.175 54.700 255.245 54.700 255.245 54.625 ;
        RECT 255.245 54.620 255.890 54.700 ;
        RECT 253.745 54.590 254.445 54.620 ;
        POLYGON 254.445 54.620 254.475 54.590 254.445 54.590 ;
        POLYGON 255.245 54.620 255.275 54.620 255.275 54.590 ;
        RECT 255.275 54.590 255.890 54.620 ;
        POLYGON 255.890 54.730 256.015 54.590 255.890 54.590 ;
        POLYGON 256.790 54.730 256.855 54.730 256.855 54.650 ;
        RECT 256.855 54.695 257.830 54.730 ;
        POLYGON 257.830 54.855 257.935 54.695 257.830 54.695 ;
        POLYGON 259.190 54.855 259.240 54.855 259.240 54.780 ;
        RECT 259.240 54.780 260.695 54.855 ;
        POLYGON 260.695 55.065 260.835 54.780 260.695 54.780 ;
        POLYGON 262.800 55.065 262.815 55.065 262.815 55.040 ;
        RECT 262.815 55.040 265.515 55.065 ;
        POLYGON 262.815 55.040 262.925 55.040 262.925 54.785 ;
        RECT 262.925 54.800 265.515 55.040 ;
        POLYGON 265.515 55.295 265.705 54.800 265.515 54.800 ;
        POLYGON 269.825 55.295 269.845 55.295 269.845 55.255 ;
        RECT 269.845 55.255 276.770 55.295 ;
        POLYGON 269.845 55.255 269.885 55.255 269.885 55.150 ;
        RECT 269.885 55.150 276.770 55.255 ;
        POLYGON 269.885 55.150 270.010 55.150 270.010 54.805 ;
        RECT 270.010 54.895 276.770 55.150 ;
        POLYGON 276.770 55.360 276.895 54.895 276.770 54.895 ;
        RECT 270.010 54.800 276.895 54.895 ;
        RECT 262.925 54.780 265.705 54.800 ;
        POLYGON 259.240 54.780 259.245 54.780 259.245 54.765 ;
        RECT 259.245 54.765 260.835 54.780 ;
        POLYGON 259.245 54.765 259.285 54.765 259.285 54.695 ;
        RECT 259.285 54.740 260.835 54.765 ;
        POLYGON 260.835 54.780 260.850 54.740 260.835 54.740 ;
        POLYGON 262.925 54.780 262.940 54.780 262.940 54.750 ;
        RECT 262.940 54.740 265.705 54.780 ;
        RECT 259.285 54.695 260.850 54.740 ;
        RECT 256.855 54.650 257.935 54.695 ;
        POLYGON 256.855 54.650 256.895 54.650 256.895 54.595 ;
        RECT 256.895 54.640 257.935 54.650 ;
        POLYGON 257.935 54.695 257.975 54.640 257.935 54.640 ;
        POLYGON 259.285 54.695 259.300 54.695 259.300 54.680 ;
        RECT 259.300 54.680 260.850 54.695 ;
        POLYGON 259.300 54.680 259.320 54.680 259.320 54.640 ;
        RECT 259.320 54.640 260.850 54.680 ;
        RECT 256.895 54.615 257.975 54.640 ;
        POLYGON 257.975 54.640 257.990 54.615 257.975 54.615 ;
        POLYGON 259.320 54.640 259.335 54.640 259.335 54.615 ;
        RECT 259.335 54.615 260.850 54.640 ;
        RECT 256.895 54.590 257.990 54.615 ;
        RECT 253.745 54.580 254.475 54.590 ;
        RECT 251.730 54.575 253.095 54.580 ;
        RECT 245.795 54.565 247.115 54.575 ;
        RECT 242.795 54.555 243.640 54.565 ;
        POLYGON 243.640 54.565 243.650 54.565 243.640 54.555 ;
        POLYGON 244.475 54.565 244.475 54.560 244.470 54.560 ;
        RECT 244.475 54.560 245.190 54.565 ;
        RECT 242.795 54.540 243.555 54.555 ;
        RECT 240.330 54.535 241.550 54.540 ;
        RECT 236.545 54.525 238.635 54.530 ;
        POLYGON 238.635 54.530 238.640 54.530 238.635 54.525 ;
        POLYGON 240.310 54.530 240.310 54.525 240.305 54.525 ;
        RECT 240.310 54.525 241.550 54.535 ;
        POLYGON 241.550 54.540 241.560 54.540 241.550 54.525 ;
        POLYGON 242.760 54.540 242.760 54.525 242.750 54.525 ;
        RECT 242.760 54.525 243.555 54.540 ;
        RECT 236.545 54.505 238.605 54.525 ;
        POLYGON 236.485 54.505 236.485 54.120 236.390 54.120 ;
        RECT 236.485 54.430 238.605 54.505 ;
        POLYGON 238.605 54.525 238.635 54.525 238.605 54.430 ;
        POLYGON 240.305 54.525 240.305 54.430 240.270 54.430 ;
        RECT 240.305 54.470 241.525 54.525 ;
        POLYGON 241.525 54.525 241.550 54.525 241.525 54.470 ;
        POLYGON 242.750 54.525 242.750 54.475 242.720 54.475 ;
        RECT 242.750 54.475 243.555 54.525 ;
        RECT 240.305 54.445 241.510 54.470 ;
        POLYGON 241.510 54.470 241.525 54.470 241.510 54.445 ;
        POLYGON 242.720 54.470 242.720 54.450 242.705 54.450 ;
        RECT 242.720 54.450 243.555 54.475 ;
        RECT 240.305 54.430 241.465 54.445 ;
        RECT 236.485 54.395 238.595 54.430 ;
        POLYGON 238.595 54.430 238.605 54.430 238.595 54.395 ;
        POLYGON 240.270 54.430 240.270 54.400 240.260 54.400 ;
        RECT 240.270 54.400 241.465 54.430 ;
        RECT 236.485 54.120 238.495 54.395 ;
        POLYGON 236.390 54.120 236.390 54.105 236.385 54.105 ;
        RECT 236.390 54.105 238.495 54.120 ;
        RECT 229.485 54.090 233.430 54.105 ;
        POLYGON 229.305 54.090 229.305 53.075 229.230 53.075 ;
        RECT 229.305 53.870 233.430 54.090 ;
        POLYGON 233.430 54.105 233.475 54.105 233.430 53.870 ;
        POLYGON 236.385 54.100 236.385 53.875 236.330 53.875 ;
        RECT 236.385 54.085 238.495 54.105 ;
        POLYGON 238.495 54.395 238.595 54.395 238.495 54.085 ;
        POLYGON 240.260 54.395 240.260 54.320 240.230 54.320 ;
        RECT 240.260 54.355 241.465 54.400 ;
        POLYGON 241.465 54.445 241.510 54.445 241.465 54.355 ;
        POLYGON 242.705 54.445 242.705 54.415 242.685 54.415 ;
        RECT 242.705 54.415 243.555 54.450 ;
        POLYGON 243.555 54.555 243.640 54.555 243.555 54.415 ;
        POLYGON 244.470 54.555 244.470 54.485 244.410 54.485 ;
        RECT 244.470 54.525 245.190 54.560 ;
        POLYGON 245.190 54.565 245.225 54.565 245.190 54.525 ;
        POLYGON 245.765 54.565 245.765 54.525 245.725 54.525 ;
        RECT 245.765 54.550 247.115 54.565 ;
        POLYGON 247.115 54.575 247.150 54.575 247.115 54.550 ;
        POLYGON 251.730 54.575 251.760 54.575 251.760 54.565 ;
        RECT 251.760 54.570 253.095 54.575 ;
        POLYGON 253.095 54.580 253.115 54.570 253.095 54.570 ;
        POLYGON 253.745 54.580 253.760 54.580 253.760 54.570 ;
        RECT 253.760 54.570 254.475 54.580 ;
        RECT 251.760 54.565 253.115 54.570 ;
        POLYGON 251.760 54.565 251.770 54.565 251.770 54.560 ;
        RECT 251.770 54.560 253.115 54.565 ;
        POLYGON 251.775 54.560 251.805 54.560 251.805 54.550 ;
        RECT 251.805 54.550 253.115 54.560 ;
        RECT 245.765 54.525 247.085 54.550 ;
        POLYGON 247.085 54.550 247.115 54.550 247.085 54.525 ;
        POLYGON 251.805 54.550 251.865 54.550 251.865 54.525 ;
        RECT 251.865 54.525 253.115 54.550 ;
        RECT 244.470 54.485 245.110 54.525 ;
        POLYGON 244.410 54.485 244.410 54.415 244.360 54.415 ;
        RECT 244.410 54.445 245.110 54.485 ;
        POLYGON 245.110 54.525 245.190 54.525 245.110 54.445 ;
        POLYGON 245.725 54.525 245.725 54.470 245.675 54.470 ;
        RECT 245.725 54.470 246.995 54.525 ;
        POLYGON 245.675 54.470 245.675 54.445 245.655 54.445 ;
        RECT 245.675 54.460 246.995 54.470 ;
        POLYGON 246.995 54.525 247.085 54.525 246.995 54.460 ;
        POLYGON 251.865 54.525 251.915 54.525 251.915 54.505 ;
        RECT 251.915 54.505 253.115 54.525 ;
        POLYGON 251.915 54.505 252.020 54.505 252.020 54.460 ;
        RECT 252.020 54.480 253.115 54.505 ;
        POLYGON 253.115 54.570 253.235 54.480 253.115 54.480 ;
        POLYGON 253.760 54.570 253.795 54.570 253.795 54.545 ;
        RECT 253.795 54.545 254.475 54.570 ;
        POLYGON 253.795 54.545 253.805 54.545 253.805 54.535 ;
        RECT 253.805 54.535 254.475 54.545 ;
        POLYGON 254.475 54.590 254.525 54.535 254.475 54.535 ;
        POLYGON 255.275 54.590 255.320 54.590 255.320 54.545 ;
        RECT 255.320 54.565 256.015 54.590 ;
        POLYGON 256.015 54.590 256.035 54.565 256.015 54.565 ;
        POLYGON 256.895 54.590 256.915 54.590 256.915 54.565 ;
        RECT 256.915 54.565 257.990 54.590 ;
        RECT 255.320 54.545 256.035 54.565 ;
        POLYGON 255.320 54.545 255.325 54.545 255.325 54.535 ;
        RECT 255.325 54.535 256.035 54.545 ;
        POLYGON 253.805 54.535 253.820 54.535 253.820 54.525 ;
        RECT 253.820 54.525 254.525 54.535 ;
        POLYGON 253.820 54.525 253.875 54.525 253.875 54.480 ;
        RECT 253.875 54.480 254.525 54.525 ;
        RECT 252.020 54.475 253.235 54.480 ;
        POLYGON 253.235 54.480 253.245 54.475 253.235 54.475 ;
        POLYGON 253.875 54.480 253.880 54.480 253.880 54.475 ;
        RECT 253.880 54.475 254.525 54.480 ;
        RECT 252.020 54.470 253.245 54.475 ;
        POLYGON 253.245 54.475 253.250 54.470 253.245 54.470 ;
        POLYGON 253.880 54.475 253.885 54.475 253.885 54.470 ;
        RECT 253.885 54.470 254.525 54.475 ;
        RECT 252.020 54.460 253.250 54.470 ;
        RECT 245.675 54.445 246.965 54.460 ;
        RECT 244.410 54.415 245.065 54.445 ;
        POLYGON 242.685 54.415 242.685 54.360 242.655 54.360 ;
        RECT 242.685 54.360 243.490 54.415 ;
        RECT 240.260 54.320 241.425 54.355 ;
        POLYGON 240.230 54.320 240.230 54.260 240.210 54.260 ;
        RECT 240.230 54.275 241.425 54.320 ;
        POLYGON 241.425 54.355 241.465 54.355 241.425 54.285 ;
        POLYGON 242.655 54.355 242.655 54.285 242.615 54.285 ;
        RECT 242.655 54.315 243.490 54.360 ;
        POLYGON 243.490 54.415 243.555 54.415 243.490 54.315 ;
        POLYGON 244.360 54.415 244.360 54.385 244.340 54.385 ;
        RECT 244.360 54.395 245.065 54.415 ;
        POLYGON 245.065 54.445 245.110 54.445 245.065 54.395 ;
        POLYGON 245.655 54.445 245.655 54.395 245.605 54.395 ;
        RECT 245.655 54.440 246.965 54.445 ;
        POLYGON 246.965 54.460 246.995 54.460 246.965 54.440 ;
        POLYGON 252.020 54.460 252.070 54.460 252.070 54.440 ;
        RECT 252.070 54.455 253.250 54.460 ;
        POLYGON 253.250 54.470 253.275 54.455 253.250 54.455 ;
        POLYGON 253.885 54.470 253.905 54.470 253.905 54.455 ;
        RECT 253.905 54.455 254.525 54.470 ;
        RECT 252.070 54.440 253.275 54.455 ;
        RECT 245.655 54.395 246.890 54.440 ;
        RECT 244.360 54.385 245.040 54.395 ;
        POLYGON 244.340 54.385 244.340 54.355 244.315 54.355 ;
        RECT 244.340 54.365 245.040 54.385 ;
        POLYGON 245.040 54.395 245.065 54.395 245.040 54.365 ;
        POLYGON 245.605 54.395 245.605 54.365 245.575 54.365 ;
        RECT 245.605 54.380 246.890 54.395 ;
        POLYGON 246.890 54.440 246.965 54.440 246.890 54.380 ;
        POLYGON 252.070 54.440 252.100 54.440 252.100 54.425 ;
        RECT 252.100 54.425 253.275 54.440 ;
        POLYGON 252.100 54.425 252.120 54.425 252.120 54.410 ;
        RECT 252.120 54.410 253.275 54.425 ;
        POLYGON 252.125 54.410 252.185 54.410 252.185 54.380 ;
        RECT 252.185 54.380 253.275 54.410 ;
        RECT 245.605 54.365 246.830 54.380 ;
        RECT 244.340 54.355 245.025 54.365 ;
        POLYGON 244.315 54.355 244.315 54.315 244.285 54.315 ;
        RECT 244.315 54.345 245.025 54.355 ;
        POLYGON 245.025 54.365 245.040 54.365 245.025 54.345 ;
        POLYGON 245.575 54.365 245.575 54.345 245.555 54.345 ;
        RECT 245.575 54.345 246.830 54.365 ;
        RECT 244.315 54.315 244.935 54.345 ;
        RECT 242.655 54.285 243.460 54.315 ;
        RECT 240.230 54.260 241.330 54.275 ;
        POLYGON 240.210 54.260 240.210 54.085 240.150 54.085 ;
        RECT 240.210 54.085 241.330 54.260 ;
        RECT 236.385 53.875 238.435 54.085 ;
        POLYGON 238.435 54.085 238.495 54.085 238.435 53.875 ;
        POLYGON 240.150 54.085 240.150 53.925 240.095 53.925 ;
        RECT 240.150 54.065 241.330 54.085 ;
        POLYGON 241.330 54.275 241.425 54.275 241.330 54.065 ;
        POLYGON 242.615 54.285 242.615 54.230 242.585 54.230 ;
        RECT 242.615 54.260 243.460 54.285 ;
        POLYGON 243.460 54.315 243.490 54.315 243.460 54.260 ;
        POLYGON 244.285 54.315 244.285 54.285 244.265 54.285 ;
        RECT 244.285 54.285 244.935 54.315 ;
        POLYGON 244.265 54.285 244.265 54.265 244.250 54.265 ;
        RECT 244.265 54.265 244.935 54.285 ;
        RECT 242.615 54.230 243.435 54.260 ;
        POLYGON 242.585 54.230 242.585 54.200 242.565 54.200 ;
        RECT 242.585 54.215 243.435 54.230 ;
        POLYGON 243.435 54.260 243.460 54.260 243.435 54.215 ;
        POLYGON 244.250 54.260 244.250 54.215 244.215 54.215 ;
        RECT 244.250 54.245 244.935 54.265 ;
        POLYGON 244.935 54.345 245.025 54.345 244.935 54.245 ;
        POLYGON 245.555 54.345 245.555 54.340 245.550 54.340 ;
        RECT 245.555 54.340 246.830 54.345 ;
        POLYGON 245.550 54.340 245.550 54.260 245.480 54.260 ;
        RECT 245.550 54.330 246.830 54.340 ;
        POLYGON 246.830 54.380 246.890 54.380 246.830 54.330 ;
        POLYGON 252.185 54.380 252.220 54.380 252.220 54.365 ;
        RECT 252.220 54.365 253.275 54.380 ;
        POLYGON 253.275 54.455 253.390 54.365 253.275 54.365 ;
        POLYGON 253.905 54.455 253.925 54.455 253.925 54.440 ;
        RECT 253.925 54.440 254.525 54.455 ;
        POLYGON 253.925 54.440 253.935 54.440 253.935 54.430 ;
        RECT 253.935 54.430 254.525 54.440 ;
        POLYGON 253.935 54.430 254.010 54.430 254.010 54.365 ;
        RECT 254.010 54.365 254.525 54.430 ;
        POLYGON 252.220 54.365 252.285 54.365 252.285 54.330 ;
        RECT 252.285 54.330 253.390 54.365 ;
        RECT 245.550 54.320 246.820 54.330 ;
        POLYGON 246.820 54.330 246.830 54.330 246.820 54.320 ;
        POLYGON 252.285 54.330 252.305 54.330 252.305 54.320 ;
        RECT 252.305 54.320 253.390 54.330 ;
        RECT 245.550 54.260 246.675 54.320 ;
        POLYGON 245.480 54.260 245.480 54.250 245.470 54.250 ;
        RECT 245.480 54.250 246.675 54.260 ;
        RECT 244.250 54.215 244.890 54.245 ;
        RECT 242.585 54.200 243.395 54.215 ;
        POLYGON 242.565 54.200 242.565 54.125 242.525 54.125 ;
        RECT 242.565 54.145 243.395 54.200 ;
        POLYGON 243.395 54.215 243.435 54.215 243.395 54.145 ;
        POLYGON 244.215 54.210 244.215 54.145 244.170 54.145 ;
        RECT 244.215 54.190 244.890 54.215 ;
        POLYGON 244.890 54.245 244.935 54.245 244.890 54.190 ;
        POLYGON 245.470 54.245 245.470 54.210 245.440 54.210 ;
        RECT 245.470 54.210 246.675 54.250 ;
        POLYGON 245.440 54.210 245.440 54.190 245.425 54.190 ;
        RECT 245.440 54.195 246.675 54.210 ;
        POLYGON 246.675 54.320 246.820 54.320 246.675 54.195 ;
        POLYGON 252.305 54.320 252.375 54.320 252.375 54.285 ;
        RECT 252.375 54.285 253.390 54.320 ;
        POLYGON 252.375 54.285 252.395 54.285 252.395 54.270 ;
        RECT 252.395 54.270 253.390 54.285 ;
        POLYGON 253.390 54.365 253.520 54.270 253.390 54.270 ;
        POLYGON 254.010 54.365 254.065 54.365 254.065 54.320 ;
        RECT 254.065 54.350 254.525 54.365 ;
        POLYGON 254.525 54.535 254.710 54.350 254.525 54.350 ;
        POLYGON 255.325 54.535 255.345 54.535 255.345 54.515 ;
        RECT 255.345 54.520 256.035 54.535 ;
        POLYGON 256.035 54.565 256.070 54.520 256.035 54.520 ;
        POLYGON 256.915 54.565 256.950 54.565 256.950 54.520 ;
        RECT 256.950 54.520 257.990 54.565 ;
        RECT 255.345 54.515 256.070 54.520 ;
        POLYGON 255.345 54.515 255.400 54.515 255.400 54.455 ;
        RECT 255.400 54.455 256.070 54.515 ;
        POLYGON 255.400 54.455 255.480 54.455 255.480 54.360 ;
        RECT 255.480 54.360 256.070 54.455 ;
        POLYGON 256.070 54.520 256.195 54.360 256.070 54.360 ;
        POLYGON 256.950 54.520 256.995 54.520 256.995 54.460 ;
        RECT 256.995 54.460 257.990 54.520 ;
        POLYGON 256.995 54.460 257.005 54.460 257.005 54.445 ;
        RECT 257.005 54.445 257.990 54.460 ;
        POLYGON 257.005 54.445 257.060 54.445 257.060 54.365 ;
        RECT 257.060 54.400 257.990 54.445 ;
        POLYGON 257.990 54.615 258.120 54.400 257.990 54.400 ;
        POLYGON 259.335 54.615 259.340 54.615 259.340 54.610 ;
        RECT 259.340 54.610 260.850 54.615 ;
        POLYGON 259.340 54.610 259.365 54.610 259.365 54.560 ;
        RECT 259.365 54.560 260.850 54.610 ;
        RECT 259.370 54.555 260.850 54.560 ;
        POLYGON 259.370 54.555 259.385 54.555 259.385 54.530 ;
        RECT 259.385 54.530 260.850 54.555 ;
        POLYGON 260.850 54.740 260.945 54.530 260.850 54.530 ;
        POLYGON 262.940 54.740 263.020 54.740 263.020 54.565 ;
        RECT 263.020 54.735 265.705 54.740 ;
        POLYGON 265.705 54.800 265.730 54.735 265.705 54.735 ;
        POLYGON 270.010 54.800 270.035 54.800 270.035 54.740 ;
        RECT 270.035 54.735 276.895 54.800 ;
        RECT 263.020 54.565 265.730 54.735 ;
        POLYGON 263.020 54.565 263.030 54.565 263.030 54.535 ;
        RECT 263.030 54.530 265.730 54.565 ;
        POLYGON 259.385 54.530 259.390 54.530 259.390 54.525 ;
        RECT 259.390 54.520 260.945 54.530 ;
        POLYGON 259.390 54.520 259.400 54.520 259.400 54.505 ;
        RECT 259.400 54.505 260.945 54.520 ;
        POLYGON 259.400 54.505 259.455 54.505 259.455 54.400 ;
        RECT 259.455 54.400 260.945 54.505 ;
        RECT 257.060 54.370 258.120 54.400 ;
        POLYGON 258.120 54.400 258.140 54.370 258.120 54.370 ;
        POLYGON 259.455 54.400 259.470 54.400 259.470 54.370 ;
        RECT 259.470 54.375 260.945 54.400 ;
        POLYGON 260.945 54.530 261.015 54.375 260.945 54.375 ;
        POLYGON 263.030 54.530 263.090 54.530 263.090 54.375 ;
        RECT 263.090 54.375 265.730 54.530 ;
        RECT 259.470 54.370 261.015 54.375 ;
        RECT 257.060 54.360 258.140 54.370 ;
        POLYGON 255.480 54.360 255.490 54.360 255.490 54.350 ;
        RECT 255.490 54.350 256.195 54.360 ;
        RECT 254.065 54.325 254.710 54.350 ;
        POLYGON 254.710 54.350 254.730 54.325 254.710 54.325 ;
        POLYGON 255.490 54.350 255.495 54.350 255.495 54.345 ;
        RECT 255.495 54.345 256.195 54.350 ;
        POLYGON 255.495 54.345 255.510 54.345 255.510 54.325 ;
        RECT 255.510 54.325 256.195 54.345 ;
        RECT 254.065 54.320 254.730 54.325 ;
        POLYGON 254.065 54.320 254.075 54.320 254.075 54.310 ;
        RECT 254.075 54.310 254.730 54.320 ;
        POLYGON 254.075 54.310 254.120 54.310 254.120 54.270 ;
        RECT 254.120 54.270 254.730 54.310 ;
        POLYGON 252.395 54.270 252.460 54.270 252.460 54.235 ;
        RECT 252.460 54.255 253.520 54.270 ;
        POLYGON 253.520 54.270 253.535 54.255 253.520 54.255 ;
        POLYGON 254.120 54.270 254.135 54.270 254.135 54.255 ;
        RECT 254.135 54.255 254.730 54.270 ;
        RECT 252.460 54.240 253.535 54.255 ;
        POLYGON 253.535 54.255 253.555 54.240 253.535 54.240 ;
        POLYGON 254.135 54.255 254.155 54.255 254.155 54.240 ;
        RECT 254.155 54.240 254.730 54.255 ;
        RECT 252.460 54.235 253.555 54.240 ;
        POLYGON 252.460 54.235 252.525 54.235 252.525 54.195 ;
        RECT 252.525 54.195 253.555 54.235 ;
        RECT 245.440 54.190 246.650 54.195 ;
        RECT 244.215 54.165 244.875 54.190 ;
        POLYGON 244.875 54.190 244.890 54.190 244.875 54.165 ;
        POLYGON 245.425 54.190 245.425 54.165 245.400 54.165 ;
        RECT 245.425 54.175 246.650 54.190 ;
        POLYGON 246.650 54.195 246.675 54.195 246.650 54.175 ;
        POLYGON 252.525 54.195 252.555 54.195 252.555 54.175 ;
        RECT 252.555 54.175 253.555 54.195 ;
        RECT 245.425 54.170 246.645 54.175 ;
        POLYGON 246.645 54.175 246.650 54.175 246.645 54.170 ;
        POLYGON 252.555 54.175 252.565 54.175 252.565 54.170 ;
        RECT 252.565 54.170 253.555 54.175 ;
        RECT 245.425 54.165 246.535 54.170 ;
        RECT 244.215 54.155 244.865 54.165 ;
        POLYGON 244.865 54.165 244.875 54.165 244.865 54.155 ;
        POLYGON 245.400 54.165 245.400 54.155 245.390 54.155 ;
        RECT 245.400 54.155 246.535 54.165 ;
        RECT 244.215 54.145 244.770 54.155 ;
        RECT 242.565 54.125 243.375 54.145 ;
        POLYGON 242.525 54.120 242.525 54.065 242.495 54.065 ;
        RECT 242.525 54.115 243.375 54.125 ;
        POLYGON 243.375 54.145 243.395 54.145 243.375 54.115 ;
        POLYGON 244.170 54.145 244.170 54.115 244.150 54.115 ;
        RECT 244.170 54.115 244.770 54.145 ;
        RECT 242.525 54.070 243.350 54.115 ;
        POLYGON 243.350 54.115 243.375 54.115 243.350 54.070 ;
        POLYGON 244.150 54.115 244.150 54.095 244.135 54.095 ;
        RECT 244.150 54.095 244.770 54.115 ;
        POLYGON 244.135 54.095 244.135 54.085 244.130 54.085 ;
        RECT 244.135 54.085 244.770 54.095 ;
        POLYGON 244.130 54.085 244.130 54.070 244.120 54.070 ;
        RECT 244.130 54.070 244.770 54.085 ;
        RECT 242.525 54.065 243.300 54.070 ;
        RECT 240.150 54.055 241.325 54.065 ;
        POLYGON 241.325 54.065 241.330 54.065 241.325 54.055 ;
        POLYGON 242.495 54.060 242.495 54.055 242.490 54.055 ;
        RECT 242.495 54.055 243.300 54.065 ;
        RECT 240.150 53.935 241.270 54.055 ;
        POLYGON 241.270 54.055 241.325 54.055 241.270 53.935 ;
        POLYGON 242.490 54.050 242.490 53.935 242.430 53.935 ;
        RECT 242.490 53.970 243.300 54.055 ;
        POLYGON 243.300 54.070 243.350 54.070 243.300 53.970 ;
        POLYGON 244.120 54.070 244.120 54.045 244.100 54.045 ;
        RECT 244.120 54.045 244.770 54.070 ;
        POLYGON 244.100 54.045 244.100 53.975 244.055 53.975 ;
        RECT 244.100 54.040 244.770 54.045 ;
        POLYGON 244.770 54.155 244.865 54.155 244.770 54.040 ;
        POLYGON 245.390 54.155 245.390 54.125 245.365 54.125 ;
        RECT 245.390 54.125 246.535 54.155 ;
        POLYGON 245.365 54.125 245.365 54.045 245.300 54.045 ;
        RECT 245.365 54.070 246.535 54.125 ;
        POLYGON 246.535 54.170 246.645 54.170 246.535 54.070 ;
        POLYGON 252.565 54.170 252.625 54.170 252.625 54.135 ;
        RECT 252.625 54.150 253.555 54.170 ;
        POLYGON 253.555 54.240 253.660 54.150 253.555 54.150 ;
        POLYGON 254.155 54.240 254.185 54.240 254.185 54.215 ;
        RECT 254.185 54.215 254.730 54.240 ;
        POLYGON 254.185 54.215 254.255 54.215 254.255 54.150 ;
        RECT 254.255 54.150 254.730 54.215 ;
        RECT 252.625 54.140 253.660 54.150 ;
        POLYGON 253.660 54.150 253.670 54.140 253.660 54.140 ;
        POLYGON 254.255 54.150 254.265 54.150 254.265 54.140 ;
        RECT 254.265 54.140 254.730 54.150 ;
        RECT 252.625 54.135 253.670 54.140 ;
        POLYGON 252.625 54.135 252.675 54.135 252.675 54.100 ;
        RECT 252.675 54.100 253.670 54.135 ;
        POLYGON 252.675 54.100 252.690 54.100 252.690 54.090 ;
        RECT 252.690 54.090 253.670 54.100 ;
        POLYGON 252.695 54.090 252.725 54.090 252.725 54.070 ;
        RECT 252.725 54.070 253.670 54.090 ;
        RECT 245.365 54.045 246.485 54.070 ;
        RECT 244.100 53.990 244.735 54.040 ;
        POLYGON 244.735 54.040 244.770 54.040 244.735 53.990 ;
        POLYGON 245.300 54.040 245.300 54.030 245.290 54.030 ;
        RECT 245.300 54.030 246.485 54.045 ;
        POLYGON 245.290 54.030 245.290 53.990 245.260 53.990 ;
        RECT 245.290 54.025 246.485 54.030 ;
        POLYGON 246.485 54.070 246.535 54.070 246.485 54.025 ;
        POLYGON 252.725 54.070 252.785 54.070 252.785 54.030 ;
        RECT 252.785 54.035 253.670 54.070 ;
        POLYGON 253.670 54.140 253.795 54.035 253.670 54.035 ;
        POLYGON 254.265 54.140 254.305 54.140 254.305 54.105 ;
        RECT 254.305 54.130 254.730 54.140 ;
        POLYGON 254.730 54.325 254.910 54.130 254.730 54.130 ;
        POLYGON 255.510 54.325 255.520 54.325 255.520 54.315 ;
        RECT 255.520 54.315 256.195 54.325 ;
        POLYGON 255.520 54.315 255.550 54.315 255.550 54.275 ;
        RECT 255.550 54.295 256.195 54.315 ;
        POLYGON 256.195 54.360 256.245 54.295 256.195 54.295 ;
        POLYGON 257.060 54.360 257.100 54.360 257.100 54.310 ;
        RECT 257.100 54.340 258.140 54.360 ;
        POLYGON 258.140 54.370 258.155 54.340 258.140 54.340 ;
        POLYGON 259.470 54.370 259.485 54.370 259.485 54.340 ;
        RECT 259.485 54.340 261.015 54.370 ;
        RECT 257.100 54.310 258.155 54.340 ;
        POLYGON 257.100 54.310 257.105 54.310 257.105 54.300 ;
        RECT 257.105 54.295 258.155 54.310 ;
        RECT 255.550 54.275 256.245 54.295 ;
        POLYGON 255.550 54.275 255.655 54.275 255.655 54.145 ;
        RECT 255.655 54.260 256.245 54.275 ;
        POLYGON 256.245 54.295 256.275 54.260 256.245 54.260 ;
        POLYGON 257.105 54.295 257.130 54.295 257.130 54.260 ;
        RECT 257.130 54.260 258.155 54.295 ;
        RECT 255.655 54.255 256.275 54.260 ;
        POLYGON 256.275 54.260 256.280 54.255 256.275 54.255 ;
        POLYGON 257.130 54.260 257.135 54.260 257.135 54.255 ;
        RECT 257.135 54.255 258.155 54.260 ;
        RECT 255.655 54.145 256.280 54.255 ;
        POLYGON 255.655 54.145 255.665 54.145 255.665 54.130 ;
        RECT 255.665 54.130 256.280 54.145 ;
        RECT 254.305 54.105 254.910 54.130 ;
        POLYGON 254.910 54.130 254.935 54.105 254.910 54.105 ;
        POLYGON 255.665 54.130 255.680 54.130 255.680 54.115 ;
        RECT 255.680 54.115 256.280 54.130 ;
        POLYGON 255.680 54.115 255.685 54.115 255.685 54.105 ;
        RECT 255.685 54.105 256.280 54.115 ;
        POLYGON 254.305 54.105 254.310 54.105 254.310 54.095 ;
        RECT 254.310 54.095 254.935 54.105 ;
        POLYGON 254.935 54.105 254.940 54.095 254.935 54.095 ;
        POLYGON 255.685 54.105 255.695 54.105 255.695 54.095 ;
        RECT 255.695 54.095 256.280 54.105 ;
        POLYGON 254.310 54.095 254.325 54.095 254.325 54.085 ;
        RECT 254.325 54.085 254.940 54.095 ;
        POLYGON 254.325 54.085 254.375 54.085 254.375 54.035 ;
        RECT 254.375 54.070 254.940 54.085 ;
        POLYGON 254.940 54.095 254.965 54.070 254.940 54.070 ;
        POLYGON 255.695 54.095 255.710 54.095 255.710 54.070 ;
        RECT 255.710 54.070 256.280 54.095 ;
        RECT 254.375 54.035 254.965 54.070 ;
        RECT 252.785 54.030 253.795 54.035 ;
        POLYGON 252.785 54.030 252.790 54.030 252.790 54.025 ;
        RECT 252.790 54.025 253.795 54.030 ;
        RECT 245.290 53.990 246.400 54.025 ;
        RECT 244.100 53.980 244.725 53.990 ;
        POLYGON 244.725 53.990 244.735 53.990 244.725 53.980 ;
        POLYGON 245.260 53.990 245.260 53.980 245.255 53.980 ;
        RECT 245.260 53.980 246.400 53.990 ;
        RECT 244.100 53.975 244.695 53.980 ;
        RECT 242.490 53.935 243.235 53.970 ;
        RECT 240.150 53.925 241.235 53.935 ;
        POLYGON 240.095 53.925 240.095 53.875 240.080 53.875 ;
        RECT 240.095 53.875 241.235 53.925 ;
        RECT 229.305 53.770 233.415 53.870 ;
        POLYGON 233.415 53.870 233.430 53.870 233.415 53.770 ;
        POLYGON 236.330 53.870 236.330 53.775 236.305 53.775 ;
        RECT 236.330 53.775 238.340 53.875 ;
        RECT 229.305 53.075 233.305 53.770 ;
        POLYGON 206.510 52.800 206.535 52.800 206.535 52.615 ;
        RECT 206.535 52.645 222.225 52.800 ;
        POLYGON 222.225 53.075 222.230 52.645 222.225 52.645 ;
        RECT 206.535 52.590 222.230 52.645 ;
        POLYGON 229.230 53.065 229.230 52.725 229.205 52.725 ;
        RECT 229.230 52.980 233.305 53.075 ;
        POLYGON 233.305 53.770 233.415 53.770 233.305 52.980 ;
        POLYGON 236.305 53.770 236.305 53.735 236.295 53.735 ;
        RECT 236.305 53.735 238.340 53.775 ;
        POLYGON 236.295 53.735 236.295 52.980 236.150 52.980 ;
        RECT 236.295 53.545 238.340 53.735 ;
        POLYGON 238.340 53.875 238.435 53.875 238.340 53.545 ;
        POLYGON 240.080 53.875 240.080 53.580 239.995 53.580 ;
        RECT 240.080 53.840 241.235 53.875 ;
        POLYGON 241.235 53.935 241.270 53.935 241.235 53.845 ;
        POLYGON 242.430 53.935 242.430 53.845 242.385 53.845 ;
        RECT 242.430 53.845 243.235 53.935 ;
        POLYGON 243.235 53.970 243.300 53.970 243.235 53.845 ;
        POLYGON 244.055 53.970 244.055 53.910 244.015 53.910 ;
        RECT 244.055 53.940 244.695 53.975 ;
        POLYGON 244.695 53.980 244.725 53.980 244.695 53.940 ;
        POLYGON 245.255 53.980 245.255 53.975 245.250 53.975 ;
        RECT 245.255 53.975 246.400 53.980 ;
        POLYGON 245.250 53.975 245.250 53.940 245.225 53.940 ;
        RECT 245.250 53.940 246.400 53.975 ;
        POLYGON 246.400 54.025 246.485 54.025 246.400 53.940 ;
        POLYGON 252.790 54.025 252.820 54.025 252.820 54.005 ;
        RECT 252.820 54.010 253.795 54.025 ;
        POLYGON 253.795 54.035 253.820 54.010 253.795 54.010 ;
        POLYGON 254.375 54.035 254.400 54.035 254.400 54.010 ;
        RECT 254.400 54.010 254.965 54.035 ;
        RECT 252.820 54.005 253.820 54.010 ;
        POLYGON 252.820 54.005 252.905 54.005 252.905 53.940 ;
        RECT 252.905 53.940 253.820 54.005 ;
        RECT 244.055 53.910 244.615 53.940 ;
        POLYGON 244.015 53.910 244.015 53.880 244.000 53.880 ;
        RECT 244.015 53.880 244.615 53.910 ;
        POLYGON 244.000 53.880 244.000 53.845 243.975 53.845 ;
        RECT 244.000 53.845 244.615 53.880 ;
        RECT 240.080 53.610 241.150 53.840 ;
        POLYGON 241.150 53.840 241.235 53.840 241.150 53.615 ;
        POLYGON 242.385 53.845 242.385 53.815 242.370 53.815 ;
        RECT 242.385 53.840 243.230 53.845 ;
        POLYGON 243.230 53.845 243.235 53.845 243.230 53.840 ;
        RECT 242.385 53.820 243.220 53.840 ;
        POLYGON 243.220 53.840 243.230 53.840 243.220 53.820 ;
        POLYGON 243.975 53.840 243.975 53.820 243.960 53.820 ;
        RECT 243.975 53.830 244.615 53.845 ;
        POLYGON 244.615 53.940 244.695 53.940 244.615 53.830 ;
        POLYGON 245.225 53.940 245.225 53.895 245.190 53.895 ;
        RECT 245.225 53.900 246.355 53.940 ;
        POLYGON 246.355 53.940 246.400 53.940 246.355 53.900 ;
        POLYGON 252.905 53.940 252.940 53.940 252.940 53.915 ;
        RECT 252.940 53.915 253.820 53.940 ;
        POLYGON 253.820 54.010 253.925 53.915 253.820 53.915 ;
        POLYGON 254.400 54.010 254.445 54.010 254.445 53.970 ;
        RECT 254.445 53.970 254.965 54.010 ;
        POLYGON 254.445 53.970 254.495 53.970 254.495 53.915 ;
        RECT 254.495 53.930 254.965 53.970 ;
        POLYGON 254.965 54.070 255.080 53.930 254.965 53.930 ;
        POLYGON 255.710 54.070 255.765 54.070 255.765 53.995 ;
        RECT 255.765 54.060 256.280 54.070 ;
        POLYGON 256.280 54.255 256.410 54.060 256.280 54.060 ;
        POLYGON 257.135 54.255 257.235 54.255 257.235 54.105 ;
        RECT 257.235 54.180 258.155 54.255 ;
        POLYGON 258.155 54.340 258.245 54.180 258.155 54.180 ;
        POLYGON 259.485 54.340 259.495 54.340 259.495 54.325 ;
        RECT 259.495 54.325 261.015 54.340 ;
        POLYGON 259.495 54.325 259.570 54.325 259.570 54.185 ;
        RECT 259.570 54.195 261.015 54.325 ;
        POLYGON 261.015 54.375 261.085 54.195 261.015 54.195 ;
        POLYGON 263.090 54.375 263.145 54.375 263.145 54.235 ;
        RECT 263.145 54.235 265.730 54.375 ;
        POLYGON 265.730 54.735 265.900 54.235 265.730 54.235 ;
        POLYGON 270.035 54.735 270.100 54.735 270.100 54.565 ;
        RECT 270.100 54.565 276.895 54.735 ;
        POLYGON 270.100 54.565 270.200 54.565 270.200 54.245 ;
        RECT 270.200 54.350 276.895 54.565 ;
        POLYGON 276.895 54.895 277.050 54.350 276.895 54.350 ;
        RECT 270.200 54.235 277.050 54.350 ;
        POLYGON 263.145 54.235 263.160 54.235 263.160 54.195 ;
        RECT 263.160 54.195 265.900 54.235 ;
        RECT 259.570 54.180 261.085 54.195 ;
        RECT 257.235 54.105 258.245 54.180 ;
        POLYGON 257.235 54.105 257.260 54.105 257.260 54.065 ;
        RECT 257.260 54.090 258.245 54.105 ;
        POLYGON 258.245 54.180 258.295 54.090 258.245 54.090 ;
        POLYGON 259.570 54.180 259.595 54.180 259.595 54.140 ;
        RECT 259.595 54.140 261.085 54.180 ;
        POLYGON 259.595 54.140 259.620 54.140 259.620 54.095 ;
        RECT 259.620 54.090 261.085 54.140 ;
        RECT 257.260 54.065 258.295 54.090 ;
        POLYGON 258.295 54.090 258.310 54.065 258.295 54.065 ;
        POLYGON 259.620 54.090 259.630 54.090 259.630 54.070 ;
        RECT 259.630 54.065 261.085 54.090 ;
        RECT 257.260 54.060 258.310 54.065 ;
        RECT 255.765 53.995 256.410 54.060 ;
        POLYGON 255.765 53.995 255.805 53.995 255.805 53.945 ;
        RECT 255.805 53.955 256.410 53.995 ;
        POLYGON 256.410 54.060 256.485 53.955 256.410 53.955 ;
        POLYGON 257.260 54.060 257.305 54.060 257.305 53.995 ;
        RECT 257.305 53.995 258.310 54.060 ;
        POLYGON 257.305 53.995 257.325 53.995 257.325 53.955 ;
        RECT 257.325 53.955 258.310 53.995 ;
        RECT 255.805 53.945 256.485 53.955 ;
        POLYGON 255.805 53.945 255.815 53.945 255.815 53.930 ;
        RECT 255.815 53.930 256.485 53.945 ;
        POLYGON 256.485 53.955 256.505 53.930 256.485 53.930 ;
        POLYGON 257.325 53.955 257.330 53.955 257.330 53.950 ;
        RECT 257.330 53.950 258.310 53.955 ;
        POLYGON 257.330 53.950 257.340 53.950 257.340 53.930 ;
        RECT 257.340 53.930 258.310 53.950 ;
        RECT 254.495 53.915 255.080 53.930 ;
        POLYGON 252.940 53.915 252.965 53.915 252.965 53.900 ;
        RECT 252.965 53.900 253.925 53.915 ;
        POLYGON 253.925 53.915 253.935 53.900 253.925 53.900 ;
        POLYGON 254.495 53.915 254.510 53.915 254.510 53.900 ;
        RECT 254.510 53.900 255.080 53.915 ;
        RECT 245.225 53.895 246.265 53.900 ;
        POLYGON 245.190 53.895 245.190 53.830 245.145 53.830 ;
        RECT 245.190 53.830 246.265 53.895 ;
        RECT 243.975 53.820 244.605 53.830 ;
        POLYGON 244.605 53.830 244.615 53.830 244.605 53.820 ;
        POLYGON 245.145 53.830 245.145 53.825 245.140 53.825 ;
        RECT 245.145 53.825 246.265 53.830 ;
        RECT 242.385 53.815 243.170 53.820 ;
        POLYGON 242.370 53.815 242.370 53.745 242.340 53.745 ;
        RECT 242.370 53.745 243.170 53.815 ;
        POLYGON 242.340 53.745 242.340 53.655 242.300 53.655 ;
        RECT 242.340 53.710 243.170 53.745 ;
        POLYGON 243.170 53.820 243.220 53.820 243.170 53.710 ;
        POLYGON 243.960 53.820 243.960 53.710 243.895 53.710 ;
        RECT 243.960 53.760 244.565 53.820 ;
        POLYGON 244.565 53.820 244.605 53.820 244.565 53.760 ;
        POLYGON 245.140 53.820 245.140 53.760 245.095 53.760 ;
        RECT 245.140 53.810 246.265 53.825 ;
        POLYGON 246.265 53.900 246.355 53.900 246.265 53.810 ;
        POLYGON 252.965 53.900 252.985 53.900 252.985 53.885 ;
        RECT 252.985 53.885 253.935 53.900 ;
        POLYGON 252.985 53.885 253.075 53.885 253.075 53.810 ;
        RECT 253.075 53.810 253.935 53.885 ;
        RECT 245.140 53.760 246.175 53.810 ;
        RECT 243.960 53.720 244.535 53.760 ;
        POLYGON 244.535 53.760 244.565 53.760 244.535 53.720 ;
        POLYGON 245.095 53.760 245.095 53.720 245.070 53.720 ;
        RECT 245.095 53.720 246.175 53.760 ;
        RECT 243.960 53.710 244.490 53.720 ;
        RECT 242.340 53.655 243.115 53.710 ;
        POLYGON 242.300 53.655 242.300 53.615 242.280 53.615 ;
        RECT 242.300 53.615 243.115 53.655 ;
        RECT 240.080 53.580 241.090 53.610 ;
        POLYGON 239.995 53.580 239.995 53.560 239.990 53.560 ;
        RECT 239.995 53.560 241.090 53.580 ;
        POLYGON 239.990 53.560 239.990 53.545 239.985 53.545 ;
        RECT 239.990 53.545 241.090 53.560 ;
        RECT 236.295 53.350 238.295 53.545 ;
        POLYGON 238.295 53.545 238.340 53.545 238.295 53.350 ;
        POLYGON 239.985 53.540 239.985 53.350 239.935 53.350 ;
        RECT 239.985 53.435 241.090 53.545 ;
        POLYGON 241.090 53.610 241.150 53.610 241.090 53.435 ;
        POLYGON 242.280 53.610 242.280 53.510 242.235 53.510 ;
        RECT 242.280 53.600 243.115 53.615 ;
        POLYGON 243.115 53.710 243.170 53.710 243.115 53.600 ;
        POLYGON 243.895 53.710 243.895 53.675 243.875 53.675 ;
        RECT 243.895 53.675 244.490 53.710 ;
        POLYGON 243.875 53.675 243.875 53.660 243.870 53.660 ;
        RECT 243.875 53.660 244.490 53.675 ;
        POLYGON 243.870 53.660 243.870 53.600 243.835 53.600 ;
        RECT 243.870 53.650 244.490 53.660 ;
        POLYGON 244.490 53.720 244.535 53.720 244.490 53.650 ;
        POLYGON 245.070 53.720 245.070 53.715 245.065 53.715 ;
        RECT 245.070 53.715 246.175 53.720 ;
        POLYGON 246.175 53.810 246.265 53.810 246.175 53.715 ;
        POLYGON 253.075 53.810 253.095 53.810 253.095 53.795 ;
        RECT 253.095 53.795 253.935 53.810 ;
        POLYGON 253.095 53.795 253.195 53.795 253.195 53.715 ;
        RECT 253.195 53.780 253.935 53.795 ;
        POLYGON 253.935 53.900 254.065 53.780 253.935 53.780 ;
        POLYGON 254.510 53.900 254.570 53.900 254.570 53.840 ;
        RECT 254.570 53.870 255.080 53.900 ;
        POLYGON 255.080 53.930 255.135 53.870 255.080 53.870 ;
        POLYGON 255.815 53.930 255.825 53.930 255.825 53.920 ;
        RECT 255.825 53.920 256.505 53.930 ;
        POLYGON 255.825 53.920 255.830 53.920 255.830 53.910 ;
        RECT 255.830 53.910 256.505 53.920 ;
        POLYGON 255.830 53.910 255.855 53.910 255.855 53.870 ;
        RECT 255.855 53.895 256.505 53.910 ;
        POLYGON 256.505 53.930 256.525 53.895 256.505 53.895 ;
        POLYGON 257.340 53.930 257.360 53.930 257.360 53.900 ;
        RECT 257.360 53.895 258.310 53.930 ;
        RECT 255.855 53.870 256.525 53.895 ;
        RECT 254.570 53.840 255.135 53.870 ;
        POLYGON 254.570 53.840 254.625 53.840 254.625 53.780 ;
        RECT 254.625 53.835 255.135 53.840 ;
        POLYGON 255.135 53.870 255.160 53.835 255.135 53.835 ;
        POLYGON 255.855 53.870 255.880 53.870 255.880 53.835 ;
        RECT 255.880 53.835 256.525 53.870 ;
        RECT 254.625 53.820 255.160 53.835 ;
        POLYGON 255.160 53.835 255.175 53.820 255.160 53.820 ;
        POLYGON 255.880 53.835 255.890 53.835 255.890 53.820 ;
        RECT 255.890 53.825 256.525 53.835 ;
        POLYGON 256.525 53.895 256.570 53.825 256.525 53.825 ;
        POLYGON 257.360 53.895 257.390 53.895 257.390 53.855 ;
        RECT 257.390 53.855 258.310 53.895 ;
        POLYGON 257.390 53.855 257.405 53.855 257.405 53.825 ;
        RECT 257.405 53.825 258.310 53.855 ;
        RECT 255.890 53.820 256.570 53.825 ;
        RECT 254.625 53.780 255.175 53.820 ;
        RECT 253.195 53.770 254.065 53.780 ;
        POLYGON 254.065 53.780 254.075 53.770 254.065 53.770 ;
        POLYGON 254.625 53.780 254.635 53.780 254.635 53.770 ;
        RECT 254.635 53.770 255.175 53.780 ;
        RECT 253.195 53.715 254.075 53.770 ;
        POLYGON 245.065 53.715 245.065 53.680 245.040 53.680 ;
        RECT 245.065 53.710 246.175 53.715 ;
        RECT 245.065 53.680 246.140 53.710 ;
        POLYGON 245.040 53.680 245.040 53.660 245.025 53.660 ;
        RECT 245.040 53.670 246.140 53.680 ;
        POLYGON 246.140 53.710 246.175 53.710 246.140 53.670 ;
        POLYGON 253.195 53.715 253.245 53.715 253.245 53.675 ;
        RECT 253.245 53.675 254.075 53.715 ;
        POLYGON 253.245 53.675 253.250 53.675 253.250 53.670 ;
        RECT 253.250 53.670 254.075 53.675 ;
        RECT 245.040 53.665 246.130 53.670 ;
        POLYGON 246.130 53.670 246.140 53.670 246.130 53.665 ;
        POLYGON 253.250 53.670 253.255 53.670 253.255 53.665 ;
        RECT 253.255 53.665 254.075 53.670 ;
        RECT 245.040 53.660 246.025 53.665 ;
        POLYGON 245.025 53.660 245.025 53.650 245.020 53.650 ;
        RECT 245.025 53.650 246.025 53.660 ;
        RECT 243.870 53.615 244.465 53.650 ;
        POLYGON 244.465 53.650 244.490 53.650 244.465 53.615 ;
        POLYGON 245.020 53.650 245.020 53.615 244.995 53.615 ;
        RECT 245.020 53.615 246.025 53.650 ;
        RECT 243.870 53.600 244.410 53.615 ;
        RECT 242.280 53.595 243.110 53.600 ;
        POLYGON 243.110 53.600 243.115 53.600 243.110 53.595 ;
        RECT 242.280 53.565 243.100 53.595 ;
        POLYGON 243.100 53.595 243.110 53.595 243.100 53.565 ;
        POLYGON 243.835 53.595 243.835 53.565 243.815 53.565 ;
        RECT 243.835 53.565 244.410 53.600 ;
        RECT 242.280 53.510 243.065 53.565 ;
        POLYGON 242.235 53.510 242.235 53.435 242.200 53.435 ;
        RECT 242.235 53.495 243.065 53.510 ;
        POLYGON 243.065 53.565 243.100 53.565 243.065 53.495 ;
        POLYGON 243.815 53.565 243.815 53.530 243.795 53.530 ;
        RECT 243.815 53.530 244.410 53.565 ;
        POLYGON 244.410 53.615 244.465 53.615 244.410 53.530 ;
        POLYGON 244.995 53.610 244.995 53.530 244.945 53.530 ;
        RECT 244.995 53.545 246.025 53.615 ;
        POLYGON 246.025 53.665 246.130 53.665 246.025 53.545 ;
        POLYGON 253.255 53.665 253.275 53.665 253.275 53.650 ;
        RECT 253.275 53.655 254.075 53.665 ;
        POLYGON 254.075 53.770 254.185 53.655 254.075 53.655 ;
        POLYGON 254.635 53.770 254.705 53.770 254.705 53.700 ;
        RECT 254.705 53.725 255.175 53.770 ;
        POLYGON 255.175 53.820 255.245 53.725 255.175 53.725 ;
        POLYGON 255.890 53.820 255.940 53.820 255.940 53.750 ;
        RECT 255.940 53.750 256.570 53.820 ;
        POLYGON 255.940 53.750 255.955 53.750 255.955 53.725 ;
        RECT 255.955 53.725 256.570 53.750 ;
        RECT 254.705 53.700 255.245 53.725 ;
        POLYGON 254.705 53.700 254.725 53.700 254.725 53.675 ;
        RECT 254.725 53.675 255.245 53.700 ;
        POLYGON 254.725 53.675 254.730 53.675 254.730 53.670 ;
        RECT 254.730 53.670 255.245 53.675 ;
        POLYGON 254.730 53.670 254.740 53.670 254.740 53.655 ;
        RECT 254.740 53.655 255.245 53.670 ;
        RECT 253.275 53.650 254.185 53.655 ;
        POLYGON 253.275 53.650 253.390 53.650 253.390 53.545 ;
        RECT 253.390 53.545 254.185 53.650 ;
        RECT 244.995 53.530 246.015 53.545 ;
        POLYGON 246.015 53.545 246.025 53.545 246.015 53.530 ;
        POLYGON 253.390 53.545 253.405 53.545 253.405 53.530 ;
        RECT 253.405 53.530 254.185 53.545 ;
        POLYGON 254.185 53.655 254.305 53.530 254.185 53.530 ;
        POLYGON 254.740 53.655 254.805 53.655 254.805 53.590 ;
        RECT 254.805 53.630 255.245 53.655 ;
        POLYGON 255.245 53.725 255.320 53.630 255.245 53.630 ;
        POLYGON 255.955 53.725 255.960 53.725 255.960 53.720 ;
        RECT 255.960 53.720 256.570 53.725 ;
        POLYGON 255.960 53.720 256.015 53.720 256.015 53.635 ;
        RECT 256.015 53.630 256.570 53.720 ;
        RECT 254.805 53.590 255.320 53.630 ;
        POLYGON 255.320 53.630 255.345 53.590 255.320 53.590 ;
        POLYGON 256.015 53.630 256.035 53.630 256.035 53.605 ;
        RECT 256.035 53.605 256.570 53.630 ;
        POLYGON 256.035 53.605 256.040 53.605 256.040 53.595 ;
        RECT 256.040 53.595 256.570 53.605 ;
        POLYGON 256.570 53.825 256.710 53.595 256.570 53.595 ;
        POLYGON 257.405 53.825 257.425 53.825 257.425 53.795 ;
        RECT 257.425 53.810 258.310 53.825 ;
        POLYGON 258.310 54.065 258.445 53.810 258.310 53.810 ;
        POLYGON 259.630 54.065 259.695 54.065 259.695 53.940 ;
        RECT 259.695 54.000 261.085 54.065 ;
        POLYGON 261.085 54.195 261.165 54.000 261.085 54.000 ;
        POLYGON 263.160 54.195 263.215 54.195 263.215 54.060 ;
        RECT 263.215 54.170 265.900 54.195 ;
        POLYGON 265.900 54.235 265.920 54.170 265.900 54.170 ;
        POLYGON 270.200 54.235 270.220 54.235 270.220 54.180 ;
        RECT 270.220 54.170 277.050 54.235 ;
        RECT 263.215 54.075 265.920 54.170 ;
        POLYGON 265.920 54.170 265.950 54.075 265.920 54.075 ;
        POLYGON 270.220 54.170 270.250 54.170 270.250 54.085 ;
        RECT 270.250 54.075 277.050 54.170 ;
        RECT 263.215 54.060 265.950 54.075 ;
        POLYGON 263.215 54.060 263.235 54.060 263.235 54.000 ;
        RECT 263.235 54.000 265.950 54.060 ;
        RECT 259.695 53.970 261.165 54.000 ;
        POLYGON 261.165 54.000 261.175 53.970 261.165 53.970 ;
        POLYGON 263.235 54.000 263.245 54.000 263.245 53.970 ;
        RECT 263.245 53.970 265.950 54.000 ;
        RECT 259.695 53.940 261.175 53.970 ;
        POLYGON 259.695 53.940 259.750 53.940 259.750 53.810 ;
        RECT 259.750 53.810 261.175 53.940 ;
        RECT 257.425 53.795 258.445 53.810 ;
        POLYGON 257.425 53.795 257.440 53.795 257.440 53.775 ;
        RECT 257.440 53.780 258.445 53.795 ;
        POLYGON 258.445 53.810 258.460 53.780 258.445 53.780 ;
        POLYGON 259.750 53.810 259.760 53.810 259.760 53.785 ;
        RECT 259.760 53.780 261.175 53.810 ;
        RECT 257.440 53.775 258.460 53.780 ;
        POLYGON 257.440 53.775 257.445 53.775 257.445 53.760 ;
        RECT 257.445 53.760 258.460 53.775 ;
        POLYGON 257.445 53.760 257.525 53.760 257.525 53.620 ;
        RECT 257.525 53.620 258.460 53.760 ;
        POLYGON 257.525 53.620 257.535 53.620 257.535 53.600 ;
        RECT 257.535 53.595 258.460 53.620 ;
        POLYGON 258.460 53.780 258.545 53.595 258.460 53.595 ;
        POLYGON 259.760 53.780 259.785 53.780 259.785 53.730 ;
        RECT 259.785 53.760 261.175 53.780 ;
        POLYGON 261.175 53.970 261.250 53.760 261.175 53.760 ;
        POLYGON 263.245 53.970 263.315 53.970 263.315 53.760 ;
        RECT 263.315 53.760 265.950 53.970 ;
        RECT 259.785 53.730 261.250 53.760 ;
        POLYGON 259.785 53.730 259.820 53.730 259.820 53.640 ;
        RECT 259.820 53.640 261.250 53.730 ;
        POLYGON 259.820 53.640 259.835 53.640 259.835 53.600 ;
        RECT 259.835 53.615 261.250 53.640 ;
        POLYGON 261.250 53.760 261.300 53.615 261.250 53.615 ;
        POLYGON 263.315 53.760 263.360 53.760 263.360 53.625 ;
        RECT 263.360 53.660 265.950 53.760 ;
        POLYGON 265.950 54.075 266.075 53.660 265.950 53.660 ;
        POLYGON 270.250 54.075 270.295 54.075 270.295 53.945 ;
        RECT 270.295 53.945 277.050 54.075 ;
        POLYGON 270.295 53.945 270.365 53.945 270.365 53.675 ;
        RECT 270.365 53.680 277.050 53.945 ;
        POLYGON 277.050 54.350 277.205 53.680 277.050 53.680 ;
        RECT 270.365 53.660 277.205 53.680 ;
        RECT 263.360 53.615 266.075 53.660 ;
        RECT 259.835 53.595 261.300 53.615 ;
        RECT 256.040 53.590 256.710 53.595 ;
        POLYGON 254.805 53.590 254.815 53.590 254.815 53.575 ;
        RECT 254.815 53.575 255.345 53.590 ;
        POLYGON 254.815 53.575 254.850 53.575 254.850 53.530 ;
        RECT 254.850 53.530 255.345 53.575 ;
        POLYGON 243.795 53.530 243.795 53.500 243.780 53.500 ;
        RECT 243.795 53.500 244.385 53.530 ;
        RECT 242.235 53.435 243.040 53.495 ;
        POLYGON 243.040 53.495 243.065 53.495 243.040 53.435 ;
        POLYGON 243.780 53.495 243.780 53.460 243.760 53.460 ;
        RECT 243.780 53.490 244.385 53.500 ;
        POLYGON 244.385 53.530 244.410 53.530 244.385 53.495 ;
        POLYGON 244.945 53.530 244.945 53.500 244.925 53.500 ;
        RECT 244.945 53.500 245.955 53.530 ;
        RECT 243.780 53.460 244.320 53.490 ;
        POLYGON 243.760 53.460 243.760 53.435 243.745 53.435 ;
        RECT 243.760 53.435 244.320 53.460 ;
        RECT 239.985 53.380 241.070 53.435 ;
        POLYGON 241.070 53.435 241.090 53.435 241.070 53.380 ;
        POLYGON 242.200 53.435 242.200 53.400 242.185 53.400 ;
        RECT 242.200 53.410 243.030 53.435 ;
        POLYGON 243.030 53.435 243.040 53.435 243.030 53.410 ;
        POLYGON 243.745 53.430 243.745 53.410 243.735 53.410 ;
        RECT 243.745 53.410 244.320 53.435 ;
        RECT 242.200 53.400 242.995 53.410 ;
        POLYGON 242.185 53.400 242.185 53.380 242.175 53.380 ;
        RECT 242.185 53.380 242.995 53.400 ;
        RECT 239.985 53.350 241.005 53.380 ;
        RECT 236.295 53.000 238.215 53.350 ;
        POLYGON 238.215 53.350 238.295 53.350 238.215 53.000 ;
        POLYGON 239.935 53.345 239.935 53.230 239.905 53.230 ;
        RECT 239.935 53.230 241.005 53.350 ;
        POLYGON 239.905 53.230 239.905 53.000 239.855 53.000 ;
        RECT 239.905 53.145 241.005 53.230 ;
        POLYGON 241.005 53.380 241.070 53.380 241.005 53.145 ;
        POLYGON 242.175 53.375 242.175 53.200 242.105 53.200 ;
        RECT 242.175 53.340 242.995 53.380 ;
        POLYGON 242.995 53.410 243.030 53.410 242.995 53.340 ;
        POLYGON 243.735 53.410 243.735 53.345 243.700 53.345 ;
        RECT 243.735 53.390 244.320 53.410 ;
        POLYGON 244.320 53.490 244.385 53.490 244.320 53.390 ;
        POLYGON 244.925 53.495 244.925 53.440 244.890 53.440 ;
        RECT 244.925 53.465 245.955 53.500 ;
        POLYGON 245.955 53.530 246.015 53.530 245.955 53.465 ;
        POLYGON 253.405 53.530 253.475 53.530 253.475 53.465 ;
        RECT 253.475 53.520 254.305 53.530 ;
        POLYGON 254.305 53.530 254.310 53.520 254.305 53.520 ;
        POLYGON 254.850 53.530 254.860 53.530 254.860 53.520 ;
        RECT 254.860 53.520 255.345 53.530 ;
        RECT 253.475 53.505 254.310 53.520 ;
        POLYGON 254.310 53.520 254.325 53.505 254.310 53.505 ;
        POLYGON 254.860 53.520 254.870 53.520 254.870 53.510 ;
        RECT 254.870 53.515 255.345 53.520 ;
        POLYGON 255.345 53.590 255.400 53.515 255.345 53.515 ;
        POLYGON 256.040 53.590 256.065 53.590 256.065 53.555 ;
        RECT 256.065 53.585 256.710 53.590 ;
        POLYGON 256.710 53.595 256.715 53.585 256.710 53.585 ;
        POLYGON 257.535 53.595 257.540 53.595 257.540 53.590 ;
        RECT 257.540 53.585 258.545 53.595 ;
        RECT 256.065 53.555 256.715 53.585 ;
        POLYGON 256.065 53.555 256.080 53.555 256.080 53.530 ;
        RECT 256.080 53.530 256.715 53.555 ;
        POLYGON 256.080 53.530 256.085 53.530 256.085 53.520 ;
        RECT 256.085 53.515 256.715 53.530 ;
        RECT 254.870 53.505 255.400 53.515 ;
        RECT 253.475 53.465 254.325 53.505 ;
        RECT 244.925 53.440 245.895 53.465 ;
        POLYGON 244.890 53.440 244.890 53.410 244.875 53.410 ;
        RECT 244.890 53.410 245.895 53.440 ;
        POLYGON 244.875 53.410 244.875 53.395 244.865 53.395 ;
        RECT 244.875 53.395 245.895 53.410 ;
        POLYGON 244.865 53.395 244.865 53.390 244.860 53.390 ;
        RECT 244.865 53.390 245.895 53.395 ;
        POLYGON 245.895 53.465 245.955 53.465 245.895 53.390 ;
        POLYGON 253.475 53.465 253.515 53.465 253.515 53.430 ;
        RECT 253.515 53.430 254.325 53.465 ;
        POLYGON 253.515 53.430 253.535 53.430 253.535 53.415 ;
        RECT 253.535 53.415 254.325 53.430 ;
        POLYGON 253.535 53.415 253.555 53.415 253.555 53.395 ;
        RECT 253.555 53.390 254.325 53.415 ;
        RECT 243.735 53.345 244.295 53.390 ;
        POLYGON 244.295 53.390 244.320 53.390 244.295 53.345 ;
        POLYGON 244.860 53.385 244.860 53.345 244.835 53.345 ;
        RECT 244.860 53.375 245.885 53.390 ;
        POLYGON 245.885 53.390 245.895 53.390 245.885 53.375 ;
        POLYGON 253.555 53.390 253.570 53.390 253.570 53.375 ;
        RECT 253.570 53.375 254.325 53.390 ;
        RECT 244.860 53.345 245.780 53.375 ;
        RECT 242.175 53.280 242.975 53.340 ;
        POLYGON 242.975 53.340 242.995 53.340 242.975 53.280 ;
        POLYGON 243.700 53.340 243.700 53.335 243.695 53.335 ;
        RECT 243.700 53.335 244.265 53.345 ;
        POLYGON 243.695 53.335 243.695 53.280 243.670 53.280 ;
        RECT 243.695 53.295 244.265 53.335 ;
        POLYGON 244.265 53.345 244.295 53.345 244.265 53.295 ;
        POLYGON 244.835 53.340 244.835 53.295 244.810 53.295 ;
        RECT 244.835 53.295 245.780 53.345 ;
        RECT 243.695 53.280 244.240 53.295 ;
        RECT 242.175 53.240 242.955 53.280 ;
        POLYGON 242.955 53.280 242.975 53.280 242.955 53.240 ;
        POLYGON 243.670 53.280 243.670 53.245 243.655 53.245 ;
        RECT 243.670 53.250 244.240 53.280 ;
        POLYGON 244.240 53.295 244.265 53.295 244.240 53.250 ;
        POLYGON 244.810 53.295 244.810 53.250 244.785 53.250 ;
        RECT 244.810 53.250 245.780 53.295 ;
        RECT 243.670 53.245 244.220 53.250 ;
        RECT 242.175 53.220 242.950 53.240 ;
        POLYGON 242.950 53.240 242.955 53.240 242.950 53.220 ;
        POLYGON 243.655 53.240 243.655 53.235 243.650 53.235 ;
        RECT 243.655 53.235 244.220 53.245 ;
        POLYGON 243.650 53.235 243.650 53.220 243.640 53.220 ;
        RECT 243.650 53.220 244.220 53.235 ;
        RECT 242.175 53.200 242.910 53.220 ;
        POLYGON 242.105 53.195 242.105 53.145 242.085 53.145 ;
        RECT 242.105 53.145 242.910 53.200 ;
        RECT 239.905 53.120 240.995 53.145 ;
        POLYGON 240.995 53.145 241.005 53.145 240.995 53.120 ;
        POLYGON 242.085 53.145 242.085 53.120 242.075 53.120 ;
        RECT 242.085 53.130 242.910 53.145 ;
        POLYGON 242.910 53.220 242.945 53.220 242.910 53.130 ;
        POLYGON 243.640 53.220 243.640 53.130 243.600 53.130 ;
        RECT 243.640 53.215 244.220 53.220 ;
        POLYGON 244.220 53.250 244.240 53.250 244.220 53.215 ;
        POLYGON 244.785 53.250 244.785 53.225 244.770 53.225 ;
        RECT 244.785 53.240 245.780 53.250 ;
        POLYGON 245.780 53.375 245.885 53.375 245.780 53.240 ;
        POLYGON 253.570 53.375 253.705 53.375 253.705 53.240 ;
        RECT 253.705 53.365 254.325 53.375 ;
        POLYGON 254.325 53.505 254.445 53.365 254.325 53.365 ;
        POLYGON 254.870 53.505 254.920 53.505 254.920 53.455 ;
        RECT 254.920 53.455 255.400 53.505 ;
        POLYGON 254.920 53.455 254.965 53.455 254.965 53.400 ;
        RECT 254.965 53.400 255.400 53.455 ;
        POLYGON 255.400 53.515 255.480 53.400 255.400 53.400 ;
        POLYGON 256.085 53.515 256.155 53.515 256.155 53.400 ;
        RECT 256.155 53.510 256.715 53.515 ;
        POLYGON 256.715 53.585 256.755 53.510 256.715 53.510 ;
        POLYGON 257.540 53.585 257.585 53.585 257.585 53.510 ;
        RECT 257.585 53.510 258.545 53.585 ;
        RECT 256.155 53.490 256.755 53.510 ;
        POLYGON 256.755 53.510 256.765 53.490 256.755 53.490 ;
        POLYGON 257.585 53.510 257.590 53.510 257.590 53.495 ;
        RECT 257.590 53.495 258.545 53.510 ;
        POLYGON 258.545 53.595 258.595 53.495 258.545 53.495 ;
        POLYGON 259.835 53.595 259.855 53.595 259.855 53.555 ;
        RECT 259.855 53.555 261.300 53.595 ;
        POLYGON 259.855 53.555 259.875 53.555 259.875 53.510 ;
        RECT 259.875 53.510 261.300 53.555 ;
        POLYGON 259.875 53.510 259.880 53.510 259.880 53.495 ;
        RECT 259.880 53.495 261.300 53.510 ;
        RECT 257.590 53.490 258.595 53.495 ;
        RECT 256.155 53.400 256.765 53.490 ;
        POLYGON 254.965 53.400 254.995 53.400 254.995 53.365 ;
        RECT 254.995 53.380 255.480 53.400 ;
        POLYGON 255.480 53.400 255.495 53.380 255.480 53.380 ;
        POLYGON 256.155 53.400 256.165 53.400 256.165 53.385 ;
        RECT 256.165 53.380 256.765 53.400 ;
        RECT 254.995 53.365 255.495 53.380 ;
        RECT 253.705 53.265 254.445 53.365 ;
        POLYGON 254.445 53.365 254.525 53.265 254.445 53.265 ;
        POLYGON 254.995 53.365 255.000 53.365 255.000 53.360 ;
        RECT 255.000 53.360 255.495 53.365 ;
        POLYGON 255.000 53.360 255.020 53.360 255.020 53.335 ;
        RECT 255.020 53.345 255.495 53.360 ;
        POLYGON 255.495 53.380 255.520 53.345 255.495 53.345 ;
        POLYGON 256.165 53.380 256.175 53.380 256.175 53.370 ;
        RECT 256.175 53.370 256.765 53.380 ;
        POLYGON 256.175 53.370 256.190 53.370 256.190 53.345 ;
        RECT 256.190 53.345 256.765 53.370 ;
        RECT 255.020 53.335 255.520 53.345 ;
        POLYGON 255.020 53.335 255.070 53.335 255.070 53.265 ;
        RECT 255.070 53.295 255.520 53.335 ;
        POLYGON 255.520 53.345 255.550 53.295 255.520 53.295 ;
        POLYGON 256.190 53.345 256.215 53.345 256.215 53.295 ;
        RECT 256.215 53.330 256.765 53.345 ;
        POLYGON 256.765 53.490 256.855 53.330 256.765 53.330 ;
        POLYGON 257.590 53.490 257.625 53.490 257.625 53.435 ;
        RECT 257.625 53.435 258.595 53.490 ;
        POLYGON 257.625 53.435 257.670 53.435 257.670 53.345 ;
        RECT 257.670 53.335 258.595 53.435 ;
        POLYGON 257.670 53.335 257.675 53.335 257.675 53.330 ;
        RECT 257.675 53.330 258.595 53.335 ;
        POLYGON 258.595 53.495 258.665 53.330 258.595 53.330 ;
        POLYGON 259.880 53.495 259.935 53.495 259.935 53.335 ;
        RECT 259.935 53.330 261.300 53.495 ;
        RECT 256.215 53.295 256.855 53.330 ;
        RECT 253.705 53.260 254.525 53.265 ;
        POLYGON 254.525 53.265 254.530 53.260 254.525 53.260 ;
        RECT 255.070 53.260 255.550 53.295 ;
        RECT 253.705 53.240 254.530 53.260 ;
        RECT 244.785 53.225 245.750 53.240 ;
        POLYGON 244.770 53.225 244.770 53.215 244.765 53.215 ;
        RECT 244.770 53.215 245.750 53.225 ;
        RECT 243.640 53.165 244.190 53.215 ;
        POLYGON 244.190 53.215 244.220 53.215 244.190 53.165 ;
        POLYGON 244.765 53.215 244.765 53.165 244.740 53.165 ;
        RECT 244.765 53.200 245.750 53.215 ;
        POLYGON 245.750 53.240 245.780 53.240 245.750 53.200 ;
        POLYGON 253.705 53.240 253.745 53.240 253.745 53.200 ;
        RECT 253.745 53.210 254.530 53.240 ;
        POLYGON 254.530 53.260 254.570 53.210 254.530 53.210 ;
        POLYGON 255.070 53.260 255.090 53.260 255.090 53.240 ;
        RECT 255.090 53.240 255.550 53.260 ;
        POLYGON 255.090 53.240 255.110 53.240 255.110 53.210 ;
        RECT 255.110 53.210 255.550 53.240 ;
        RECT 253.745 53.200 254.570 53.210 ;
        RECT 244.765 53.165 245.715 53.200 ;
        RECT 243.640 53.130 244.155 53.165 ;
        RECT 242.085 53.120 242.880 53.130 ;
        RECT 239.905 53.000 240.930 53.120 ;
        RECT 236.295 52.980 238.190 53.000 ;
        RECT 229.230 52.840 233.290 52.980 ;
        POLYGON 233.290 52.980 233.305 52.980 233.290 52.840 ;
        POLYGON 236.150 52.980 236.150 52.955 236.145 52.955 ;
        RECT 236.150 52.955 238.190 52.980 ;
        POLYGON 236.145 52.955 236.145 52.840 236.130 52.840 ;
        RECT 236.145 52.870 238.190 52.955 ;
        POLYGON 238.190 53.000 238.215 53.000 238.190 52.870 ;
        POLYGON 239.855 52.995 239.855 52.875 239.830 52.875 ;
        RECT 239.855 52.890 240.930 53.000 ;
        POLYGON 240.930 53.120 240.995 53.120 240.930 52.890 ;
        POLYGON 242.075 53.120 242.075 53.055 242.050 53.055 ;
        RECT 242.075 53.055 242.880 53.120 ;
        POLYGON 242.050 53.055 242.050 52.895 241.995 52.895 ;
        RECT 242.050 53.045 242.880 53.055 ;
        POLYGON 242.880 53.130 242.910 53.130 242.880 53.045 ;
        POLYGON 243.600 53.130 243.600 53.045 243.560 53.045 ;
        RECT 243.600 53.100 244.155 53.130 ;
        POLYGON 244.155 53.165 244.190 53.165 244.155 53.100 ;
        POLYGON 244.740 53.165 244.740 53.135 244.725 53.135 ;
        RECT 244.740 53.150 245.715 53.165 ;
        POLYGON 245.715 53.200 245.750 53.200 245.715 53.150 ;
        POLYGON 253.745 53.200 253.770 53.200 253.770 53.175 ;
        RECT 253.770 53.175 254.570 53.200 ;
        POLYGON 253.770 53.175 253.785 53.175 253.785 53.155 ;
        RECT 253.785 53.150 254.570 53.175 ;
        RECT 244.740 53.135 245.670 53.150 ;
        POLYGON 244.725 53.135 244.725 53.100 244.705 53.100 ;
        RECT 244.725 53.100 245.670 53.135 ;
        RECT 243.600 53.050 244.130 53.100 ;
        POLYGON 244.130 53.100 244.155 53.100 244.130 53.050 ;
        POLYGON 244.705 53.100 244.705 53.050 244.680 53.050 ;
        RECT 244.705 53.090 245.670 53.100 ;
        POLYGON 245.670 53.150 245.715 53.150 245.670 53.090 ;
        POLYGON 253.785 53.150 253.820 53.150 253.820 53.115 ;
        RECT 253.820 53.115 254.570 53.150 ;
        POLYGON 253.820 53.115 253.840 53.115 253.840 53.090 ;
        RECT 253.840 53.090 254.570 53.115 ;
        RECT 244.705 53.050 245.620 53.090 ;
        RECT 243.600 53.045 244.105 53.050 ;
        RECT 242.050 52.990 242.860 53.045 ;
        POLYGON 242.860 53.045 242.880 53.045 242.860 52.990 ;
        POLYGON 243.560 53.040 243.560 52.990 243.535 52.990 ;
        RECT 243.560 53.005 244.105 53.045 ;
        POLYGON 244.105 53.050 244.130 53.050 244.105 53.005 ;
        POLYGON 244.680 53.045 244.680 53.005 244.660 53.005 ;
        RECT 244.680 53.025 245.620 53.050 ;
        POLYGON 245.620 53.090 245.670 53.090 245.620 53.025 ;
        POLYGON 253.840 53.090 253.895 53.090 253.895 53.025 ;
        RECT 253.895 53.030 254.570 53.090 ;
        POLYGON 254.570 53.210 254.705 53.030 254.570 53.030 ;
        POLYGON 255.110 53.210 255.160 53.210 255.160 53.145 ;
        RECT 255.160 53.145 255.550 53.210 ;
        POLYGON 255.160 53.145 255.175 53.145 255.175 53.125 ;
        RECT 255.175 53.130 255.550 53.145 ;
        POLYGON 255.550 53.295 255.655 53.130 255.550 53.130 ;
        POLYGON 256.215 53.295 256.270 53.295 256.270 53.195 ;
        RECT 256.270 53.250 256.855 53.295 ;
        POLYGON 256.855 53.330 256.895 53.250 256.855 53.250 ;
        POLYGON 257.675 53.330 257.680 53.330 257.680 53.325 ;
        RECT 257.680 53.325 258.665 53.330 ;
        POLYGON 257.680 53.325 257.715 53.325 257.715 53.250 ;
        RECT 257.715 53.250 258.665 53.325 ;
        RECT 256.270 53.195 256.895 53.250 ;
        POLYGON 256.270 53.195 256.280 53.195 256.280 53.180 ;
        RECT 256.280 53.180 256.895 53.195 ;
        POLYGON 256.280 53.180 256.285 53.180 256.285 53.170 ;
        RECT 256.285 53.170 256.895 53.180 ;
        POLYGON 256.285 53.170 256.305 53.170 256.305 53.135 ;
        RECT 256.305 53.130 256.895 53.170 ;
        RECT 255.175 53.125 255.655 53.130 ;
        POLYGON 255.175 53.125 255.210 53.125 255.210 53.075 ;
        RECT 255.210 53.095 255.655 53.125 ;
        POLYGON 255.655 53.130 255.680 53.095 255.655 53.095 ;
        POLYGON 256.305 53.130 256.325 53.130 256.325 53.095 ;
        RECT 256.325 53.095 256.895 53.130 ;
        RECT 255.210 53.075 255.680 53.095 ;
        POLYGON 255.210 53.075 255.235 53.075 255.235 53.045 ;
        RECT 255.235 53.065 255.680 53.075 ;
        POLYGON 255.680 53.095 255.695 53.065 255.680 53.065 ;
        POLYGON 256.325 53.095 256.340 53.095 256.340 53.065 ;
        RECT 256.340 53.065 256.895 53.095 ;
        POLYGON 256.895 53.250 256.980 53.065 256.895 53.065 ;
        POLYGON 257.715 53.250 257.795 53.250 257.795 53.080 ;
        RECT 257.795 53.240 258.665 53.250 ;
        POLYGON 258.665 53.330 258.705 53.240 258.665 53.240 ;
        POLYGON 259.935 53.330 259.955 53.330 259.955 53.280 ;
        RECT 259.955 53.280 261.300 53.330 ;
        POLYGON 259.955 53.280 259.965 53.280 259.965 53.245 ;
        RECT 259.965 53.240 261.300 53.280 ;
        RECT 257.795 53.205 258.705 53.240 ;
        POLYGON 258.705 53.240 258.720 53.205 258.705 53.205 ;
        POLYGON 259.965 53.240 259.975 53.240 259.975 53.210 ;
        RECT 259.975 53.225 261.300 53.240 ;
        POLYGON 261.300 53.615 261.425 53.225 261.300 53.225 ;
        POLYGON 263.360 53.615 263.385 53.615 263.385 53.555 ;
        RECT 263.385 53.595 266.075 53.615 ;
        POLYGON 266.075 53.660 266.095 53.595 266.075 53.595 ;
        POLYGON 270.365 53.660 270.375 53.660 270.375 53.640 ;
        RECT 270.375 53.640 277.205 53.660 ;
        POLYGON 270.375 53.640 270.385 53.640 270.385 53.595 ;
        RECT 270.385 53.595 277.205 53.640 ;
        RECT 263.385 53.555 266.095 53.595 ;
        POLYGON 263.385 53.555 263.480 53.555 263.480 53.225 ;
        RECT 263.480 53.225 266.095 53.555 ;
        RECT 259.975 53.205 261.425 53.225 ;
        RECT 257.795 53.080 258.720 53.205 ;
        POLYGON 257.795 53.080 257.800 53.080 257.800 53.070 ;
        RECT 257.800 53.065 258.720 53.080 ;
        RECT 255.235 53.045 255.695 53.065 ;
        POLYGON 255.235 53.045 255.245 53.045 255.245 53.030 ;
        RECT 255.245 53.030 255.695 53.045 ;
        RECT 253.895 53.025 254.705 53.030 ;
        RECT 244.680 53.005 245.565 53.025 ;
        RECT 243.560 53.000 244.100 53.005 ;
        POLYGON 244.100 53.005 244.105 53.005 244.100 53.000 ;
        RECT 243.560 52.990 244.070 53.000 ;
        RECT 242.050 52.965 242.850 52.990 ;
        POLYGON 242.850 52.990 242.860 52.990 242.850 52.965 ;
        POLYGON 243.535 52.985 243.535 52.965 243.525 52.965 ;
        RECT 243.535 52.965 244.070 52.990 ;
        RECT 242.050 52.895 242.805 52.965 ;
        RECT 239.855 52.875 240.915 52.890 ;
        RECT 236.145 52.840 238.180 52.870 ;
        RECT 229.230 52.725 233.270 52.840 ;
        RECT 229.205 52.590 233.270 52.725 ;
        POLYGON 233.270 52.840 233.290 52.840 233.270 52.605 ;
        POLYGON 236.130 52.835 236.130 52.605 236.100 52.605 ;
        RECT 236.130 52.830 238.180 52.840 ;
        POLYGON 238.180 52.870 238.190 52.870 238.180 52.830 ;
        POLYGON 239.830 52.870 239.830 52.830 239.820 52.830 ;
        RECT 239.830 52.830 240.915 52.875 ;
        RECT 236.130 52.605 238.135 52.830 ;
        RECT 236.100 52.590 238.135 52.605 ;
        POLYGON 238.135 52.830 238.180 52.830 238.135 52.590 ;
        RECT 239.820 52.825 240.915 52.830 ;
        POLYGON 240.915 52.890 240.930 52.890 240.915 52.825 ;
        POLYGON 241.995 52.890 241.995 52.880 241.990 52.880 ;
        RECT 241.995 52.880 242.805 52.895 ;
        POLYGON 241.990 52.880 241.990 52.825 241.970 52.825 ;
        RECT 241.990 52.845 242.805 52.880 ;
        POLYGON 242.805 52.965 242.850 52.965 242.805 52.845 ;
        POLYGON 243.525 52.965 243.525 52.885 243.490 52.885 ;
        RECT 243.525 52.935 244.070 52.965 ;
        POLYGON 244.070 53.000 244.100 53.000 244.070 52.935 ;
        POLYGON 244.660 53.000 244.660 52.940 244.630 52.940 ;
        RECT 244.660 52.940 245.565 53.005 ;
        POLYGON 245.565 53.025 245.620 53.025 245.565 52.940 ;
        POLYGON 253.895 53.025 253.935 53.025 253.935 52.980 ;
        RECT 253.935 52.995 254.705 53.025 ;
        POLYGON 254.705 53.030 254.725 52.995 254.705 52.995 ;
        POLYGON 255.245 53.030 255.255 53.030 255.255 53.015 ;
        RECT 255.255 53.015 255.695 53.030 ;
        POLYGON 255.255 53.015 255.265 53.015 255.265 52.995 ;
        RECT 255.265 52.995 255.695 53.015 ;
        RECT 253.935 52.990 254.725 52.995 ;
        POLYGON 254.725 52.995 254.730 52.990 254.725 52.990 ;
        POLYGON 255.265 52.995 255.270 52.995 255.270 52.990 ;
        RECT 255.270 52.990 255.695 52.995 ;
        RECT 253.935 52.980 254.730 52.990 ;
        POLYGON 253.935 52.980 253.965 52.980 253.965 52.945 ;
        RECT 253.965 52.940 254.730 52.980 ;
        RECT 243.525 52.890 244.045 52.935 ;
        POLYGON 244.045 52.935 244.065 52.935 244.045 52.890 ;
        POLYGON 244.630 52.935 244.630 52.905 244.615 52.905 ;
        RECT 244.630 52.920 245.550 52.940 ;
        POLYGON 245.550 52.940 245.565 52.940 245.550 52.920 ;
        POLYGON 253.965 52.940 253.985 52.940 253.985 52.920 ;
        RECT 253.985 52.920 254.730 52.940 ;
        RECT 244.630 52.905 245.520 52.920 ;
        POLYGON 244.615 52.905 244.615 52.890 244.605 52.890 ;
        RECT 244.615 52.890 245.520 52.905 ;
        RECT 243.525 52.885 244.040 52.890 ;
        POLYGON 243.490 52.885 243.490 52.850 243.475 52.850 ;
        RECT 243.490 52.875 244.040 52.885 ;
        POLYGON 244.040 52.890 244.045 52.890 244.040 52.875 ;
        POLYGON 244.605 52.890 244.605 52.880 244.600 52.880 ;
        RECT 244.605 52.880 245.520 52.890 ;
        RECT 244.600 52.875 245.520 52.880 ;
        POLYGON 245.520 52.920 245.550 52.920 245.520 52.875 ;
        POLYGON 253.985 52.920 254.000 52.920 254.000 52.905 ;
        RECT 254.000 52.905 254.730 52.920 ;
        POLYGON 254.000 52.905 254.020 52.905 254.020 52.880 ;
        RECT 254.020 52.880 254.730 52.905 ;
        POLYGON 254.730 52.990 254.805 52.880 254.730 52.880 ;
        POLYGON 255.270 52.990 255.300 52.990 255.300 52.945 ;
        RECT 255.300 52.945 255.695 52.990 ;
        POLYGON 255.300 52.945 255.325 52.945 255.325 52.910 ;
        RECT 255.325 52.940 255.695 52.945 ;
        POLYGON 255.695 53.065 255.765 52.940 255.695 52.940 ;
        POLYGON 256.340 53.065 256.355 53.065 256.355 53.035 ;
        RECT 256.355 53.035 256.980 53.065 ;
        POLYGON 256.355 53.035 256.365 53.035 256.365 53.010 ;
        RECT 256.365 53.030 256.980 53.035 ;
        POLYGON 256.980 53.065 256.995 53.030 256.980 53.030 ;
        POLYGON 257.800 53.065 257.805 53.065 257.805 53.060 ;
        RECT 257.805 53.060 258.720 53.065 ;
        POLYGON 257.805 53.060 257.815 53.060 257.815 53.030 ;
        RECT 257.815 53.030 258.720 53.060 ;
        RECT 256.365 53.010 256.995 53.030 ;
        POLYGON 256.995 53.030 257.005 53.010 256.995 53.010 ;
        POLYGON 257.815 53.030 257.820 53.030 257.820 53.020 ;
        RECT 257.820 53.010 258.720 53.030 ;
        POLYGON 256.365 53.010 256.400 53.010 256.400 52.940 ;
        RECT 256.400 52.940 257.005 53.010 ;
        RECT 255.325 52.910 255.765 52.940 ;
        POLYGON 255.325 52.910 255.340 52.910 255.340 52.880 ;
        RECT 255.340 52.880 255.765 52.910 ;
        RECT 254.020 52.875 254.805 52.880 ;
        RECT 243.490 52.850 244.000 52.875 ;
        RECT 241.990 52.825 242.780 52.845 ;
        POLYGON 239.820 52.825 239.820 52.590 239.770 52.590 ;
        RECT 239.820 52.625 240.870 52.825 ;
        POLYGON 240.870 52.825 240.915 52.825 240.870 52.625 ;
        POLYGON 241.970 52.820 241.970 52.625 241.905 52.625 ;
        RECT 241.970 52.780 242.780 52.825 ;
        POLYGON 242.780 52.845 242.805 52.845 242.780 52.780 ;
        POLYGON 243.475 52.845 243.475 52.810 243.460 52.810 ;
        RECT 243.475 52.810 244.000 52.850 ;
        POLYGON 243.460 52.810 243.460 52.785 243.450 52.785 ;
        RECT 243.460 52.790 244.000 52.810 ;
        POLYGON 244.000 52.875 244.040 52.875 244.000 52.790 ;
        POLYGON 244.600 52.875 244.600 52.790 244.565 52.790 ;
        RECT 244.600 52.840 245.500 52.875 ;
        POLYGON 245.500 52.875 245.520 52.875 245.500 52.840 ;
        POLYGON 254.020 52.875 254.050 52.875 254.050 52.840 ;
        RECT 254.050 52.860 254.805 52.875 ;
        POLYGON 254.805 52.880 254.815 52.860 254.805 52.860 ;
        POLYGON 255.340 52.880 255.345 52.880 255.345 52.875 ;
        RECT 255.345 52.875 255.765 52.880 ;
        POLYGON 255.765 52.940 255.805 52.875 255.765 52.875 ;
        POLYGON 256.400 52.940 256.405 52.940 256.405 52.935 ;
        RECT 256.405 52.935 257.005 52.940 ;
        POLYGON 256.405 52.935 256.425 52.935 256.425 52.885 ;
        RECT 256.425 52.895 257.005 52.935 ;
        POLYGON 257.005 53.010 257.060 52.895 257.005 52.895 ;
        POLYGON 257.820 53.010 257.870 53.010 257.870 52.900 ;
        RECT 257.870 52.945 258.720 53.010 ;
        POLYGON 258.720 53.205 258.820 52.945 258.720 52.945 ;
        POLYGON 259.975 53.205 260.055 53.205 260.055 52.950 ;
        RECT 260.055 53.000 261.425 53.205 ;
        POLYGON 261.425 53.225 261.485 53.000 261.425 53.000 ;
        POLYGON 263.480 53.225 263.495 53.225 263.495 53.175 ;
        RECT 263.495 53.175 266.095 53.225 ;
        POLYGON 263.495 53.175 263.535 53.175 263.535 53.050 ;
        RECT 263.535 53.080 266.095 53.175 ;
        POLYGON 266.095 53.595 266.230 53.080 266.095 53.080 ;
        POLYGON 270.385 53.595 270.445 53.595 270.445 53.335 ;
        RECT 270.445 53.335 277.205 53.595 ;
        POLYGON 270.445 53.335 270.485 53.335 270.485 53.095 ;
        RECT 270.485 53.320 277.205 53.335 ;
        POLYGON 277.205 53.680 277.290 53.320 277.205 53.320 ;
        RECT 270.485 53.080 277.290 53.320 ;
        RECT 263.535 53.050 266.230 53.080 ;
        POLYGON 263.535 53.050 263.545 53.050 263.545 53.010 ;
        RECT 263.545 53.015 266.230 53.050 ;
        POLYGON 266.230 53.080 266.245 53.015 266.230 53.015 ;
        POLYGON 270.485 53.080 270.495 53.080 270.495 53.035 ;
        RECT 270.495 53.015 277.290 53.080 ;
        RECT 263.545 53.000 266.245 53.015 ;
        RECT 260.055 52.975 261.485 53.000 ;
        POLYGON 261.485 53.000 261.495 52.975 261.485 52.975 ;
        POLYGON 263.545 53.000 263.550 53.000 263.550 52.990 ;
        RECT 263.550 52.975 266.245 53.000 ;
        RECT 260.055 52.945 261.495 52.975 ;
        RECT 257.870 52.910 258.820 52.945 ;
        POLYGON 258.820 52.945 258.830 52.910 258.820 52.910 ;
        POLYGON 260.055 52.945 260.065 52.945 260.065 52.915 ;
        RECT 260.065 52.910 261.495 52.945 ;
        RECT 257.870 52.895 258.830 52.910 ;
        RECT 256.425 52.885 257.060 52.895 ;
        POLYGON 256.425 52.885 256.430 52.885 256.430 52.875 ;
        RECT 256.430 52.875 257.060 52.885 ;
        POLYGON 255.345 52.875 255.350 52.875 255.350 52.865 ;
        RECT 255.350 52.860 255.805 52.875 ;
        RECT 254.050 52.840 254.815 52.860 ;
        RECT 244.600 52.790 245.465 52.840 ;
        RECT 243.460 52.785 243.995 52.790 ;
        POLYGON 243.995 52.790 244.000 52.790 243.995 52.785 ;
        RECT 244.565 52.785 245.465 52.790 ;
        POLYGON 245.465 52.840 245.500 52.840 245.465 52.785 ;
        POLYGON 254.050 52.840 254.065 52.840 254.065 52.825 ;
        RECT 254.065 52.825 254.815 52.840 ;
        POLYGON 254.065 52.825 254.075 52.825 254.075 52.810 ;
        RECT 254.075 52.810 254.815 52.825 ;
        POLYGON 254.075 52.810 254.090 52.810 254.090 52.790 ;
        RECT 254.090 52.785 254.815 52.810 ;
        RECT 241.970 52.625 242.720 52.780 ;
        RECT 239.820 52.590 240.865 52.625 ;
        POLYGON 240.865 52.625 240.870 52.625 240.865 52.600 ;
        POLYGON 241.905 52.625 241.905 52.600 241.895 52.600 ;
        RECT 241.905 52.600 242.720 52.625 ;
        RECT 182.485 52.390 196.860 52.590 ;
        RECT 171.405 52.225 175.575 52.390 ;
        POLYGON 168.755 52.225 168.795 52.035 168.755 52.035 ;
        POLYGON 171.405 52.225 171.435 52.225 171.435 52.070 ;
        RECT 171.435 52.070 175.575 52.225 ;
        POLYGON 171.435 52.070 171.440 52.070 171.440 52.045 ;
        RECT 171.440 52.035 175.575 52.070 ;
        RECT 166.720 52.005 168.795 52.035 ;
        POLYGON 166.720 52.005 166.730 52.005 166.730 51.940 ;
        RECT 166.730 51.935 168.795 52.005 ;
        RECT 164.140 51.860 165.290 51.935 ;
        RECT 162.440 51.785 163.245 51.860 ;
        RECT 161.280 51.770 161.805 51.785 ;
        RECT 160.350 51.740 160.795 51.770 ;
        RECT 149.995 51.705 159.705 51.740 ;
        POLYGON 149.920 51.705 149.920 51.660 149.905 51.660 ;
        RECT 149.920 51.690 159.705 51.705 ;
        POLYGON 159.705 51.740 159.720 51.690 159.705 51.690 ;
        POLYGON 160.350 51.740 160.370 51.740 160.370 51.695 ;
        RECT 160.370 51.690 160.795 51.740 ;
        RECT 149.920 51.660 159.720 51.690 ;
        RECT 148.620 51.630 149.155 51.660 ;
        RECT 117.205 51.455 148.050 51.625 ;
        RECT 53.295 50.930 111.645 51.455 ;
        POLYGON 111.645 51.455 111.745 50.930 111.645 50.930 ;
        RECT 117.195 51.450 148.050 51.455 ;
        POLYGON 148.050 51.625 148.085 51.625 148.050 51.450 ;
        POLYGON 148.605 51.625 148.605 51.595 148.595 51.595 ;
        RECT 148.605 51.595 149.155 51.630 ;
        POLYGON 148.595 51.595 148.595 51.565 148.590 51.565 ;
        RECT 148.595 51.565 149.155 51.595 ;
        POLYGON 148.590 51.565 148.590 51.450 148.560 51.450 ;
        RECT 148.590 51.500 149.155 51.565 ;
        POLYGON 149.155 51.660 149.185 51.660 149.155 51.500 ;
        POLYGON 149.905 51.660 149.905 51.520 149.860 51.520 ;
        RECT 149.905 51.650 159.720 51.660 ;
        POLYGON 159.720 51.690 159.735 51.650 159.720 51.650 ;
        POLYGON 160.370 51.690 160.380 51.690 160.380 51.670 ;
        RECT 160.380 51.670 160.795 51.690 ;
        POLYGON 160.380 51.670 160.385 51.670 160.385 51.655 ;
        RECT 160.385 51.660 160.795 51.670 ;
        POLYGON 160.795 51.770 160.820 51.660 160.795 51.660 ;
        RECT 160.385 51.650 160.820 51.660 ;
        POLYGON 161.280 51.770 161.315 51.770 161.315 51.650 ;
        RECT 161.315 51.650 161.805 51.770 ;
        RECT 149.905 51.590 159.735 51.650 ;
        POLYGON 159.735 51.650 159.760 51.590 159.735 51.590 ;
        POLYGON 160.385 51.650 160.405 51.650 160.405 51.590 ;
        RECT 160.405 51.590 160.820 51.650 ;
        RECT 149.905 51.520 159.760 51.590 ;
        POLYGON 149.860 51.520 149.860 51.510 149.855 51.510 ;
        RECT 149.860 51.510 159.760 51.520 ;
        POLYGON 159.760 51.590 159.785 51.510 159.760 51.510 ;
        POLYGON 160.405 51.590 160.430 51.590 160.430 51.510 ;
        RECT 160.430 51.510 160.820 51.590 ;
        RECT 148.590 51.450 149.140 51.500 ;
        RECT 117.195 51.395 148.040 51.450 ;
        POLYGON 148.040 51.450 148.050 51.450 148.040 51.395 ;
        POLYGON 148.560 51.440 148.560 51.400 148.550 51.400 ;
        RECT 148.560 51.435 149.140 51.450 ;
        POLYGON 149.140 51.500 149.155 51.500 149.140 51.435 ;
        POLYGON 149.855 51.500 149.855 51.435 149.835 51.435 ;
        RECT 149.855 51.475 159.785 51.510 ;
        POLYGON 159.785 51.510 159.795 51.475 159.785 51.475 ;
        POLYGON 160.430 51.510 160.440 51.510 160.440 51.480 ;
        RECT 160.440 51.475 160.820 51.510 ;
        RECT 149.855 51.435 159.795 51.475 ;
        POLYGON 159.795 51.475 159.810 51.435 159.795 51.435 ;
        POLYGON 160.440 51.475 160.450 51.475 160.450 51.450 ;
        RECT 160.450 51.450 160.820 51.475 ;
        POLYGON 160.820 51.650 160.860 51.450 160.820 51.450 ;
        POLYGON 161.315 51.650 161.325 51.650 161.325 51.620 ;
        RECT 161.325 51.620 161.805 51.650 ;
        POLYGON 161.805 51.785 161.850 51.620 161.805 51.620 ;
        POLYGON 162.440 51.785 162.465 51.785 162.465 51.695 ;
        RECT 162.465 51.765 163.245 51.785 ;
        POLYGON 163.245 51.860 163.270 51.765 163.245 51.765 ;
        POLYGON 164.140 51.860 164.155 51.860 164.155 51.805 ;
        RECT 164.155 51.795 165.290 51.860 ;
        POLYGON 164.155 51.795 164.160 51.795 164.160 51.770 ;
        RECT 164.160 51.765 165.290 51.795 ;
        RECT 162.465 51.695 163.270 51.765 ;
        POLYGON 162.465 51.695 162.480 51.695 162.480 51.630 ;
        RECT 162.480 51.620 163.270 51.695 ;
        POLYGON 161.325 51.620 161.360 51.620 161.360 51.505 ;
        RECT 161.360 51.505 161.850 51.620 ;
        POLYGON 161.360 51.505 161.370 51.505 161.370 51.465 ;
        RECT 161.370 51.480 161.850 51.505 ;
        POLYGON 161.850 51.620 161.885 51.480 161.850 51.480 ;
        POLYGON 162.480 51.620 162.515 51.620 162.515 51.490 ;
        RECT 162.515 51.480 163.270 51.620 ;
        RECT 161.370 51.450 161.885 51.480 ;
        RECT 148.560 51.420 149.135 51.435 ;
        POLYGON 149.135 51.435 149.140 51.435 149.135 51.420 ;
        POLYGON 149.835 51.435 149.835 51.420 149.830 51.420 ;
        RECT 149.835 51.420 159.810 51.435 ;
        POLYGON 160.450 51.450 160.455 51.450 160.455 51.430 ;
        RECT 160.455 51.430 160.860 51.450 ;
        RECT 148.560 51.400 149.090 51.420 ;
        RECT 117.195 51.335 148.030 51.395 ;
        POLYGON 148.030 51.395 148.040 51.395 148.030 51.335 ;
        POLYGON 148.550 51.395 148.550 51.335 148.540 51.335 ;
        RECT 148.550 51.335 149.090 51.400 ;
        POLYGON 117.195 51.330 117.195 50.930 117.185 50.930 ;
        RECT 117.195 51.220 148.010 51.335 ;
        POLYGON 148.010 51.335 148.030 51.335 148.010 51.220 ;
        POLYGON 148.540 51.330 148.540 51.230 148.520 51.230 ;
        RECT 148.540 51.230 149.090 51.335 ;
        RECT 117.195 51.155 148.005 51.220 ;
        POLYGON 148.005 51.220 148.010 51.220 148.005 51.155 ;
        POLYGON 148.520 51.220 148.520 51.205 148.515 51.205 ;
        RECT 148.520 51.205 149.090 51.230 ;
        POLYGON 148.515 51.205 148.515 51.170 148.510 51.170 ;
        RECT 148.515 51.170 149.090 51.205 ;
        RECT 117.195 51.115 148.000 51.155 ;
        POLYGON 148.000 51.155 148.005 51.155 148.000 51.125 ;
        POLYGON 148.000 51.125 148.005 51.115 148.000 51.115 ;
        POLYGON 148.510 51.155 148.510 51.125 148.505 51.125 ;
        RECT 148.510 51.125 149.090 51.170 ;
        RECT 117.195 51.015 148.005 51.115 ;
        POLYGON 148.005 51.115 148.040 51.015 148.005 51.015 ;
        RECT 117.195 50.985 148.040 51.015 ;
        POLYGON 148.505 51.115 148.505 51.005 148.485 51.005 ;
        RECT 148.505 51.110 149.090 51.125 ;
        POLYGON 149.090 51.420 149.135 51.420 149.090 51.120 ;
        POLYGON 149.830 51.415 149.830 51.315 149.800 51.315 ;
        RECT 149.830 51.365 159.810 51.420 ;
        POLYGON 159.810 51.430 159.830 51.365 159.810 51.365 ;
        POLYGON 160.455 51.430 160.470 51.430 160.470 51.370 ;
        RECT 160.470 51.365 160.860 51.430 ;
        RECT 149.830 51.315 159.830 51.365 ;
        POLYGON 149.800 51.315 149.800 51.300 149.795 51.300 ;
        RECT 149.800 51.300 159.830 51.315 ;
        POLYGON 149.795 51.300 149.795 51.120 149.755 51.120 ;
        RECT 149.795 51.205 159.830 51.300 ;
        POLYGON 159.830 51.365 159.870 51.205 159.830 51.205 ;
        POLYGON 160.470 51.365 160.475 51.365 160.475 51.355 ;
        RECT 160.475 51.355 160.860 51.365 ;
        POLYGON 160.475 51.355 160.510 51.355 160.510 51.230 ;
        RECT 160.510 51.335 160.860 51.355 ;
        POLYGON 160.860 51.450 160.875 51.335 160.860 51.335 ;
        POLYGON 161.370 51.450 161.400 51.450 161.400 51.345 ;
        RECT 161.400 51.335 161.885 51.450 ;
        POLYGON 161.885 51.480 161.920 51.335 161.885 51.335 ;
        POLYGON 162.515 51.480 162.540 51.480 162.540 51.390 ;
        RECT 162.540 51.435 163.270 51.480 ;
        POLYGON 163.270 51.765 163.350 51.435 163.270 51.435 ;
        POLYGON 164.160 51.765 164.225 51.765 164.225 51.445 ;
        RECT 164.225 51.760 165.290 51.765 ;
        POLYGON 165.290 51.935 165.325 51.760 165.290 51.760 ;
        POLYGON 166.730 51.935 166.760 51.935 166.760 51.760 ;
        RECT 166.760 51.810 168.795 51.935 ;
        POLYGON 168.795 52.035 168.840 51.810 168.795 51.810 ;
        POLYGON 171.440 52.035 171.485 52.035 171.485 51.825 ;
        RECT 171.485 51.810 175.575 52.035 ;
        RECT 166.760 51.770 168.840 51.810 ;
        POLYGON 168.840 51.810 168.850 51.770 168.840 51.770 ;
        POLYGON 171.485 51.810 171.490 51.810 171.490 51.805 ;
        RECT 171.490 51.805 175.575 51.810 ;
        POLYGON 171.490 51.805 171.495 51.805 171.495 51.770 ;
        RECT 171.495 51.770 175.575 51.805 ;
        RECT 166.760 51.760 168.850 51.770 ;
        RECT 164.225 51.435 165.325 51.760 ;
        RECT 162.540 51.390 163.350 51.435 ;
        POLYGON 162.540 51.390 162.550 51.390 162.550 51.335 ;
        RECT 162.550 51.335 163.350 51.390 ;
        POLYGON 163.350 51.435 163.370 51.335 163.350 51.335 ;
        POLYGON 164.225 51.435 164.240 51.435 164.240 51.375 ;
        RECT 164.240 51.375 165.325 51.435 ;
        POLYGON 164.240 51.375 164.245 51.375 164.245 51.340 ;
        RECT 164.245 51.335 165.325 51.375 ;
        RECT 160.510 51.230 160.875 51.335 ;
        POLYGON 160.510 51.230 160.515 51.230 160.515 51.205 ;
        RECT 160.515 51.205 160.875 51.230 ;
        RECT 149.795 51.140 159.870 51.205 ;
        POLYGON 159.870 51.205 159.880 51.140 159.870 51.140 ;
        POLYGON 160.515 51.205 160.525 51.205 160.525 51.165 ;
        RECT 160.525 51.165 160.875 51.205 ;
        POLYGON 160.525 51.165 160.530 51.165 160.530 51.140 ;
        RECT 160.530 51.140 160.875 51.165 ;
        RECT 149.795 51.120 159.880 51.140 ;
        RECT 148.505 51.030 149.080 51.110 ;
        POLYGON 149.080 51.110 149.090 51.110 149.080 51.030 ;
        POLYGON 149.755 51.120 149.755 51.035 149.740 51.035 ;
        RECT 149.755 51.065 159.880 51.120 ;
        POLYGON 159.880 51.140 159.895 51.065 159.880 51.065 ;
        POLYGON 160.530 51.140 160.545 51.140 160.545 51.075 ;
        RECT 160.545 51.115 160.875 51.140 ;
        POLYGON 160.875 51.335 160.910 51.115 160.875 51.115 ;
        POLYGON 161.400 51.335 161.430 51.335 161.430 51.225 ;
        RECT 161.430 51.310 161.920 51.335 ;
        POLYGON 161.920 51.335 161.925 51.310 161.920 51.310 ;
        RECT 162.550 51.310 163.370 51.335 ;
        RECT 161.430 51.225 161.925 51.310 ;
        POLYGON 161.430 51.225 161.455 51.225 161.455 51.115 ;
        RECT 161.455 51.165 161.925 51.225 ;
        POLYGON 161.925 51.310 161.960 51.165 161.925 51.165 ;
        POLYGON 162.550 51.310 162.580 51.310 162.580 51.170 ;
        RECT 162.580 51.205 163.370 51.310 ;
        POLYGON 163.370 51.335 163.395 51.205 163.370 51.205 ;
        POLYGON 164.245 51.335 164.260 51.335 164.260 51.240 ;
        RECT 164.260 51.330 165.325 51.335 ;
        POLYGON 165.325 51.760 165.385 51.330 165.325 51.330 ;
        POLYGON 166.760 51.760 166.790 51.760 166.790 51.580 ;
        RECT 166.790 51.580 168.850 51.760 ;
        POLYGON 166.790 51.580 166.825 51.580 166.825 51.350 ;
        RECT 166.825 51.535 168.850 51.580 ;
        POLYGON 168.850 51.770 168.890 51.535 168.850 51.535 ;
        POLYGON 171.495 51.770 171.530 51.770 171.530 51.540 ;
        RECT 171.530 51.535 175.575 51.770 ;
        RECT 166.825 51.330 168.890 51.535 ;
        RECT 164.260 51.240 165.385 51.330 ;
        POLYGON 164.260 51.240 164.265 51.240 164.265 51.205 ;
        RECT 164.265 51.210 165.385 51.240 ;
        POLYGON 165.385 51.330 165.400 51.210 165.385 51.210 ;
        POLYGON 166.825 51.330 166.840 51.330 166.840 51.230 ;
        RECT 166.840 51.290 168.890 51.330 ;
        POLYGON 168.890 51.535 168.930 51.290 168.890 51.290 ;
        POLYGON 171.530 51.535 171.565 51.535 171.565 51.310 ;
        RECT 171.565 51.290 175.575 51.535 ;
        RECT 166.840 51.210 168.930 51.290 ;
        RECT 164.265 51.205 165.400 51.210 ;
        RECT 162.580 51.165 163.395 51.205 ;
        RECT 161.455 51.115 161.960 51.165 ;
        RECT 160.545 51.065 160.910 51.115 ;
        RECT 149.755 51.035 159.895 51.065 ;
        RECT 148.505 51.005 149.055 51.030 ;
        POLYGON 148.040 51.005 148.050 50.985 148.040 50.985 ;
        POLYGON 148.485 51.005 148.485 50.985 148.480 50.985 ;
        RECT 148.485 50.985 149.055 51.005 ;
        RECT 117.195 50.970 148.050 50.985 ;
        POLYGON 148.050 50.985 148.055 50.970 148.050 50.970 ;
        RECT 117.195 50.930 148.055 50.970 ;
        POLYGON 148.055 50.965 148.070 50.930 148.055 50.930 ;
        RECT 53.295 50.000 111.745 50.930 ;
        POLYGON 13.270 50.000 13.355 50.000 13.355 44.770 ;
        RECT 13.355 44.770 22.040 50.000 ;
        POLYGON 13.355 44.770 13.610 44.770 13.610 39.610 ;
        RECT 13.610 42.000 22.040 44.770 ;
        POLYGON 22.040 50.000 22.195 42.000 22.040 42.000 ;
        POLYGON 53.295 50.000 53.325 50.000 53.325 49.915 ;
        RECT 53.325 49.915 111.745 50.000 ;
        POLYGON 53.325 49.915 53.440 49.915 53.440 49.575 ;
        RECT 53.440 49.575 111.745 49.915 ;
        POLYGON 53.440 49.575 54.910 49.575 54.910 45.915 ;
        RECT 54.910 49.500 111.745 49.575 ;
        POLYGON 111.745 50.930 112.015 49.500 111.745 49.500 ;
        RECT 117.185 50.815 148.070 50.930 ;
        POLYGON 148.480 50.965 148.480 50.925 148.475 50.925 ;
        RECT 148.480 50.925 149.055 50.985 ;
        POLYGON 148.070 50.925 148.110 50.815 148.070 50.815 ;
        POLYGON 117.185 50.800 117.185 50.535 117.180 50.535 ;
        RECT 117.185 50.760 148.110 50.815 ;
        POLYGON 148.475 50.925 148.475 50.810 148.460 50.810 ;
        RECT 148.475 50.810 149.055 50.925 ;
        POLYGON 148.110 50.810 148.130 50.760 148.110 50.760 ;
        RECT 117.185 50.690 148.130 50.760 ;
        POLYGON 148.460 50.810 148.460 50.765 148.455 50.765 ;
        RECT 148.460 50.795 149.055 50.810 ;
        POLYGON 149.055 51.030 149.080 51.030 149.055 50.795 ;
        POLYGON 149.740 51.030 149.740 50.925 149.720 50.925 ;
        RECT 149.740 51.015 159.895 51.035 ;
        POLYGON 159.895 51.065 159.900 51.015 159.895 51.015 ;
        POLYGON 160.545 51.065 160.555 51.065 160.555 51.030 ;
        RECT 160.555 51.015 160.910 51.065 ;
        RECT 149.740 50.925 159.900 51.015 ;
        POLYGON 149.720 50.925 149.720 50.815 149.705 50.815 ;
        RECT 149.720 50.845 159.900 50.925 ;
        POLYGON 159.900 51.015 159.930 50.845 159.900 50.845 ;
        POLYGON 160.555 51.015 160.560 51.015 160.560 51.010 ;
        RECT 160.560 51.010 160.910 51.015 ;
        POLYGON 160.560 51.010 160.580 51.010 160.580 50.915 ;
        RECT 160.580 50.980 160.910 51.010 ;
        POLYGON 160.910 51.115 160.925 50.980 160.910 50.980 ;
        POLYGON 161.455 51.115 161.480 51.115 161.480 50.995 ;
        RECT 161.480 51.025 161.960 51.115 ;
        POLYGON 161.960 51.165 161.985 51.025 161.960 51.025 ;
        POLYGON 162.580 51.165 162.585 51.165 162.585 51.145 ;
        RECT 162.585 51.145 163.395 51.165 ;
        POLYGON 162.585 51.145 162.600 51.145 162.600 51.080 ;
        RECT 162.600 51.085 163.395 51.145 ;
        POLYGON 163.395 51.205 163.420 51.085 163.395 51.085 ;
        POLYGON 164.265 51.205 164.280 51.205 164.280 51.105 ;
        RECT 164.280 51.085 165.400 51.205 ;
        RECT 162.600 51.080 163.420 51.085 ;
        POLYGON 162.600 51.080 162.605 51.080 162.605 51.040 ;
        RECT 162.605 51.025 163.420 51.080 ;
        RECT 161.480 50.980 161.985 51.025 ;
        RECT 160.580 50.915 160.925 50.980 ;
        POLYGON 160.580 50.915 160.590 50.915 160.590 50.865 ;
        RECT 160.590 50.845 160.925 50.915 ;
        RECT 149.720 50.815 159.930 50.845 ;
        POLYGON 149.705 50.815 149.705 50.795 149.700 50.795 ;
        RECT 149.705 50.795 159.930 50.815 ;
        RECT 148.460 50.765 149.030 50.795 ;
        POLYGON 148.130 50.755 148.155 50.690 148.130 50.690 ;
        RECT 117.185 50.675 148.155 50.690 ;
        POLYGON 148.455 50.755 148.455 50.685 148.445 50.685 ;
        RECT 148.455 50.685 149.030 50.765 ;
        POLYGON 148.155 50.685 148.160 50.675 148.155 50.675 ;
        RECT 117.185 50.620 148.160 50.675 ;
        POLYGON 148.160 50.670 148.180 50.620 148.160 50.620 ;
        RECT 117.185 50.535 148.180 50.620 ;
        POLYGON 148.445 50.670 148.445 50.610 148.440 50.610 ;
        RECT 148.445 50.610 149.030 50.685 ;
        RECT 117.180 50.520 148.180 50.535 ;
        POLYGON 148.180 50.610 148.215 50.520 148.180 50.520 ;
        POLYGON 148.440 50.610 148.440 50.540 148.435 50.540 ;
        RECT 148.440 50.540 149.030 50.610 ;
        POLYGON 117.180 50.495 117.180 50.000 117.170 50.000 ;
        RECT 117.180 50.450 148.215 50.520 ;
        POLYGON 148.215 50.520 148.240 50.450 148.215 50.450 ;
        RECT 117.180 50.320 148.240 50.450 ;
        POLYGON 148.435 50.520 148.435 50.475 148.430 50.475 ;
        RECT 148.435 50.475 149.030 50.540 ;
        POLYGON 148.240 50.440 148.285 50.320 148.240 50.320 ;
        RECT 117.180 50.020 148.285 50.320 ;
        POLYGON 148.430 50.440 148.430 50.405 148.425 50.405 ;
        RECT 148.430 50.425 149.030 50.475 ;
        POLYGON 149.030 50.795 149.055 50.795 149.030 50.465 ;
        POLYGON 149.700 50.785 149.700 50.725 149.690 50.725 ;
        RECT 149.700 50.780 159.930 50.795 ;
        POLYGON 159.930 50.845 159.940 50.780 159.930 50.780 ;
        POLYGON 160.590 50.845 160.605 50.845 160.605 50.790 ;
        RECT 160.605 50.780 160.925 50.845 ;
        RECT 149.700 50.725 159.940 50.780 ;
        POLYGON 149.690 50.725 149.690 50.530 149.675 50.530 ;
        RECT 149.690 50.655 159.940 50.725 ;
        POLYGON 159.940 50.780 159.955 50.655 159.940 50.655 ;
        POLYGON 160.605 50.780 160.610 50.780 160.610 50.750 ;
        RECT 160.610 50.760 160.925 50.780 ;
        POLYGON 160.925 50.980 160.945 50.760 160.925 50.760 ;
        POLYGON 161.480 50.980 161.490 50.980 161.490 50.950 ;
        RECT 161.490 50.950 161.985 50.980 ;
        POLYGON 161.490 50.950 161.515 50.950 161.515 50.775 ;
        RECT 161.515 50.865 161.985 50.950 ;
        POLYGON 161.985 51.025 162.015 50.865 161.985 50.865 ;
        POLYGON 162.605 51.025 162.630 51.025 162.630 50.865 ;
        RECT 162.630 51.010 163.420 51.025 ;
        POLYGON 163.420 51.085 163.435 51.010 163.420 51.010 ;
        POLYGON 164.280 51.085 164.290 51.085 164.290 51.040 ;
        RECT 164.290 51.010 165.400 51.085 ;
        RECT 162.630 50.910 163.435 51.010 ;
        POLYGON 163.435 51.010 163.450 50.910 163.435 50.910 ;
        POLYGON 164.290 51.010 164.305 51.010 164.305 50.940 ;
        RECT 164.305 50.910 165.400 51.010 ;
        RECT 162.630 50.865 163.450 50.910 ;
        RECT 161.515 50.760 162.015 50.865 ;
        RECT 160.610 50.750 160.945 50.760 ;
        POLYGON 160.610 50.750 160.620 50.750 160.620 50.680 ;
        RECT 160.620 50.655 160.945 50.750 ;
        RECT 149.690 50.530 159.955 50.655 ;
        RECT 149.675 50.480 159.955 50.530 ;
        POLYGON 159.955 50.655 159.975 50.480 159.955 50.480 ;
        POLYGON 160.620 50.655 160.630 50.655 160.630 50.615 ;
        RECT 160.630 50.630 160.945 50.655 ;
        POLYGON 160.945 50.760 160.955 50.630 160.945 50.630 ;
        POLYGON 161.515 50.760 161.530 50.760 161.530 50.670 ;
        RECT 161.530 50.740 162.015 50.760 ;
        POLYGON 162.015 50.865 162.030 50.740 162.015 50.740 ;
        POLYGON 162.630 50.865 162.645 50.865 162.645 50.770 ;
        RECT 162.645 50.740 163.450 50.865 ;
        RECT 161.530 50.670 162.030 50.740 ;
        POLYGON 161.530 50.670 161.535 50.670 161.535 50.630 ;
        RECT 160.630 50.615 160.955 50.630 ;
        POLYGON 160.630 50.615 160.635 50.615 160.635 50.570 ;
        RECT 160.635 50.570 160.955 50.615 ;
        RECT 161.535 50.610 162.030 50.670 ;
        POLYGON 160.635 50.570 160.645 50.570 160.645 50.485 ;
        RECT 160.645 50.480 160.955 50.570 ;
        RECT 148.430 50.405 149.025 50.425 ;
        POLYGON 148.285 50.315 148.390 50.020 148.285 50.020 ;
        RECT 117.180 50.000 148.390 50.020 ;
        POLYGON 148.425 50.315 148.425 50.205 148.420 50.205 ;
        RECT 148.425 50.205 149.025 50.405 ;
        POLYGON 117.170 50.000 117.175 50.000 117.175 49.730 ;
        RECT 117.175 49.935 148.390 50.000 ;
        POLYGON 148.390 50.015 148.420 49.935 148.390 49.935 ;
        RECT 148.420 50.005 149.025 50.205 ;
        POLYGON 149.025 50.425 149.030 50.425 149.025 50.130 ;
        POLYGON 148.420 50.005 148.425 50.005 148.425 49.935 ;
        RECT 117.175 49.925 148.420 49.935 ;
        POLYGON 148.420 49.935 148.425 49.925 148.420 49.925 ;
        RECT 148.425 49.925 149.025 50.005 ;
        RECT 117.175 49.800 149.025 49.925 ;
        POLYGON 149.025 50.130 149.030 49.800 149.025 49.800 ;
        POLYGON 149.675 50.465 149.675 50.335 149.670 50.335 ;
        RECT 149.675 50.435 159.975 50.480 ;
        POLYGON 159.975 50.480 159.980 50.435 159.975 50.435 ;
        POLYGON 160.645 50.480 160.650 50.480 160.650 50.445 ;
        RECT 160.650 50.435 160.955 50.480 ;
        POLYGON 149.670 50.335 149.675 50.335 149.675 50.110 ;
        RECT 149.675 50.285 159.980 50.435 ;
        POLYGON 159.980 50.435 159.985 50.285 159.980 50.285 ;
        POLYGON 160.650 50.435 160.660 50.435 160.660 50.365 ;
        RECT 160.660 50.395 160.955 50.435 ;
        POLYGON 160.955 50.610 160.970 50.395 160.955 50.395 ;
        POLYGON 161.535 50.610 161.560 50.610 161.560 50.430 ;
        RECT 161.560 50.585 162.030 50.610 ;
        POLYGON 162.030 50.740 162.055 50.585 162.030 50.585 ;
        POLYGON 162.645 50.740 162.665 50.740 162.665 50.590 ;
        RECT 161.560 50.440 162.055 50.585 ;
        RECT 162.665 50.585 163.450 50.740 ;
        POLYGON 163.450 50.910 163.495 50.585 163.450 50.585 ;
        POLYGON 164.305 50.910 164.340 50.910 164.340 50.595 ;
        RECT 164.340 50.755 165.400 50.910 ;
        POLYGON 165.400 51.210 165.445 50.755 165.400 50.755 ;
        POLYGON 166.840 51.210 166.850 51.210 166.850 51.150 ;
        RECT 166.850 51.150 168.930 51.210 ;
        POLYGON 166.850 51.150 166.885 51.150 166.885 50.765 ;
        RECT 166.885 51.035 168.930 51.150 ;
        POLYGON 168.930 51.290 168.965 51.035 168.930 51.035 ;
        POLYGON 171.565 51.290 171.600 51.290 171.600 51.080 ;
        RECT 171.600 51.035 175.575 51.290 ;
        RECT 166.885 50.805 168.965 51.035 ;
        POLYGON 168.965 51.035 168.995 50.805 168.965 50.805 ;
        POLYGON 171.600 51.035 171.625 51.035 171.625 50.835 ;
        RECT 171.625 50.970 175.575 51.035 ;
        POLYGON 175.575 52.390 175.670 50.970 175.575 50.970 ;
        POLYGON 182.485 52.390 182.620 52.390 182.620 51.635 ;
        RECT 182.620 51.635 196.860 52.390 ;
        POLYGON 182.620 51.635 182.665 51.635 182.665 51.260 ;
        RECT 182.665 51.515 196.860 51.635 ;
        POLYGON 196.860 52.590 197.095 51.515 196.860 51.515 ;
        POLYGON 206.535 52.590 206.685 52.590 206.685 51.525 ;
        RECT 182.665 51.505 197.095 51.515 ;
        POLYGON 197.095 51.515 197.100 51.505 197.095 51.505 ;
        RECT 206.685 51.505 222.230 52.590 ;
        RECT 182.665 51.260 197.100 51.505 ;
        POLYGON 182.665 51.260 182.700 51.260 182.700 50.970 ;
        RECT 182.700 51.030 197.100 51.260 ;
        POLYGON 197.100 51.505 197.200 51.030 197.100 51.030 ;
        POLYGON 206.685 51.505 206.695 51.505 206.695 51.455 ;
        RECT 206.695 51.455 222.230 51.505 ;
        POLYGON 206.695 51.455 206.775 51.455 206.775 51.035 ;
        RECT 206.775 51.030 222.230 51.455 ;
        RECT 182.700 50.970 197.200 51.030 ;
        RECT 171.625 50.805 175.670 50.970 ;
        RECT 166.885 50.755 168.995 50.805 ;
        RECT 164.340 50.640 165.445 50.755 ;
        POLYGON 165.445 50.755 165.455 50.640 165.445 50.640 ;
        POLYGON 166.885 50.755 166.895 50.755 166.895 50.660 ;
        RECT 166.895 50.640 168.995 50.755 ;
        RECT 164.340 50.585 165.455 50.640 ;
        RECT 162.665 50.570 163.495 50.585 ;
        POLYGON 162.055 50.570 162.065 50.440 162.055 50.440 ;
        POLYGON 162.665 50.570 162.680 50.570 162.680 50.455 ;
        RECT 162.680 50.470 163.495 50.570 ;
        POLYGON 163.495 50.585 163.505 50.470 163.495 50.470 ;
        POLYGON 164.340 50.585 164.350 50.585 164.350 50.500 ;
        RECT 164.350 50.470 165.455 50.585 ;
        RECT 162.680 50.440 163.505 50.470 ;
        RECT 161.560 50.395 162.065 50.440 ;
        RECT 160.660 50.285 160.970 50.395 ;
        RECT 149.675 50.135 159.985 50.285 ;
        POLYGON 159.985 50.285 159.995 50.135 159.985 50.135 ;
        RECT 149.675 50.070 159.995 50.135 ;
        POLYGON 160.660 50.285 160.675 50.285 160.675 50.125 ;
        RECT 160.675 50.190 160.970 50.285 ;
        POLYGON 160.970 50.395 160.975 50.190 160.970 50.190 ;
        POLYGON 161.560 50.395 161.565 50.395 161.565 50.390 ;
        RECT 161.565 50.390 162.065 50.395 ;
        POLYGON 161.565 50.390 161.570 50.390 161.570 50.265 ;
        RECT 161.570 50.270 162.065 50.390 ;
        POLYGON 162.065 50.440 162.085 50.270 162.065 50.270 ;
        POLYGON 162.680 50.440 162.690 50.440 162.690 50.295 ;
        RECT 162.690 50.270 163.505 50.440 ;
        RECT 161.570 50.265 162.085 50.270 ;
        POLYGON 149.675 50.070 149.685 50.070 149.685 49.890 ;
        RECT 149.685 49.890 159.995 50.070 ;
        POLYGON 149.685 49.890 149.690 49.890 149.690 49.825 ;
        RECT 117.175 49.575 149.030 49.800 ;
        RECT 149.690 49.790 159.995 49.890 ;
        POLYGON 149.030 49.790 149.045 49.575 149.030 49.575 ;
        POLYGON 149.690 49.790 149.705 49.790 149.705 49.685 ;
        RECT 149.705 49.765 159.995 49.790 ;
        RECT 149.705 49.675 159.975 49.765 ;
        POLYGON 149.705 49.675 149.715 49.675 149.715 49.600 ;
        RECT 149.715 49.575 159.975 49.675 ;
        RECT 117.175 49.500 149.045 49.575 ;
        RECT 54.910 48.615 112.015 49.500 ;
        POLYGON 112.015 49.500 112.180 48.615 112.015 48.615 ;
        POLYGON 117.175 49.500 117.195 49.500 117.195 48.665 ;
        RECT 117.195 49.480 149.045 49.500 ;
        POLYGON 149.045 49.575 149.055 49.480 149.045 49.480 ;
        POLYGON 149.715 49.575 149.720 49.575 149.720 49.565 ;
        RECT 149.720 49.565 159.975 49.575 ;
        POLYGON 149.720 49.565 149.725 49.565 149.725 49.510 ;
        RECT 149.725 49.480 159.975 49.565 ;
        RECT 117.195 49.250 149.055 49.480 ;
        POLYGON 149.055 49.480 149.080 49.250 149.055 49.250 ;
        POLYGON 149.725 49.480 149.730 49.480 149.730 49.460 ;
        RECT 149.730 49.460 159.975 49.480 ;
        POLYGON 149.730 49.460 149.765 49.460 149.765 49.250 ;
        RECT 149.765 49.445 159.975 49.460 ;
        POLYGON 159.975 49.765 159.995 49.765 159.975 49.445 ;
        RECT 160.675 50.085 160.975 50.190 ;
        POLYGON 161.570 50.265 161.580 50.265 161.580 50.110 ;
        RECT 161.580 50.130 162.085 50.265 ;
        POLYGON 162.085 50.270 162.090 50.130 162.085 50.130 ;
        POLYGON 162.690 50.270 162.700 50.270 162.700 50.140 ;
        RECT 162.700 50.155 163.505 50.270 ;
        POLYGON 163.505 50.470 163.535 50.155 163.505 50.155 ;
        POLYGON 164.350 50.470 164.365 50.470 164.365 50.235 ;
        RECT 164.365 50.355 165.455 50.470 ;
        POLYGON 165.455 50.640 165.475 50.355 165.455 50.355 ;
        POLYGON 166.895 50.640 166.920 50.640 166.920 50.385 ;
        RECT 166.920 50.530 168.995 50.640 ;
        POLYGON 168.995 50.805 169.020 50.530 168.995 50.530 ;
        POLYGON 171.625 50.805 171.655 50.805 171.655 50.540 ;
        RECT 171.655 50.530 175.670 50.805 ;
        RECT 166.920 50.355 169.020 50.530 ;
        RECT 164.365 50.160 165.475 50.355 ;
        POLYGON 165.475 50.355 165.485 50.160 165.475 50.160 ;
        POLYGON 166.920 50.355 166.930 50.355 166.930 50.280 ;
        RECT 166.930 50.320 169.020 50.355 ;
        POLYGON 169.020 50.530 169.040 50.320 169.020 50.320 ;
        POLYGON 171.655 50.530 171.675 50.530 171.675 50.350 ;
        RECT 171.675 50.320 175.670 50.530 ;
        RECT 166.930 50.160 169.040 50.320 ;
        RECT 164.365 50.155 165.485 50.160 ;
        RECT 162.700 50.130 163.535 50.155 ;
        RECT 161.580 50.110 162.090 50.130 ;
        POLYGON 160.675 50.085 160.680 50.085 160.680 49.900 ;
        POLYGON 160.680 49.900 160.680 49.680 160.675 49.680 ;
        RECT 160.680 49.680 160.975 50.085 ;
        RECT 160.675 49.650 160.975 49.680 ;
        POLYGON 160.675 49.645 160.675 49.460 160.665 49.460 ;
        RECT 160.675 49.460 160.955 49.650 ;
        RECT 149.765 49.285 159.955 49.445 ;
        POLYGON 159.955 49.445 159.975 49.445 159.955 49.285 ;
        POLYGON 160.665 49.445 160.665 49.405 160.660 49.405 ;
        RECT 160.665 49.405 160.955 49.460 ;
        POLYGON 160.660 49.385 160.660 49.290 160.650 49.290 ;
        RECT 160.660 49.290 160.955 49.405 ;
        RECT 149.765 49.250 159.930 49.285 ;
        RECT 117.195 49.170 149.080 49.250 ;
        POLYGON 149.080 49.250 149.090 49.170 149.080 49.170 ;
        POLYGON 149.765 49.250 149.780 49.250 149.780 49.170 ;
        RECT 117.195 48.860 149.090 49.170 ;
        RECT 149.780 49.160 159.930 49.250 ;
        POLYGON 149.090 49.160 149.135 48.860 149.090 48.860 ;
        POLYGON 149.780 49.160 149.800 49.160 149.800 49.065 ;
        RECT 149.800 49.130 159.930 49.160 ;
        POLYGON 159.930 49.285 159.955 49.285 159.930 49.130 ;
        POLYGON 160.650 49.285 160.650 49.240 160.645 49.240 ;
        RECT 160.650 49.275 160.955 49.290 ;
        POLYGON 160.955 49.650 160.975 49.650 160.955 49.275 ;
        POLYGON 161.580 50.110 161.585 50.110 161.585 49.825 ;
        RECT 161.585 49.975 162.090 50.110 ;
        POLYGON 162.090 50.130 162.100 49.975 162.090 49.975 ;
        POLYGON 161.585 49.825 161.585 49.585 161.580 49.585 ;
        RECT 161.585 49.675 162.100 49.975 ;
        RECT 161.585 49.585 162.090 49.675 ;
        POLYGON 161.580 49.545 161.580 49.425 161.570 49.425 ;
        RECT 161.580 49.425 162.090 49.585 ;
        POLYGON 161.570 49.425 161.570 49.320 161.565 49.320 ;
        RECT 161.570 49.380 162.090 49.425 ;
        POLYGON 162.090 49.675 162.100 49.675 162.090 49.380 ;
        POLYGON 162.700 50.130 162.705 50.130 162.705 49.825 ;
        RECT 162.705 50.005 163.535 50.130 ;
        POLYGON 163.535 50.155 163.540 50.005 163.535 50.005 ;
        POLYGON 164.365 50.155 164.375 50.155 164.375 50.060 ;
        RECT 164.375 50.070 165.485 50.155 ;
        POLYGON 165.485 50.160 165.490 50.070 165.485 50.070 ;
        POLYGON 166.930 50.160 166.935 50.160 166.935 50.110 ;
        RECT 164.375 50.005 165.490 50.070 ;
        RECT 166.935 50.025 169.040 50.160 ;
        POLYGON 169.040 50.320 169.060 50.025 169.040 50.025 ;
        POLYGON 171.675 50.320 171.695 50.320 171.695 50.055 ;
        RECT 171.695 50.025 175.670 50.320 ;
        RECT 166.935 50.005 169.060 50.025 ;
        POLYGON 162.705 49.825 162.705 49.510 162.700 49.510 ;
        RECT 162.705 49.510 163.540 50.005 ;
        POLYGON 163.540 50.005 163.545 49.730 163.540 49.730 ;
        POLYGON 162.700 49.475 162.700 49.380 162.695 49.380 ;
        RECT 162.700 49.380 163.540 49.510 ;
        RECT 161.570 49.320 162.065 49.380 ;
        POLYGON 161.565 49.320 161.565 49.275 161.560 49.275 ;
        RECT 161.565 49.275 162.065 49.320 ;
        RECT 160.650 49.240 160.925 49.275 ;
        POLYGON 160.645 49.240 160.645 49.180 160.635 49.180 ;
        RECT 160.645 49.180 160.925 49.240 ;
        POLYGON 160.635 49.180 160.635 49.130 160.630 49.130 ;
        RECT 160.635 49.130 160.925 49.180 ;
        RECT 149.800 49.065 159.910 49.130 ;
        POLYGON 149.800 49.065 149.805 49.065 149.805 49.045 ;
        RECT 149.805 49.045 159.910 49.065 ;
        POLYGON 149.805 49.045 149.845 49.045 149.845 48.865 ;
        RECT 149.845 49.030 159.910 49.045 ;
        POLYGON 159.910 49.130 159.930 49.130 159.910 49.030 ;
        POLYGON 160.630 49.130 160.630 49.030 160.615 49.030 ;
        RECT 160.630 49.030 160.925 49.130 ;
        RECT 149.845 48.975 159.900 49.030 ;
        POLYGON 159.900 49.030 159.910 49.030 159.900 48.975 ;
        POLYGON 160.615 49.020 160.615 48.990 160.610 48.990 ;
        RECT 160.615 48.990 160.925 49.030 ;
        RECT 117.195 48.850 149.135 48.860 ;
        POLYGON 149.135 48.860 149.140 48.850 149.135 48.850 ;
        RECT 149.845 48.850 159.870 48.975 ;
        RECT 117.195 48.785 149.140 48.850 ;
        POLYGON 149.140 48.850 149.155 48.785 149.140 48.785 ;
        POLYGON 149.845 48.850 149.850 48.850 149.850 48.845 ;
        RECT 149.850 48.845 159.870 48.850 ;
        POLYGON 149.850 48.845 149.855 48.845 149.855 48.835 ;
        RECT 149.855 48.825 159.870 48.845 ;
        POLYGON 159.870 48.975 159.900 48.975 159.870 48.825 ;
        POLYGON 160.610 48.975 160.610 48.955 160.605 48.955 ;
        RECT 160.610 48.955 160.925 48.990 ;
        POLYGON 160.605 48.955 160.605 48.825 160.580 48.825 ;
        RECT 160.605 48.910 160.925 48.955 ;
        POLYGON 160.925 49.275 160.955 49.275 160.925 48.910 ;
        POLYGON 161.560 49.265 161.560 49.035 161.530 49.035 ;
        RECT 161.560 49.085 162.065 49.275 ;
        POLYGON 162.065 49.380 162.090 49.380 162.065 49.085 ;
        POLYGON 162.695 49.380 162.695 49.190 162.685 49.190 ;
        RECT 162.695 49.300 163.540 49.380 ;
        POLYGON 163.540 49.730 163.545 49.730 163.540 49.300 ;
        POLYGON 164.375 50.005 164.380 50.005 164.380 49.620 ;
        POLYGON 164.380 49.620 164.380 49.500 164.375 49.500 ;
        RECT 164.380 49.500 165.490 50.005 ;
        POLYGON 164.375 49.500 164.375 49.340 164.370 49.340 ;
        RECT 164.375 49.490 165.490 49.500 ;
        POLYGON 165.490 50.005 165.500 49.490 165.490 49.490 ;
        RECT 164.375 49.340 165.485 49.490 ;
        RECT 162.695 49.190 163.505 49.300 ;
        POLYGON 162.685 49.190 162.685 49.140 162.680 49.140 ;
        RECT 162.685 49.140 163.505 49.190 ;
        POLYGON 162.680 49.140 162.680 49.095 162.675 49.095 ;
        RECT 162.680 49.095 163.505 49.140 ;
        RECT 161.560 49.035 162.030 49.085 ;
        POLYGON 161.530 49.035 161.530 48.985 161.525 48.985 ;
        RECT 161.530 48.985 162.030 49.035 ;
        POLYGON 161.525 48.985 161.525 48.920 161.515 48.920 ;
        RECT 161.525 48.920 162.030 48.985 ;
        RECT 160.605 48.825 160.880 48.910 ;
        POLYGON 149.855 48.825 149.865 48.825 149.865 48.785 ;
        RECT 149.865 48.785 159.830 48.825 ;
        RECT 117.195 48.625 149.155 48.785 ;
        POLYGON 149.155 48.785 149.185 48.625 149.155 48.625 ;
        POLYGON 149.865 48.785 149.905 48.785 149.905 48.645 ;
        RECT 149.905 48.675 159.830 48.785 ;
        POLYGON 159.830 48.825 159.870 48.825 159.830 48.675 ;
        POLYGON 160.580 48.820 160.580 48.800 160.575 48.800 ;
        RECT 160.580 48.800 160.880 48.825 ;
        POLYGON 160.575 48.800 160.575 48.735 160.560 48.735 ;
        RECT 160.575 48.735 160.880 48.800 ;
        POLYGON 160.560 48.735 160.560 48.720 160.555 48.720 ;
        RECT 160.560 48.720 160.880 48.735 ;
        POLYGON 160.555 48.720 160.555 48.675 160.545 48.675 ;
        RECT 160.555 48.675 160.880 48.720 ;
        RECT 149.905 48.645 159.795 48.675 ;
        POLYGON 149.905 48.645 149.910 48.645 149.910 48.625 ;
        RECT 149.910 48.625 159.795 48.645 ;
        RECT 117.195 48.615 149.185 48.625 ;
        RECT 54.910 48.295 112.180 48.615 ;
        POLYGON 112.180 48.615 112.260 48.295 112.180 48.295 ;
        POLYGON 117.195 48.615 117.200 48.615 117.200 48.400 ;
        RECT 117.200 48.560 149.185 48.615 ;
        POLYGON 149.185 48.625 149.200 48.560 149.185 48.560 ;
        POLYGON 149.910 48.625 149.920 48.625 149.920 48.595 ;
        RECT 149.920 48.595 159.795 48.625 ;
        POLYGON 149.920 48.595 149.930 48.595 149.930 48.560 ;
        RECT 149.930 48.570 159.795 48.595 ;
        POLYGON 159.795 48.675 159.830 48.675 159.795 48.570 ;
        POLYGON 160.545 48.675 160.545 48.585 160.525 48.585 ;
        RECT 160.545 48.585 160.880 48.675 ;
        RECT 160.525 48.580 160.880 48.585 ;
        POLYGON 160.880 48.910 160.925 48.910 160.880 48.580 ;
        POLYGON 161.515 48.910 161.515 48.755 161.490 48.755 ;
        RECT 161.515 48.795 162.030 48.920 ;
        POLYGON 162.030 49.085 162.065 49.085 162.030 48.795 ;
        POLYGON 162.675 49.085 162.675 48.875 162.650 48.875 ;
        RECT 162.675 48.875 163.505 49.095 ;
        POLYGON 162.650 48.875 162.650 48.820 162.645 48.820 ;
        RECT 162.650 48.870 163.505 48.875 ;
        POLYGON 163.505 49.300 163.540 49.300 163.505 48.870 ;
        POLYGON 164.370 49.300 164.370 49.180 164.365 49.180 ;
        RECT 164.370 49.180 165.485 49.340 ;
        POLYGON 164.365 49.180 164.365 49.005 164.350 49.005 ;
        RECT 164.365 49.005 165.485 49.180 ;
        POLYGON 164.350 49.005 164.350 48.875 164.340 48.875 ;
        RECT 164.350 48.915 165.485 49.005 ;
        POLYGON 165.485 49.490 165.500 49.490 165.485 48.915 ;
        POLYGON 166.935 50.005 166.960 50.005 166.960 49.350 ;
        RECT 166.960 49.830 169.060 50.005 ;
        POLYGON 169.060 50.025 169.070 49.830 169.060 49.830 ;
        POLYGON 171.695 50.025 171.710 50.025 171.710 49.835 ;
        RECT 171.710 49.850 175.670 50.025 ;
        POLYGON 175.670 50.970 175.685 49.850 175.670 49.850 ;
        POLYGON 182.700 50.970 182.765 50.970 182.765 50.435 ;
        RECT 182.765 50.435 197.200 50.970 ;
        POLYGON 182.765 50.435 182.795 50.435 182.795 50.185 ;
        RECT 182.795 50.185 197.200 50.435 ;
        POLYGON 182.795 50.185 182.815 50.185 182.815 49.900 ;
        RECT 182.815 49.850 197.200 50.185 ;
        RECT 171.710 49.830 175.685 49.850 ;
        RECT 166.960 49.490 169.070 49.830 ;
        POLYGON 169.070 49.830 169.080 49.490 169.070 49.490 ;
        POLYGON 171.710 49.830 171.725 49.830 171.725 49.615 ;
        RECT 171.725 49.490 175.685 49.830 ;
        POLYGON 166.960 49.350 166.960 48.915 166.955 48.915 ;
        RECT 166.960 48.915 169.080 49.490 ;
        POLYGON 169.080 49.490 169.085 49.340 169.080 49.340 ;
        RECT 164.350 48.875 165.475 48.915 ;
        RECT 162.650 48.820 163.450 48.870 ;
        POLYGON 162.645 48.820 162.645 48.795 162.640 48.795 ;
        RECT 162.645 48.795 163.450 48.820 ;
        RECT 161.515 48.755 161.985 48.795 ;
        POLYGON 161.490 48.755 161.490 48.580 161.455 48.580 ;
        RECT 161.490 48.580 161.985 48.755 ;
        RECT 149.930 48.560 159.785 48.570 ;
        RECT 117.200 48.545 149.200 48.560 ;
        POLYGON 149.200 48.560 149.205 48.545 149.200 48.545 ;
        POLYGON 149.930 48.560 149.935 48.560 149.935 48.545 ;
        RECT 149.935 48.545 159.785 48.560 ;
        RECT 117.200 48.295 149.205 48.545 ;
        RECT 54.910 45.915 112.260 48.295 ;
        POLYGON 54.910 45.915 55.200 45.915 55.200 45.200 ;
        RECT 55.200 45.840 112.260 45.915 ;
        POLYGON 112.260 48.295 112.885 45.840 112.260 45.840 ;
        POLYGON 117.200 48.295 117.205 48.295 117.205 48.135 ;
        RECT 117.205 48.270 149.205 48.295 ;
        POLYGON 149.205 48.545 149.275 48.270 149.205 48.270 ;
        POLYGON 149.935 48.545 149.965 48.545 149.965 48.450 ;
        RECT 149.965 48.525 159.785 48.545 ;
        POLYGON 159.785 48.570 159.795 48.570 159.785 48.525 ;
        POLYGON 160.525 48.570 160.525 48.535 160.515 48.535 ;
        RECT 160.525 48.550 160.875 48.580 ;
        POLYGON 160.875 48.580 160.880 48.580 160.875 48.550 ;
        POLYGON 161.455 48.580 161.455 48.560 161.450 48.560 ;
        RECT 161.455 48.560 161.985 48.580 ;
        RECT 160.525 48.535 160.820 48.550 ;
        RECT 149.965 48.485 159.770 48.525 ;
        POLYGON 159.770 48.525 159.785 48.525 159.770 48.485 ;
        POLYGON 160.515 48.525 160.515 48.515 160.510 48.515 ;
        RECT 160.515 48.515 160.820 48.535 ;
        POLYGON 160.510 48.515 160.510 48.485 160.500 48.485 ;
        RECT 160.510 48.485 160.820 48.515 ;
        RECT 149.965 48.450 159.735 48.485 ;
        POLYGON 149.965 48.450 149.995 48.450 149.995 48.370 ;
        RECT 149.995 48.380 159.735 48.450 ;
        POLYGON 159.735 48.485 159.770 48.485 159.735 48.380 ;
        POLYGON 160.500 48.480 160.500 48.385 160.475 48.385 ;
        RECT 160.500 48.385 160.820 48.485 ;
        RECT 149.995 48.370 159.680 48.380 ;
        POLYGON 149.995 48.370 150.025 48.370 150.025 48.280 ;
        RECT 150.025 48.270 159.680 48.370 ;
        RECT 117.205 48.180 149.275 48.270 ;
        POLYGON 149.275 48.270 149.305 48.180 149.275 48.180 ;
        POLYGON 150.025 48.270 150.030 48.270 150.030 48.265 ;
        RECT 150.030 48.265 159.680 48.270 ;
        POLYGON 150.030 48.265 150.060 48.265 150.060 48.185 ;
        RECT 150.060 48.235 159.680 48.265 ;
        POLYGON 159.680 48.380 159.735 48.380 159.680 48.235 ;
        POLYGON 160.475 48.380 160.475 48.365 160.470 48.365 ;
        RECT 160.475 48.365 160.820 48.385 ;
        POLYGON 160.470 48.365 160.470 48.315 160.455 48.315 ;
        RECT 160.470 48.315 160.820 48.365 ;
        POLYGON 160.455 48.315 160.455 48.295 160.450 48.295 ;
        RECT 160.455 48.295 160.820 48.315 ;
        POLYGON 160.450 48.295 160.450 48.235 160.430 48.235 ;
        RECT 160.450 48.235 160.820 48.295 ;
        RECT 150.060 48.180 159.625 48.235 ;
        RECT 117.205 48.035 149.305 48.180 ;
        POLYGON 149.305 48.180 149.350 48.035 149.305 48.035 ;
        POLYGON 150.060 48.180 150.075 48.180 150.075 48.150 ;
        RECT 150.075 48.150 159.625 48.180 ;
        POLYGON 150.075 48.150 150.105 48.150 150.105 48.080 ;
        RECT 150.105 48.095 159.625 48.150 ;
        POLYGON 159.625 48.235 159.680 48.235 159.625 48.095 ;
        POLYGON 160.430 48.235 160.430 48.155 160.405 48.155 ;
        RECT 160.430 48.210 160.820 48.235 ;
        POLYGON 160.820 48.550 160.875 48.550 160.820 48.210 ;
        POLYGON 161.450 48.550 161.450 48.475 161.430 48.475 ;
        RECT 161.450 48.505 161.985 48.560 ;
        POLYGON 161.985 48.795 162.030 48.795 161.985 48.505 ;
        POLYGON 162.640 48.785 162.640 48.720 162.630 48.720 ;
        RECT 162.640 48.720 163.450 48.795 ;
        POLYGON 162.630 48.720 162.630 48.555 162.605 48.555 ;
        RECT 162.630 48.555 163.450 48.720 ;
        POLYGON 162.605 48.555 162.605 48.510 162.600 48.510 ;
        RECT 162.605 48.510 163.450 48.555 ;
        RECT 161.450 48.475 161.925 48.505 ;
        POLYGON 161.430 48.475 161.430 48.425 161.420 48.425 ;
        RECT 161.430 48.425 161.925 48.475 ;
        POLYGON 161.420 48.425 161.420 48.215 161.365 48.215 ;
        RECT 161.420 48.220 161.925 48.425 ;
        POLYGON 161.925 48.505 161.985 48.505 161.925 48.220 ;
        POLYGON 162.600 48.505 162.600 48.445 162.585 48.445 ;
        RECT 162.600 48.445 163.450 48.510 ;
        POLYGON 163.450 48.870 163.505 48.870 163.450 48.445 ;
        POLYGON 164.340 48.870 164.340 48.740 164.330 48.740 ;
        RECT 164.340 48.745 165.475 48.875 ;
        POLYGON 165.475 48.915 165.485 48.915 165.475 48.795 ;
        RECT 166.955 48.845 169.080 48.915 ;
        POLYGON 169.080 49.340 169.085 49.340 169.080 48.845 ;
        POLYGON 171.725 49.490 171.745 49.490 171.745 48.880 ;
        RECT 164.340 48.740 165.445 48.745 ;
        POLYGON 164.330 48.740 164.330 48.550 164.305 48.550 ;
        RECT 164.330 48.550 165.445 48.740 ;
        POLYGON 164.305 48.550 164.305 48.445 164.290 48.445 ;
        RECT 164.305 48.445 165.445 48.550 ;
        POLYGON 162.585 48.445 162.585 48.240 162.550 48.240 ;
        RECT 162.585 48.385 163.440 48.445 ;
        POLYGON 163.440 48.445 163.450 48.445 163.440 48.385 ;
        POLYGON 164.290 48.425 164.290 48.385 164.285 48.385 ;
        RECT 164.290 48.385 165.445 48.445 ;
        RECT 162.585 48.240 163.395 48.385 ;
        POLYGON 162.550 48.240 162.550 48.220 162.545 48.220 ;
        RECT 162.550 48.220 163.395 48.240 ;
        RECT 161.420 48.215 161.905 48.220 ;
        RECT 160.430 48.155 160.760 48.210 ;
        POLYGON 160.405 48.155 160.405 48.095 160.385 48.095 ;
        RECT 160.405 48.095 160.760 48.155 ;
        RECT 150.105 48.090 159.620 48.095 ;
        POLYGON 159.620 48.095 159.625 48.095 159.620 48.090 ;
        RECT 150.105 48.080 159.565 48.090 ;
        POLYGON 150.105 48.080 150.120 48.080 150.120 48.040 ;
        RECT 150.120 48.035 159.565 48.080 ;
        RECT 117.205 47.985 149.350 48.035 ;
        POLYGON 149.350 48.035 149.365 47.985 149.350 47.985 ;
        POLYGON 150.120 48.035 150.140 48.035 150.140 47.990 ;
        RECT 150.140 47.985 159.565 48.035 ;
        RECT 117.205 47.965 149.365 47.985 ;
        POLYGON 149.365 47.985 149.370 47.965 149.365 47.965 ;
        POLYGON 150.140 47.985 150.150 47.985 150.150 47.965 ;
        RECT 150.150 47.965 159.565 47.985 ;
        POLYGON 159.565 48.090 159.620 48.090 159.565 47.965 ;
        POLYGON 160.385 48.090 160.385 48.080 160.380 48.080 ;
        RECT 160.385 48.080 160.760 48.095 ;
        POLYGON 160.380 48.080 160.380 47.965 160.335 47.965 ;
        RECT 160.380 47.965 160.760 48.080 ;
        RECT 117.205 47.870 149.370 47.965 ;
        POLYGON 117.205 47.870 117.220 47.870 117.220 47.335 ;
        RECT 117.220 47.805 149.370 47.870 ;
        POLYGON 149.370 47.965 149.430 47.805 149.370 47.805 ;
        POLYGON 150.150 47.965 150.180 47.965 150.180 47.895 ;
        RECT 150.180 47.950 159.560 47.965 ;
        POLYGON 159.560 47.965 159.565 47.965 159.560 47.950 ;
        POLYGON 160.335 47.960 160.335 47.950 160.330 47.950 ;
        RECT 160.335 47.950 160.760 47.965 ;
        RECT 150.180 47.895 159.490 47.950 ;
        POLYGON 150.180 47.895 150.225 47.895 150.225 47.805 ;
        RECT 150.225 47.810 159.490 47.895 ;
        POLYGON 159.490 47.950 159.560 47.950 159.490 47.810 ;
        RECT 160.330 47.945 160.760 47.950 ;
        POLYGON 160.760 48.210 160.820 48.210 160.760 47.945 ;
        POLYGON 161.365 48.210 161.365 48.195 161.360 48.195 ;
        RECT 161.365 48.195 161.905 48.215 ;
        POLYGON 161.360 48.195 161.360 48.150 161.350 48.150 ;
        RECT 161.360 48.150 161.905 48.195 ;
        POLYGON 161.350 48.150 161.350 48.075 161.325 48.075 ;
        RECT 161.350 48.145 161.905 48.150 ;
        POLYGON 161.905 48.220 161.925 48.220 161.905 48.145 ;
        POLYGON 162.545 48.220 162.545 48.200 162.540 48.200 ;
        RECT 162.545 48.200 163.395 48.220 ;
        POLYGON 162.540 48.200 162.540 48.145 162.525 48.145 ;
        RECT 162.540 48.160 163.395 48.200 ;
        POLYGON 163.395 48.385 163.440 48.385 163.395 48.160 ;
        POLYGON 164.285 48.385 164.285 48.300 164.275 48.300 ;
        RECT 164.285 48.340 165.445 48.385 ;
        POLYGON 165.445 48.745 165.475 48.745 165.445 48.340 ;
        POLYGON 166.955 48.520 166.955 48.380 166.950 48.380 ;
        RECT 166.955 48.380 169.060 48.845 ;
        RECT 166.950 48.355 169.060 48.380 ;
        POLYGON 169.060 48.845 169.080 48.845 169.060 48.355 ;
        POLYGON 171.745 48.845 171.745 48.385 171.735 48.385 ;
        RECT 171.745 48.385 175.685 49.490 ;
        RECT 164.285 48.300 165.385 48.340 ;
        POLYGON 164.275 48.300 164.275 48.225 164.260 48.225 ;
        RECT 164.275 48.225 165.385 48.300 ;
        POLYGON 164.260 48.225 164.260 48.170 164.250 48.170 ;
        RECT 164.260 48.170 165.385 48.225 ;
        RECT 162.540 48.145 163.370 48.160 ;
        RECT 161.350 48.075 161.855 48.145 ;
        POLYGON 161.325 48.075 161.325 47.945 161.285 47.945 ;
        RECT 161.325 47.945 161.855 48.075 ;
        POLYGON 160.330 47.945 160.330 47.865 160.300 47.865 ;
        RECT 160.330 47.885 160.745 47.945 ;
        POLYGON 160.745 47.945 160.760 47.945 160.745 47.885 ;
        RECT 161.285 47.935 161.855 47.945 ;
        POLYGON 161.855 48.145 161.905 48.145 161.855 47.935 ;
        POLYGON 162.525 48.140 162.525 47.935 162.475 47.935 ;
        RECT 162.525 48.020 163.370 48.145 ;
        POLYGON 163.370 48.160 163.395 48.160 163.370 48.020 ;
        POLYGON 164.250 48.160 164.250 48.110 164.240 48.110 ;
        RECT 164.250 48.110 165.385 48.170 ;
        POLYGON 164.240 48.110 164.240 48.025 164.225 48.025 ;
        RECT 164.240 48.025 165.385 48.110 ;
        RECT 162.525 47.935 163.270 48.020 ;
        POLYGON 161.285 47.935 161.285 47.890 161.270 47.890 ;
        RECT 161.285 47.920 161.850 47.935 ;
        POLYGON 161.850 47.935 161.855 47.935 161.850 47.920 ;
        RECT 161.285 47.890 161.770 47.920 ;
        RECT 160.330 47.865 160.710 47.885 ;
        POLYGON 160.300 47.865 160.300 47.855 160.295 47.855 ;
        RECT 160.300 47.855 160.710 47.865 ;
        POLYGON 160.295 47.855 160.295 47.815 160.280 47.815 ;
        RECT 160.295 47.815 160.710 47.855 ;
        RECT 150.225 47.805 159.415 47.810 ;
        RECT 117.220 47.710 149.430 47.805 ;
        POLYGON 149.430 47.805 149.465 47.710 149.430 47.710 ;
        POLYGON 150.225 47.805 150.265 47.805 150.265 47.725 ;
        RECT 150.265 47.720 159.415 47.805 ;
        POLYGON 150.265 47.720 150.270 47.720 150.270 47.710 ;
        RECT 150.270 47.710 159.415 47.720 ;
        RECT 117.220 47.685 149.465 47.710 ;
        POLYGON 149.465 47.710 149.475 47.685 149.465 47.685 ;
        POLYGON 150.270 47.710 150.280 47.710 150.280 47.690 ;
        RECT 150.280 47.685 159.415 47.710 ;
        RECT 117.220 47.480 149.475 47.685 ;
        POLYGON 149.475 47.685 149.560 47.480 149.475 47.480 ;
        POLYGON 150.280 47.685 150.340 47.685 150.340 47.575 ;
        RECT 150.340 47.675 159.415 47.685 ;
        POLYGON 159.415 47.810 159.490 47.810 159.415 47.675 ;
        POLYGON 160.280 47.810 160.280 47.735 160.250 47.735 ;
        RECT 160.280 47.765 160.710 47.815 ;
        POLYGON 160.710 47.885 160.745 47.885 160.710 47.765 ;
        POLYGON 161.270 47.885 161.270 47.875 161.265 47.875 ;
        RECT 161.270 47.875 161.770 47.890 ;
        POLYGON 161.265 47.875 161.265 47.765 161.225 47.765 ;
        RECT 161.265 47.765 161.770 47.875 ;
        RECT 160.280 47.735 160.705 47.765 ;
        POLYGON 160.250 47.735 160.250 47.680 160.225 47.680 ;
        RECT 160.250 47.730 160.705 47.735 ;
        POLYGON 160.705 47.765 160.710 47.765 160.705 47.730 ;
        POLYGON 161.225 47.765 161.225 47.735 161.215 47.735 ;
        RECT 161.225 47.735 161.770 47.765 ;
        RECT 160.250 47.680 160.660 47.730 ;
        RECT 150.340 47.575 159.335 47.675 ;
        POLYGON 150.340 47.575 150.355 47.575 150.355 47.550 ;
        RECT 150.355 47.550 159.335 47.575 ;
        POLYGON 150.355 47.550 150.370 47.550 150.370 47.520 ;
        RECT 150.370 47.540 159.335 47.550 ;
        POLYGON 159.335 47.675 159.415 47.675 159.335 47.540 ;
        POLYGON 160.225 47.675 160.225 47.655 160.215 47.655 ;
        RECT 160.225 47.655 160.660 47.680 ;
        POLYGON 160.215 47.655 160.215 47.640 160.205 47.640 ;
        RECT 160.215 47.640 160.660 47.655 ;
        POLYGON 160.205 47.640 160.205 47.550 160.165 47.550 ;
        RECT 160.205 47.585 160.660 47.640 ;
        POLYGON 160.660 47.730 160.705 47.730 160.660 47.585 ;
        POLYGON 161.215 47.730 161.215 47.665 161.190 47.665 ;
        RECT 161.215 47.665 161.770 47.735 ;
        POLYGON 161.190 47.665 161.190 47.605 161.170 47.605 ;
        RECT 161.190 47.655 161.770 47.665 ;
        POLYGON 161.770 47.920 161.850 47.920 161.770 47.655 ;
        POLYGON 162.475 47.920 162.475 47.890 162.465 47.890 ;
        RECT 162.475 47.890 163.270 47.935 ;
        POLYGON 162.465 47.890 162.465 47.690 162.410 47.690 ;
        RECT 162.465 47.690 163.270 47.890 ;
        POLYGON 162.410 47.690 162.410 47.655 162.400 47.655 ;
        RECT 162.410 47.655 163.270 47.690 ;
        RECT 161.190 47.605 161.675 47.655 ;
        POLYGON 161.170 47.605 161.170 47.585 161.160 47.585 ;
        RECT 161.170 47.585 161.675 47.605 ;
        RECT 160.205 47.550 160.585 47.585 ;
        POLYGON 160.165 47.550 160.165 47.540 160.160 47.540 ;
        RECT 160.165 47.540 160.585 47.550 ;
        RECT 150.370 47.520 159.320 47.540 ;
        POLYGON 150.370 47.520 150.390 47.520 150.390 47.485 ;
        RECT 150.390 47.515 159.320 47.520 ;
        POLYGON 159.320 47.540 159.335 47.540 159.320 47.515 ;
        POLYGON 160.160 47.540 160.160 47.520 160.150 47.520 ;
        RECT 160.160 47.520 160.585 47.540 ;
        RECT 150.390 47.480 159.300 47.515 ;
        POLYGON 159.300 47.515 159.320 47.515 159.300 47.480 ;
        POLYGON 160.150 47.515 160.150 47.480 160.130 47.480 ;
        RECT 160.150 47.480 160.585 47.520 ;
        RECT 117.220 47.445 149.565 47.480 ;
        POLYGON 149.565 47.480 149.580 47.445 149.565 47.445 ;
        POLYGON 150.390 47.480 150.410 47.480 150.410 47.450 ;
        RECT 150.410 47.445 159.250 47.480 ;
        RECT 117.220 47.420 149.580 47.445 ;
        POLYGON 149.580 47.445 149.590 47.420 149.580 47.420 ;
        POLYGON 150.410 47.445 150.425 47.445 150.425 47.420 ;
        RECT 150.425 47.420 159.250 47.445 ;
        RECT 117.220 47.250 149.590 47.420 ;
        POLYGON 149.590 47.420 149.670 47.250 149.590 47.250 ;
        POLYGON 150.425 47.420 150.450 47.420 150.450 47.380 ;
        RECT 150.450 47.405 159.250 47.420 ;
        POLYGON 159.250 47.480 159.300 47.480 159.250 47.405 ;
        POLYGON 160.130 47.475 160.130 47.405 160.095 47.405 ;
        RECT 160.130 47.405 160.585 47.480 ;
        RECT 150.450 47.380 159.130 47.405 ;
        POLYGON 150.450 47.380 150.485 47.380 150.485 47.325 ;
        RECT 150.485 47.325 159.130 47.380 ;
        POLYGON 150.485 47.325 150.530 47.325 150.530 47.250 ;
        RECT 150.530 47.250 159.130 47.325 ;
        RECT 117.220 47.245 149.670 47.250 ;
        POLYGON 149.670 47.250 149.675 47.245 149.670 47.245 ;
        RECT 117.220 47.220 149.675 47.245 ;
        POLYGON 150.530 47.250 150.535 47.250 150.535 47.240 ;
        RECT 150.535 47.240 159.130 47.250 ;
        POLYGON 149.675 47.240 149.685 47.220 149.675 47.220 ;
        POLYGON 150.535 47.240 150.550 47.240 150.550 47.220 ;
        RECT 150.550 47.230 159.130 47.240 ;
        POLYGON 159.130 47.405 159.250 47.405 159.130 47.230 ;
        POLYGON 160.095 47.405 160.095 47.325 160.055 47.325 ;
        RECT 160.095 47.375 160.585 47.405 ;
        POLYGON 160.585 47.585 160.660 47.585 160.585 47.375 ;
        POLYGON 161.160 47.580 161.160 47.385 161.080 47.385 ;
        RECT 161.160 47.385 161.675 47.585 ;
        POLYGON 161.080 47.385 161.080 47.380 161.075 47.380 ;
        RECT 161.080 47.380 161.675 47.385 ;
        POLYGON 161.675 47.655 161.770 47.655 161.675 47.380 ;
        POLYGON 162.400 47.655 162.400 47.615 162.390 47.615 ;
        RECT 162.400 47.615 163.270 47.655 ;
        POLYGON 162.390 47.615 162.390 47.585 162.380 47.585 ;
        RECT 162.390 47.595 163.270 47.615 ;
        POLYGON 163.270 48.020 163.370 48.020 163.270 47.595 ;
        POLYGON 164.225 48.020 164.225 47.860 164.195 47.860 ;
        RECT 164.225 47.860 165.385 48.025 ;
        POLYGON 164.195 47.860 164.195 47.680 164.155 47.680 ;
        RECT 164.195 47.780 165.385 47.860 ;
        POLYGON 165.385 48.340 165.445 48.340 165.385 47.780 ;
        POLYGON 166.950 48.340 166.950 47.830 166.930 47.830 ;
        RECT 166.950 47.860 169.020 48.355 ;
        POLYGON 169.020 48.355 169.060 48.355 169.020 47.860 ;
        POLYGON 171.735 48.355 171.735 48.140 171.730 48.140 ;
        RECT 171.735 48.140 175.685 48.385 ;
        POLYGON 175.685 49.850 175.700 48.380 175.685 48.380 ;
        POLYGON 182.815 49.850 182.900 49.850 182.900 48.705 ;
        RECT 182.900 49.260 197.200 49.850 ;
        POLYGON 197.200 51.030 197.510 49.260 197.200 49.260 ;
        POLYGON 206.775 51.030 206.795 51.030 206.795 50.930 ;
        RECT 206.795 50.930 222.230 51.030 ;
        RECT 182.900 48.835 197.510 49.260 ;
        POLYGON 206.795 50.930 207.110 50.930 207.110 49.250 ;
        RECT 207.110 50.495 222.230 50.930 ;
        POLYGON 222.230 52.590 222.255 50.495 222.230 50.495 ;
        POLYGON 229.205 52.590 229.205 51.355 229.190 51.355 ;
        RECT 229.205 52.080 233.225 52.590 ;
        POLYGON 233.225 52.590 233.270 52.590 233.225 52.080 ;
        POLYGON 236.100 52.590 236.100 52.240 236.055 52.240 ;
        RECT 236.100 52.455 238.110 52.590 ;
        POLYGON 238.110 52.590 238.135 52.590 238.110 52.455 ;
        POLYGON 239.770 52.580 239.770 52.530 239.760 52.530 ;
        RECT 239.770 52.530 240.820 52.590 ;
        POLYGON 239.760 52.510 239.760 52.455 239.750 52.455 ;
        RECT 239.760 52.455 240.820 52.530 ;
        RECT 236.100 52.300 238.090 52.455 ;
        POLYGON 238.090 52.455 238.110 52.455 238.090 52.300 ;
        POLYGON 239.750 52.440 239.750 52.305 239.730 52.305 ;
        RECT 239.750 52.385 240.820 52.455 ;
        POLYGON 240.820 52.590 240.865 52.590 240.820 52.385 ;
        POLYGON 241.895 52.590 241.895 52.565 241.885 52.565 ;
        RECT 241.895 52.585 242.720 52.600 ;
        POLYGON 242.720 52.780 242.780 52.780 242.720 52.590 ;
        POLYGON 243.450 52.780 243.450 52.745 243.435 52.745 ;
        RECT 243.450 52.745 243.975 52.785 ;
        POLYGON 243.435 52.745 243.435 52.635 243.395 52.635 ;
        RECT 243.435 52.735 243.975 52.745 ;
        POLYGON 243.975 52.785 243.995 52.785 243.975 52.735 ;
        POLYGON 244.565 52.785 244.565 52.735 244.540 52.735 ;
        RECT 244.565 52.735 245.385 52.785 ;
        RECT 243.435 52.695 243.955 52.735 ;
        POLYGON 243.955 52.735 243.975 52.735 243.955 52.695 ;
        POLYGON 244.540 52.735 244.540 52.725 244.535 52.725 ;
        RECT 244.540 52.725 245.385 52.735 ;
        POLYGON 244.535 52.725 244.535 52.700 244.525 52.700 ;
        RECT 244.535 52.700 245.385 52.725 ;
        RECT 243.435 52.635 243.910 52.695 ;
        POLYGON 243.395 52.635 243.395 52.590 243.375 52.590 ;
        RECT 243.395 52.590 243.910 52.635 ;
        POLYGON 243.910 52.695 243.955 52.695 243.910 52.595 ;
        POLYGON 244.525 52.695 244.525 52.615 244.490 52.615 ;
        RECT 244.525 52.660 245.385 52.700 ;
        POLYGON 245.385 52.785 245.465 52.785 245.385 52.660 ;
        POLYGON 254.090 52.785 254.110 52.785 254.110 52.765 ;
        RECT 254.110 52.765 254.815 52.785 ;
        POLYGON 254.110 52.765 254.185 52.765 254.185 52.665 ;
        RECT 254.185 52.725 254.815 52.765 ;
        POLYGON 254.815 52.860 254.900 52.725 254.815 52.725 ;
        POLYGON 255.350 52.860 255.360 52.860 255.360 52.850 ;
        RECT 255.360 52.850 255.805 52.860 ;
        POLYGON 255.360 52.850 255.385 52.850 255.385 52.815 ;
        RECT 255.385 52.840 255.805 52.850 ;
        POLYGON 255.805 52.875 255.825 52.840 255.805 52.840 ;
        POLYGON 256.430 52.875 256.435 52.875 256.435 52.865 ;
        RECT 256.435 52.865 257.060 52.875 ;
        POLYGON 256.435 52.865 256.445 52.865 256.445 52.840 ;
        RECT 256.445 52.840 257.060 52.865 ;
        RECT 255.385 52.825 255.825 52.840 ;
        POLYGON 255.825 52.840 255.830 52.825 255.825 52.825 ;
        POLYGON 256.445 52.840 256.450 52.840 256.450 52.830 ;
        RECT 256.450 52.825 257.060 52.840 ;
        RECT 255.385 52.815 255.830 52.825 ;
        POLYGON 255.385 52.815 255.390 52.815 255.390 52.805 ;
        RECT 255.390 52.805 255.830 52.815 ;
        POLYGON 255.390 52.805 255.435 52.805 255.435 52.725 ;
        RECT 255.435 52.725 255.830 52.805 ;
        RECT 254.185 52.695 254.900 52.725 ;
        POLYGON 254.900 52.725 254.920 52.695 254.900 52.695 ;
        POLYGON 255.435 52.725 255.445 52.725 255.445 52.710 ;
        RECT 255.445 52.710 255.830 52.725 ;
        POLYGON 255.445 52.710 255.450 52.710 255.450 52.700 ;
        RECT 255.450 52.695 255.830 52.710 ;
        RECT 254.185 52.660 254.920 52.695 ;
        RECT 244.525 52.630 245.370 52.660 ;
        POLYGON 245.370 52.660 245.385 52.660 245.370 52.630 ;
        POLYGON 254.185 52.660 254.210 52.660 254.210 52.630 ;
        RECT 254.210 52.630 254.920 52.660 ;
        RECT 244.525 52.625 245.365 52.630 ;
        POLYGON 245.365 52.630 245.370 52.630 245.365 52.625 ;
        POLYGON 254.210 52.630 254.215 52.630 254.215 52.625 ;
        RECT 254.215 52.625 254.920 52.630 ;
        RECT 244.525 52.615 245.345 52.625 ;
        POLYGON 244.490 52.615 244.490 52.600 244.485 52.600 ;
        RECT 244.490 52.600 245.345 52.615 ;
        RECT 241.895 52.565 242.710 52.585 ;
        POLYGON 241.885 52.565 241.885 52.555 241.880 52.555 ;
        RECT 241.885 52.555 242.710 52.565 ;
        POLYGON 242.710 52.585 242.720 52.585 242.710 52.555 ;
        POLYGON 243.375 52.590 243.375 52.560 243.365 52.560 ;
        RECT 243.375 52.560 243.875 52.590 ;
        POLYGON 241.880 52.555 241.880 52.390 241.835 52.390 ;
        RECT 241.880 52.515 242.695 52.555 ;
        POLYGON 242.695 52.555 242.710 52.555 242.695 52.515 ;
        POLYGON 243.365 52.555 243.365 52.515 243.350 52.515 ;
        RECT 243.365 52.515 243.875 52.560 ;
        POLYGON 243.875 52.590 243.910 52.590 243.875 52.515 ;
        POLYGON 244.485 52.595 244.485 52.590 244.480 52.590 ;
        RECT 244.485 52.590 245.345 52.600 ;
        POLYGON 245.345 52.625 245.365 52.625 245.345 52.590 ;
        POLYGON 254.215 52.625 254.235 52.625 254.235 52.595 ;
        RECT 254.235 52.610 254.920 52.625 ;
        POLYGON 254.920 52.695 254.965 52.610 254.920 52.610 ;
        POLYGON 255.450 52.695 255.470 52.695 255.470 52.675 ;
        RECT 255.470 52.675 255.830 52.695 ;
        POLYGON 255.470 52.675 255.500 52.675 255.500 52.620 ;
        RECT 255.500 52.620 255.830 52.675 ;
        POLYGON 255.500 52.620 255.505 52.620 255.505 52.610 ;
        RECT 255.505 52.615 255.830 52.620 ;
        POLYGON 255.830 52.825 255.940 52.615 255.830 52.615 ;
        POLYGON 256.450 52.825 256.485 52.825 256.485 52.755 ;
        RECT 256.485 52.800 257.060 52.825 ;
        POLYGON 257.060 52.895 257.100 52.800 257.060 52.800 ;
        POLYGON 257.870 52.895 257.910 52.895 257.910 52.810 ;
        RECT 257.910 52.800 258.830 52.895 ;
        RECT 256.485 52.755 257.100 52.800 ;
        POLYGON 256.485 52.755 256.490 52.755 256.490 52.740 ;
        RECT 256.490 52.740 257.100 52.755 ;
        POLYGON 256.490 52.740 256.495 52.740 256.495 52.730 ;
        RECT 256.495 52.730 257.100 52.740 ;
        POLYGON 256.495 52.730 256.505 52.730 256.505 52.715 ;
        RECT 256.505 52.715 257.100 52.730 ;
        POLYGON 256.505 52.715 256.530 52.715 256.530 52.650 ;
        RECT 256.530 52.650 257.100 52.715 ;
        POLYGON 256.530 52.650 256.535 52.650 256.535 52.635 ;
        RECT 256.535 52.635 257.100 52.650 ;
        POLYGON 256.535 52.635 256.545 52.635 256.545 52.615 ;
        RECT 256.545 52.615 257.100 52.635 ;
        RECT 255.505 52.610 255.940 52.615 ;
        RECT 254.235 52.590 254.965 52.610 ;
        POLYGON 254.965 52.610 254.975 52.590 254.965 52.590 ;
        POLYGON 255.505 52.610 255.515 52.610 255.515 52.590 ;
        RECT 255.515 52.595 255.940 52.610 ;
        POLYGON 255.940 52.615 255.950 52.595 255.940 52.595 ;
        POLYGON 256.545 52.615 256.555 52.615 256.555 52.595 ;
        RECT 255.515 52.590 255.950 52.595 ;
        RECT 256.555 52.590 257.100 52.615 ;
        POLYGON 257.100 52.800 257.180 52.590 257.100 52.590 ;
        POLYGON 257.910 52.800 257.955 52.800 257.955 52.705 ;
        RECT 257.955 52.705 258.830 52.800 ;
        POLYGON 257.955 52.705 257.975 52.705 257.975 52.660 ;
        RECT 257.975 52.665 258.830 52.705 ;
        POLYGON 258.830 52.910 258.920 52.665 258.830 52.665 ;
        POLYGON 260.065 52.910 260.080 52.910 260.080 52.870 ;
        RECT 260.080 52.870 261.495 52.910 ;
        POLYGON 260.080 52.870 260.100 52.870 260.100 52.800 ;
        RECT 260.100 52.825 261.495 52.870 ;
        POLYGON 261.495 52.975 261.535 52.825 261.495 52.825 ;
        POLYGON 263.550 52.975 263.590 52.975 263.590 52.835 ;
        RECT 263.590 52.970 266.245 52.975 ;
        POLYGON 266.245 53.015 266.255 52.970 266.245 52.970 ;
        POLYGON 270.495 53.015 270.500 53.015 270.500 53.010 ;
        RECT 270.500 53.010 277.290 53.015 ;
        POLYGON 270.500 53.010 270.505 53.010 270.505 52.975 ;
        RECT 270.505 52.970 277.290 53.010 ;
        RECT 263.590 52.825 266.255 52.970 ;
        RECT 260.100 52.800 261.535 52.825 ;
        POLYGON 260.100 52.800 260.130 52.800 260.130 52.675 ;
        RECT 260.130 52.665 261.535 52.800 ;
        RECT 257.975 52.660 258.920 52.665 ;
        POLYGON 257.975 52.660 257.995 52.660 257.995 52.600 ;
        RECT 257.995 52.650 258.920 52.660 ;
        POLYGON 258.920 52.665 258.925 52.650 258.920 52.650 ;
        POLYGON 260.130 52.665 260.135 52.665 260.135 52.650 ;
        RECT 260.135 52.650 261.535 52.665 ;
        RECT 257.995 52.615 258.925 52.650 ;
        POLYGON 258.925 52.650 258.935 52.615 258.925 52.615 ;
        POLYGON 260.135 52.650 260.140 52.650 260.140 52.630 ;
        RECT 260.140 52.630 261.535 52.650 ;
        POLYGON 261.535 52.825 261.580 52.630 261.535 52.630 ;
        POLYGON 263.590 52.825 263.600 52.825 263.600 52.800 ;
        RECT 263.600 52.800 266.255 52.825 ;
        POLYGON 263.600 52.800 263.640 52.800 263.640 52.635 ;
        RECT 263.640 52.630 266.255 52.800 ;
        RECT 260.140 52.615 261.580 52.630 ;
        RECT 257.995 52.595 258.935 52.615 ;
        POLYGON 258.935 52.615 258.940 52.595 258.935 52.595 ;
        RECT 257.995 52.590 258.940 52.595 ;
        POLYGON 260.140 52.615 260.150 52.615 260.150 52.590 ;
        RECT 260.150 52.590 261.580 52.615 ;
        POLYGON 261.580 52.630 261.590 52.590 261.580 52.590 ;
        POLYGON 263.640 52.630 263.650 52.630 263.650 52.595 ;
        RECT 263.650 52.600 266.255 52.630 ;
        POLYGON 266.255 52.970 266.340 52.600 266.255 52.600 ;
        POLYGON 270.505 52.970 270.550 52.970 270.550 52.670 ;
        RECT 270.550 52.670 277.290 52.970 ;
        RECT 263.650 52.590 266.340 52.600 ;
        POLYGON 270.550 52.670 270.555 52.670 270.555 52.595 ;
        RECT 270.555 52.610 277.290 52.670 ;
        POLYGON 277.290 53.320 277.425 52.610 277.290 52.610 ;
        RECT 270.555 52.590 277.425 52.610 ;
        POLYGON 244.480 52.585 244.480 52.540 244.465 52.540 ;
        RECT 244.480 52.575 245.335 52.590 ;
        POLYGON 245.335 52.590 245.345 52.590 245.335 52.575 ;
        POLYGON 254.235 52.590 254.245 52.590 254.245 52.580 ;
        RECT 254.245 52.575 254.975 52.590 ;
        RECT 244.480 52.540 245.280 52.575 ;
        POLYGON 244.465 52.540 244.465 52.515 244.455 52.515 ;
        RECT 244.465 52.515 245.280 52.540 ;
        RECT 241.880 52.390 242.625 52.515 ;
        RECT 239.750 52.305 240.775 52.385 ;
        RECT 236.100 52.240 238.035 52.300 ;
        POLYGON 236.055 52.240 236.055 52.170 236.045 52.170 ;
        RECT 236.055 52.170 238.035 52.240 ;
        POLYGON 236.045 52.170 236.045 52.105 236.040 52.105 ;
        RECT 236.045 52.105 238.035 52.170 ;
        RECT 229.205 51.865 233.220 52.080 ;
        POLYGON 233.220 52.080 233.225 52.080 233.220 51.865 ;
        POLYGON 236.040 52.080 236.040 51.865 236.020 51.865 ;
        RECT 236.040 51.915 238.035 52.105 ;
        POLYGON 238.035 52.300 238.090 52.300 238.035 51.915 ;
        POLYGON 239.730 52.300 239.730 52.030 239.690 52.030 ;
        RECT 239.730 52.110 240.775 52.305 ;
        POLYGON 240.775 52.385 240.820 52.385 240.775 52.110 ;
        POLYGON 241.835 52.385 241.835 52.355 241.825 52.355 ;
        RECT 241.835 52.355 242.625 52.390 ;
        POLYGON 241.825 52.355 241.825 52.245 241.790 52.245 ;
        RECT 241.825 52.270 242.625 52.355 ;
        POLYGON 242.625 52.515 242.695 52.515 242.625 52.270 ;
        POLYGON 243.350 52.515 243.350 52.365 243.300 52.365 ;
        RECT 243.350 52.505 243.875 52.515 ;
        RECT 243.350 52.455 243.850 52.505 ;
        POLYGON 243.850 52.505 243.875 52.505 243.850 52.455 ;
        POLYGON 244.455 52.515 244.455 52.455 244.430 52.455 ;
        RECT 244.455 52.470 245.280 52.515 ;
        POLYGON 245.280 52.575 245.335 52.575 245.280 52.470 ;
        POLYGON 254.245 52.575 254.305 52.575 254.305 52.495 ;
        RECT 254.305 52.550 254.975 52.575 ;
        POLYGON 254.975 52.590 255.000 52.550 254.975 52.550 ;
        POLYGON 255.515 52.590 255.520 52.590 255.520 52.580 ;
        RECT 255.520 52.580 255.950 52.590 ;
        POLYGON 255.520 52.580 255.530 52.580 255.530 52.555 ;
        RECT 255.530 52.575 255.950 52.580 ;
        POLYGON 255.950 52.590 255.960 52.575 255.950 52.575 ;
        POLYGON 256.555 52.590 256.565 52.590 256.565 52.575 ;
        RECT 255.530 52.550 255.960 52.575 ;
        RECT 254.305 52.510 255.000 52.550 ;
        POLYGON 255.000 52.550 255.020 52.510 255.000 52.510 ;
        POLYGON 255.530 52.550 255.540 52.550 255.540 52.535 ;
        RECT 255.540 52.535 255.960 52.550 ;
        POLYGON 255.540 52.535 255.555 52.535 255.555 52.510 ;
        RECT 255.555 52.510 255.960 52.535 ;
        RECT 254.305 52.495 255.020 52.510 ;
        POLYGON 254.305 52.495 254.310 52.495 254.310 52.480 ;
        RECT 254.310 52.480 255.020 52.495 ;
        POLYGON 254.315 52.480 254.320 52.480 254.320 52.470 ;
        RECT 254.320 52.470 255.020 52.480 ;
        RECT 244.455 52.455 245.195 52.470 ;
        RECT 243.350 52.365 243.765 52.455 ;
        POLYGON 243.300 52.365 243.300 52.270 243.270 52.270 ;
        RECT 243.300 52.270 243.765 52.365 ;
        RECT 241.825 52.245 242.615 52.270 ;
        POLYGON 242.615 52.270 242.625 52.270 242.615 52.245 ;
        POLYGON 243.270 52.265 243.270 52.250 243.265 52.250 ;
        RECT 243.270 52.250 243.765 52.270 ;
        POLYGON 241.790 52.245 241.790 52.110 241.755 52.110 ;
        RECT 241.790 52.195 242.605 52.245 ;
        POLYGON 242.605 52.245 242.615 52.245 242.605 52.195 ;
        POLYGON 243.265 52.245 243.265 52.200 243.250 52.200 ;
        RECT 243.265 52.235 243.765 52.250 ;
        POLYGON 243.765 52.455 243.850 52.455 243.765 52.235 ;
        POLYGON 244.430 52.450 244.430 52.400 244.410 52.400 ;
        RECT 244.430 52.400 245.195 52.455 ;
        POLYGON 244.410 52.400 244.410 52.330 244.385 52.330 ;
        RECT 244.410 52.330 245.195 52.400 ;
        POLYGON 244.385 52.325 244.385 52.235 244.355 52.235 ;
        RECT 244.385 52.310 245.195 52.330 ;
        POLYGON 245.195 52.470 245.280 52.470 245.195 52.310 ;
        POLYGON 254.320 52.470 254.405 52.470 254.405 52.335 ;
        RECT 254.405 52.385 255.020 52.470 ;
        POLYGON 255.020 52.510 255.085 52.385 255.020 52.385 ;
        POLYGON 255.555 52.510 255.580 52.510 255.580 52.455 ;
        RECT 255.580 52.455 255.960 52.510 ;
        POLYGON 255.580 52.455 255.590 52.455 255.590 52.435 ;
        RECT 255.590 52.435 255.960 52.455 ;
        POLYGON 255.590 52.435 255.605 52.435 255.605 52.390 ;
        RECT 255.605 52.415 255.960 52.435 ;
        POLYGON 255.960 52.575 256.035 52.415 255.960 52.415 ;
        RECT 256.565 52.565 257.180 52.590 ;
        POLYGON 256.565 52.565 256.585 52.565 256.585 52.525 ;
        RECT 256.585 52.525 257.180 52.565 ;
        POLYGON 257.180 52.590 257.205 52.525 257.180 52.525 ;
        POLYGON 257.995 52.590 258.020 52.590 258.020 52.530 ;
        RECT 258.020 52.525 258.940 52.590 ;
        RECT 256.585 52.520 257.205 52.525 ;
        POLYGON 256.585 52.520 256.590 52.520 256.590 52.505 ;
        RECT 256.590 52.505 257.205 52.520 ;
        POLYGON 256.590 52.505 256.625 52.505 256.625 52.415 ;
        RECT 256.625 52.435 257.205 52.505 ;
        POLYGON 257.205 52.525 257.235 52.435 257.205 52.435 ;
        POLYGON 258.020 52.525 258.050 52.525 258.050 52.445 ;
        RECT 258.050 52.435 258.940 52.525 ;
        RECT 256.625 52.415 257.235 52.435 ;
        RECT 255.605 52.385 256.035 52.415 ;
        RECT 254.405 52.370 255.085 52.385 ;
        POLYGON 255.085 52.385 255.090 52.370 255.085 52.370 ;
        POLYGON 255.605 52.385 255.610 52.385 255.610 52.380 ;
        RECT 255.610 52.370 256.035 52.385 ;
        RECT 254.405 52.335 255.090 52.370 ;
        POLYGON 254.405 52.335 254.415 52.335 254.415 52.315 ;
        RECT 254.415 52.310 255.090 52.335 ;
        RECT 244.385 52.300 245.190 52.310 ;
        POLYGON 245.190 52.310 245.195 52.310 245.190 52.300 ;
        POLYGON 254.415 52.310 254.420 52.310 254.420 52.305 ;
        RECT 254.420 52.300 255.090 52.310 ;
        RECT 244.385 52.285 245.180 52.300 ;
        POLYGON 245.180 52.300 245.190 52.300 245.180 52.285 ;
        POLYGON 254.420 52.300 254.430 52.300 254.430 52.290 ;
        RECT 254.430 52.285 255.090 52.300 ;
        RECT 244.385 52.255 245.165 52.285 ;
        POLYGON 245.165 52.285 245.180 52.285 245.165 52.255 ;
        POLYGON 254.430 52.285 254.450 52.285 254.450 52.255 ;
        RECT 254.450 52.255 255.090 52.285 ;
        RECT 244.385 52.235 245.115 52.255 ;
        RECT 243.265 52.220 243.760 52.235 ;
        POLYGON 243.760 52.235 243.765 52.235 243.760 52.220 ;
        POLYGON 244.355 52.235 244.355 52.220 244.350 52.220 ;
        RECT 244.355 52.220 245.115 52.235 ;
        RECT 243.265 52.210 243.755 52.220 ;
        POLYGON 243.755 52.220 243.760 52.220 243.755 52.210 ;
        RECT 243.265 52.200 243.735 52.210 ;
        RECT 241.790 52.110 242.550 52.195 ;
        RECT 239.730 52.030 240.755 52.110 ;
        POLYGON 239.690 52.030 239.690 51.930 239.675 51.930 ;
        RECT 239.690 51.990 240.755 52.030 ;
        POLYGON 240.755 52.110 240.775 52.110 240.755 52.000 ;
        POLYGON 241.755 52.105 241.755 52.000 241.730 52.000 ;
        RECT 241.755 52.000 242.550 52.110 ;
        RECT 239.690 51.930 240.735 51.990 ;
        RECT 236.040 51.865 238.020 51.915 ;
        POLYGON 229.190 51.355 229.205 51.355 229.205 50.965 ;
        RECT 229.205 50.965 233.200 51.865 ;
        POLYGON 233.200 51.865 233.220 51.865 233.200 51.175 ;
        POLYGON 236.020 51.840 236.020 51.645 236.005 51.645 ;
        RECT 236.020 51.765 238.020 51.865 ;
        POLYGON 238.020 51.915 238.035 51.915 238.020 51.765 ;
        POLYGON 239.675 51.915 239.675 51.800 239.655 51.800 ;
        RECT 239.675 51.865 240.735 51.930 ;
        POLYGON 240.735 51.990 240.755 51.990 240.735 51.865 ;
        POLYGON 241.730 52.000 241.730 51.920 241.710 51.920 ;
        RECT 241.730 51.970 242.550 52.000 ;
        POLYGON 242.550 52.195 242.605 52.195 242.550 51.980 ;
        POLYGON 243.250 52.195 243.250 52.150 243.235 52.150 ;
        RECT 243.250 52.150 243.735 52.200 ;
        POLYGON 243.735 52.210 243.755 52.210 243.735 52.150 ;
        POLYGON 244.350 52.210 244.350 52.155 244.330 52.155 ;
        RECT 244.350 52.155 245.115 52.220 ;
        RECT 244.330 52.150 245.115 52.155 ;
        POLYGON 245.115 52.255 245.165 52.255 245.115 52.150 ;
        POLYGON 254.450 52.255 254.490 52.255 254.490 52.185 ;
        RECT 254.490 52.220 255.090 52.255 ;
        POLYGON 255.090 52.370 255.160 52.220 255.090 52.220 ;
        POLYGON 255.610 52.370 255.615 52.370 255.615 52.365 ;
        RECT 255.615 52.365 256.035 52.370 ;
        POLYGON 255.615 52.365 255.635 52.365 255.635 52.325 ;
        RECT 255.635 52.350 256.035 52.365 ;
        POLYGON 256.035 52.415 256.065 52.350 256.035 52.350 ;
        POLYGON 256.625 52.415 256.650 52.415 256.650 52.350 ;
        RECT 256.650 52.350 257.235 52.415 ;
        RECT 255.635 52.320 256.065 52.350 ;
        POLYGON 255.635 52.320 255.640 52.320 255.640 52.310 ;
        RECT 255.640 52.315 256.065 52.320 ;
        POLYGON 256.065 52.350 256.080 52.315 256.065 52.315 ;
        POLYGON 256.650 52.350 256.665 52.350 256.665 52.315 ;
        RECT 255.640 52.310 256.080 52.315 ;
        RECT 256.665 52.310 257.235 52.350 ;
        POLYGON 255.640 52.310 255.655 52.310 255.655 52.270 ;
        RECT 255.655 52.265 256.080 52.310 ;
        POLYGON 255.655 52.265 255.665 52.265 255.665 52.235 ;
        RECT 255.665 52.235 256.080 52.265 ;
        POLYGON 255.665 52.235 255.670 52.235 255.670 52.230 ;
        RECT 255.670 52.220 256.080 52.235 ;
        RECT 254.490 52.190 255.160 52.220 ;
        POLYGON 255.160 52.220 255.175 52.190 255.160 52.190 ;
        POLYGON 255.670 52.220 255.675 52.220 255.675 52.215 ;
        RECT 255.675 52.215 256.080 52.220 ;
        POLYGON 255.675 52.215 255.680 52.215 255.680 52.205 ;
        RECT 255.680 52.190 256.080 52.215 ;
        RECT 254.490 52.185 255.175 52.190 ;
        POLYGON 254.490 52.185 254.505 52.185 254.505 52.155 ;
        RECT 254.505 52.150 255.175 52.185 ;
        POLYGON 243.235 52.150 243.235 52.140 243.230 52.140 ;
        RECT 243.235 52.140 243.675 52.150 ;
        POLYGON 243.230 52.140 243.230 52.105 243.220 52.105 ;
        RECT 243.230 52.105 243.675 52.140 ;
        POLYGON 243.220 52.105 243.220 51.990 243.190 51.990 ;
        RECT 243.220 51.990 243.675 52.105 ;
        RECT 241.730 51.920 242.525 51.970 ;
        POLYGON 241.710 51.920 241.710 51.870 241.700 51.870 ;
        RECT 241.710 51.870 242.525 51.920 ;
        RECT 239.675 51.800 240.700 51.865 ;
        POLYGON 239.655 51.800 239.655 51.765 239.650 51.765 ;
        RECT 239.655 51.765 240.700 51.800 ;
        RECT 236.020 51.645 237.985 51.765 ;
        POLYGON 236.005 51.645 236.005 51.390 235.985 51.390 ;
        RECT 236.005 51.390 237.985 51.645 ;
        POLYGON 229.205 50.965 229.225 50.965 229.225 50.525 ;
        RECT 229.225 50.495 233.200 50.965 ;
        RECT 207.110 49.245 222.255 50.495 ;
        POLYGON 197.510 49.245 197.580 48.835 197.510 48.835 ;
        POLYGON 207.110 49.245 207.185 49.245 207.185 48.850 ;
        RECT 207.185 48.835 222.255 49.245 ;
        RECT 182.900 48.720 197.580 48.835 ;
        POLYGON 197.580 48.835 197.600 48.720 197.580 48.720 ;
        POLYGON 207.185 48.835 207.210 48.835 207.210 48.720 ;
        RECT 207.210 48.720 222.255 48.835 ;
        RECT 182.900 48.705 197.600 48.720 ;
        POLYGON 171.730 48.140 171.730 48.075 171.725 48.075 ;
        RECT 171.730 48.075 175.685 48.140 ;
        POLYGON 171.725 48.075 171.725 47.860 171.710 47.860 ;
        RECT 171.725 47.860 175.685 48.075 ;
        RECT 166.950 47.830 168.965 47.860 ;
        RECT 164.195 47.680 165.300 47.780 ;
        POLYGON 164.155 47.675 164.155 47.595 164.135 47.595 ;
        RECT 164.155 47.595 165.300 47.680 ;
        RECT 162.390 47.585 163.145 47.595 ;
        POLYGON 162.380 47.585 162.380 47.525 162.365 47.525 ;
        RECT 162.380 47.525 163.145 47.585 ;
        POLYGON 162.365 47.525 162.365 47.385 162.320 47.385 ;
        RECT 162.365 47.385 163.145 47.525 ;
        RECT 160.095 47.325 160.555 47.375 ;
        POLYGON 160.055 47.325 160.055 47.300 160.045 47.300 ;
        RECT 160.055 47.310 160.555 47.325 ;
        POLYGON 160.555 47.375 160.585 47.375 160.555 47.310 ;
        POLYGON 161.075 47.375 161.075 47.335 161.060 47.335 ;
        RECT 161.075 47.335 161.620 47.380 ;
        POLYGON 161.060 47.335 161.060 47.315 161.050 47.315 ;
        RECT 161.060 47.315 161.620 47.335 ;
        RECT 160.055 47.300 160.535 47.310 ;
        POLYGON 160.045 47.300 160.045 47.240 160.010 47.240 ;
        RECT 160.045 47.260 160.535 47.300 ;
        POLYGON 160.535 47.310 160.555 47.310 160.535 47.260 ;
        POLYGON 161.050 47.310 161.050 47.295 161.040 47.295 ;
        RECT 161.050 47.295 161.620 47.315 ;
        POLYGON 161.040 47.295 161.040 47.265 161.025 47.265 ;
        RECT 161.040 47.265 161.620 47.295 ;
        RECT 160.045 47.240 160.475 47.260 ;
        POLYGON 160.010 47.235 160.010 47.230 160.005 47.230 ;
        RECT 160.010 47.230 160.475 47.240 ;
        RECT 150.550 47.220 159.065 47.230 ;
        RECT 117.220 47.205 149.685 47.220 ;
        POLYGON 149.685 47.220 149.690 47.205 149.685 47.205 ;
        POLYGON 150.550 47.220 150.555 47.220 150.555 47.210 ;
        RECT 150.555 47.205 159.065 47.220 ;
        RECT 117.220 47.185 149.690 47.205 ;
        POLYGON 149.690 47.205 149.705 47.185 149.690 47.185 ;
        RECT 117.220 47.155 149.705 47.185 ;
        POLYGON 150.555 47.205 150.575 47.205 150.575 47.180 ;
        RECT 150.575 47.180 159.065 47.205 ;
        POLYGON 149.705 47.180 149.720 47.155 149.705 47.155 ;
        POLYGON 150.575 47.180 150.590 47.180 150.590 47.155 ;
        RECT 150.590 47.155 159.065 47.180 ;
        RECT 117.220 47.140 149.720 47.155 ;
        POLYGON 117.220 47.140 117.235 47.140 117.235 46.535 ;
        RECT 117.235 47.135 149.720 47.140 ;
        POLYGON 149.720 47.155 149.730 47.135 149.720 47.135 ;
        POLYGON 150.590 47.155 150.605 47.155 150.605 47.135 ;
        RECT 150.605 47.135 159.065 47.155 ;
        POLYGON 159.065 47.230 159.130 47.230 159.065 47.135 ;
        POLYGON 160.005 47.230 160.005 47.215 159.995 47.215 ;
        RECT 160.005 47.215 160.475 47.230 ;
        POLYGON 159.995 47.210 159.995 47.195 159.985 47.195 ;
        RECT 159.995 47.195 160.475 47.215 ;
        POLYGON 159.985 47.195 159.985 47.170 159.975 47.170 ;
        RECT 159.985 47.170 160.475 47.195 ;
        POLYGON 159.975 47.170 159.975 47.135 159.955 47.135 ;
        RECT 159.975 47.135 160.475 47.170 ;
        RECT 117.235 47.090 149.730 47.135 ;
        POLYGON 149.730 47.135 149.755 47.090 149.730 47.090 ;
        POLYGON 150.605 47.135 150.635 47.135 150.635 47.090 ;
        RECT 150.635 47.130 159.060 47.135 ;
        POLYGON 159.060 47.135 159.065 47.135 159.060 47.130 ;
        RECT 159.955 47.130 160.475 47.135 ;
        POLYGON 160.475 47.260 160.535 47.260 160.475 47.130 ;
        POLYGON 161.025 47.260 161.025 47.160 160.975 47.160 ;
        RECT 161.025 47.230 161.620 47.265 ;
        POLYGON 161.620 47.380 161.675 47.380 161.620 47.230 ;
        POLYGON 162.320 47.380 162.320 47.305 162.295 47.305 ;
        RECT 162.320 47.305 163.145 47.385 ;
        POLYGON 162.295 47.305 162.295 47.230 162.265 47.230 ;
        RECT 162.295 47.230 163.145 47.305 ;
        RECT 161.025 47.160 161.570 47.230 ;
        POLYGON 160.975 47.150 160.975 47.135 160.965 47.135 ;
        RECT 160.975 47.135 161.570 47.160 ;
        RECT 150.635 47.090 158.950 47.130 ;
        RECT 117.235 47.075 149.755 47.090 ;
        POLYGON 149.755 47.090 149.765 47.075 149.755 47.075 ;
        POLYGON 150.635 47.090 150.645 47.090 150.645 47.075 ;
        RECT 150.645 47.075 158.950 47.090 ;
        RECT 117.235 47.010 149.765 47.075 ;
        POLYGON 149.765 47.075 149.800 47.010 149.765 47.010 ;
        POLYGON 150.645 47.075 150.655 47.075 150.655 47.060 ;
        RECT 150.655 47.060 158.950 47.075 ;
        POLYGON 150.655 47.060 150.690 47.060 150.690 47.010 ;
        RECT 150.690 47.010 158.950 47.060 ;
        RECT 117.235 47.000 149.800 47.010 ;
        POLYGON 149.800 47.010 149.805 47.000 149.800 47.000 ;
        POLYGON 150.690 47.010 150.695 47.010 150.695 47.005 ;
        RECT 150.695 47.000 158.950 47.010 ;
        RECT 117.235 46.935 149.805 47.000 ;
        POLYGON 149.805 47.000 149.840 46.935 149.805 46.935 ;
        POLYGON 150.695 47.000 150.735 47.000 150.735 46.955 ;
        RECT 150.735 46.995 158.950 47.000 ;
        POLYGON 158.950 47.130 159.060 47.130 158.950 46.995 ;
        POLYGON 159.955 47.130 159.955 47.125 159.950 47.125 ;
        RECT 159.955 47.125 160.400 47.130 ;
        POLYGON 159.950 47.125 159.950 47.050 159.900 47.050 ;
        RECT 159.950 47.050 160.400 47.125 ;
        POLYGON 159.900 47.050 159.900 47.000 159.875 47.000 ;
        RECT 159.900 47.000 160.400 47.050 ;
        RECT 150.735 46.955 158.855 46.995 ;
        POLYGON 150.735 46.955 150.745 46.955 150.745 46.940 ;
        RECT 150.745 46.935 158.855 46.955 ;
        RECT 117.235 46.920 149.840 46.935 ;
        POLYGON 149.840 46.935 149.850 46.920 149.840 46.920 ;
        POLYGON 150.745 46.935 150.755 46.935 150.755 46.925 ;
        RECT 150.755 46.920 158.855 46.935 ;
        RECT 117.235 46.915 149.850 46.920 ;
        POLYGON 149.850 46.920 149.855 46.915 149.850 46.915 ;
        RECT 117.235 46.830 149.855 46.915 ;
        POLYGON 150.755 46.920 150.765 46.920 150.765 46.910 ;
        RECT 150.765 46.910 158.855 46.920 ;
        POLYGON 149.855 46.910 149.905 46.830 149.855 46.830 ;
        POLYGON 150.765 46.910 150.825 46.910 150.825 46.830 ;
        RECT 150.825 46.875 158.855 46.910 ;
        POLYGON 158.855 46.995 158.950 46.995 158.855 46.875 ;
        POLYGON 159.875 46.995 159.875 46.990 159.870 46.990 ;
        RECT 159.875 46.990 160.400 47.000 ;
        POLYGON 159.870 46.990 159.870 46.930 159.830 46.930 ;
        RECT 159.870 46.985 160.400 46.990 ;
        POLYGON 160.400 47.130 160.475 47.130 160.400 46.985 ;
        POLYGON 160.965 47.130 160.965 47.115 160.955 47.115 ;
        RECT 160.965 47.115 161.570 47.135 ;
        POLYGON 160.955 47.115 160.955 47.070 160.935 47.070 ;
        RECT 160.955 47.110 161.570 47.115 ;
        POLYGON 161.570 47.230 161.620 47.230 161.570 47.110 ;
        POLYGON 162.265 47.225 162.265 47.110 162.220 47.110 ;
        RECT 162.265 47.175 163.145 47.230 ;
        POLYGON 163.145 47.595 163.270 47.595 163.145 47.175 ;
        POLYGON 164.135 47.585 164.135 47.430 164.100 47.430 ;
        RECT 164.135 47.430 165.300 47.595 ;
        POLYGON 164.100 47.430 164.100 47.240 164.050 47.240 ;
        RECT 164.100 47.240 165.300 47.430 ;
        POLYGON 164.050 47.240 164.050 47.180 164.035 47.180 ;
        RECT 164.050 47.235 165.300 47.240 ;
        POLYGON 165.300 47.780 165.385 47.780 165.300 47.235 ;
        POLYGON 166.930 47.780 166.930 47.520 166.910 47.520 ;
        RECT 166.930 47.520 168.965 47.830 ;
        POLYGON 166.910 47.520 166.910 47.235 166.880 47.235 ;
        RECT 166.910 47.365 168.965 47.520 ;
        POLYGON 168.965 47.860 169.020 47.860 168.965 47.365 ;
        POLYGON 171.710 47.825 171.710 47.405 171.685 47.405 ;
        RECT 171.710 47.405 175.685 47.860 ;
        POLYGON 171.685 47.405 171.685 47.365 171.680 47.365 ;
        RECT 171.685 47.365 175.685 47.405 ;
        RECT 166.910 47.235 168.890 47.365 ;
        RECT 164.050 47.180 165.190 47.235 ;
        RECT 162.265 47.125 163.125 47.175 ;
        POLYGON 163.125 47.175 163.145 47.175 163.125 47.125 ;
        POLYGON 164.035 47.175 164.035 47.125 164.020 47.125 ;
        RECT 164.035 47.125 165.190 47.180 ;
        RECT 162.265 47.110 163.120 47.125 ;
        RECT 160.955 47.075 161.555 47.110 ;
        POLYGON 161.555 47.110 161.570 47.110 161.555 47.075 ;
        RECT 162.220 47.105 163.120 47.110 ;
        POLYGON 163.120 47.125 163.125 47.125 163.120 47.105 ;
        POLYGON 164.020 47.125 164.020 47.105 164.015 47.105 ;
        RECT 164.020 47.105 165.190 47.125 ;
        POLYGON 162.220 47.105 162.220 47.080 162.210 47.080 ;
        RECT 162.220 47.080 162.995 47.105 ;
        RECT 160.955 47.070 161.455 47.075 ;
        POLYGON 160.935 47.070 160.935 47.045 160.925 47.045 ;
        RECT 160.935 47.045 161.455 47.070 ;
        POLYGON 160.925 47.045 160.925 46.985 160.890 46.985 ;
        RECT 160.925 46.985 161.455 47.045 ;
        RECT 159.870 46.950 160.385 46.985 ;
        POLYGON 160.385 46.985 160.400 46.985 160.385 46.950 ;
        POLYGON 160.890 46.985 160.890 46.965 160.880 46.965 ;
        RECT 160.890 46.965 161.455 46.985 ;
        POLYGON 160.880 46.965 160.880 46.960 160.875 46.960 ;
        RECT 160.880 46.960 161.455 46.965 ;
        POLYGON 160.875 46.960 160.875 46.950 160.870 46.950 ;
        RECT 160.875 46.950 161.455 46.960 ;
        RECT 159.870 46.930 160.345 46.950 ;
        POLYGON 159.830 46.925 159.830 46.875 159.795 46.875 ;
        RECT 159.830 46.880 160.345 46.930 ;
        POLYGON 160.345 46.950 160.385 46.950 160.345 46.880 ;
        POLYGON 160.870 46.950 160.870 46.880 160.835 46.880 ;
        RECT 160.870 46.880 161.455 46.950 ;
        RECT 159.830 46.875 160.280 46.880 ;
        RECT 150.825 46.830 158.790 46.875 ;
        RECT 117.235 46.805 149.905 46.830 ;
        POLYGON 149.905 46.830 149.920 46.805 149.905 46.805 ;
        POLYGON 150.825 46.830 150.845 46.830 150.845 46.805 ;
        RECT 150.845 46.805 158.790 46.830 ;
        RECT 117.235 46.790 149.920 46.805 ;
        POLYGON 149.920 46.805 149.930 46.790 149.920 46.790 ;
        POLYGON 150.845 46.805 150.855 46.805 150.855 46.790 ;
        RECT 150.855 46.800 158.790 46.805 ;
        POLYGON 158.790 46.875 158.855 46.875 158.790 46.800 ;
        POLYGON 159.795 46.875 159.795 46.860 159.785 46.860 ;
        RECT 159.795 46.860 160.280 46.875 ;
        POLYGON 159.785 46.860 159.785 46.835 159.770 46.835 ;
        RECT 159.785 46.835 160.280 46.860 ;
        POLYGON 159.770 46.835 159.770 46.800 159.745 46.800 ;
        RECT 159.770 46.800 160.280 46.835 ;
        RECT 150.855 46.790 158.630 46.800 ;
        RECT 117.235 46.735 149.930 46.790 ;
        POLYGON 149.930 46.790 149.965 46.735 149.930 46.735 ;
        POLYGON 150.855 46.790 150.870 46.790 150.870 46.775 ;
        RECT 150.870 46.775 158.630 46.790 ;
        POLYGON 150.870 46.775 150.880 46.775 150.880 46.760 ;
        RECT 150.880 46.760 158.630 46.775 ;
        POLYGON 150.880 46.760 150.900 46.760 150.900 46.735 ;
        RECT 150.900 46.735 158.630 46.760 ;
        RECT 117.235 46.695 149.965 46.735 ;
        POLYGON 149.965 46.735 149.990 46.695 149.965 46.695 ;
        POLYGON 150.900 46.735 150.935 46.735 150.935 46.695 ;
        RECT 150.935 46.695 158.630 46.735 ;
        RECT 117.235 46.690 149.990 46.695 ;
        POLYGON 149.990 46.695 149.995 46.690 149.990 46.690 ;
        POLYGON 150.935 46.695 150.940 46.695 150.940 46.690 ;
        RECT 150.940 46.690 158.630 46.695 ;
        RECT 117.235 46.665 149.995 46.690 ;
        POLYGON 149.995 46.690 150.010 46.665 149.995 46.665 ;
        POLYGON 150.940 46.690 150.960 46.690 150.960 46.665 ;
        RECT 150.960 46.665 158.630 46.690 ;
        RECT 117.235 46.635 150.010 46.665 ;
        POLYGON 150.010 46.665 150.030 46.635 150.010 46.635 ;
        POLYGON 150.960 46.665 150.985 46.665 150.985 46.635 ;
        RECT 150.985 46.635 158.630 46.665 ;
        RECT 117.235 46.570 150.030 46.635 ;
        POLYGON 150.030 46.635 150.075 46.570 150.030 46.570 ;
        POLYGON 150.985 46.635 151.000 46.635 151.000 46.620 ;
        RECT 151.000 46.620 158.630 46.635 ;
        POLYGON 158.630 46.800 158.790 46.800 158.630 46.620 ;
        POLYGON 159.745 46.800 159.745 46.785 159.735 46.785 ;
        RECT 159.745 46.785 160.280 46.800 ;
        POLYGON 159.735 46.785 159.735 46.735 159.705 46.735 ;
        RECT 159.735 46.775 160.280 46.785 ;
        POLYGON 160.280 46.880 160.345 46.880 160.280 46.775 ;
        POLYGON 160.835 46.875 160.835 46.845 160.820 46.845 ;
        RECT 160.835 46.845 161.455 46.880 ;
        POLYGON 160.820 46.845 160.820 46.775 160.780 46.775 ;
        RECT 160.820 46.840 161.455 46.845 ;
        POLYGON 161.455 47.075 161.555 47.075 161.455 46.840 ;
        POLYGON 162.210 47.075 162.210 47.000 162.180 47.000 ;
        RECT 162.210 47.000 162.995 47.080 ;
        POLYGON 162.180 47.000 162.180 46.970 162.170 46.970 ;
        RECT 162.180 46.970 162.995 47.000 ;
        POLYGON 162.170 46.970 162.170 46.840 162.115 46.840 ;
        RECT 162.170 46.840 162.995 46.970 ;
        RECT 160.820 46.775 161.325 46.840 ;
        RECT 159.735 46.735 160.205 46.775 ;
        POLYGON 159.705 46.735 159.705 46.705 159.680 46.705 ;
        RECT 159.705 46.705 160.205 46.735 ;
        POLYGON 159.680 46.705 159.680 46.620 159.625 46.620 ;
        RECT 159.680 46.660 160.205 46.705 ;
        POLYGON 160.205 46.775 160.280 46.775 160.205 46.660 ;
        POLYGON 160.780 46.775 160.780 46.735 160.760 46.735 ;
        RECT 160.780 46.735 161.325 46.775 ;
        POLYGON 160.760 46.735 160.760 46.715 160.745 46.715 ;
        RECT 160.760 46.715 161.325 46.735 ;
        POLYGON 160.745 46.715 160.745 46.665 160.715 46.665 ;
        RECT 160.745 46.665 161.325 46.715 ;
        RECT 159.680 46.620 160.165 46.660 ;
        POLYGON 151.000 46.620 151.010 46.620 151.010 46.605 ;
        RECT 151.010 46.605 158.580 46.620 ;
        POLYGON 151.010 46.605 151.045 46.605 151.045 46.570 ;
        RECT 151.045 46.575 158.580 46.605 ;
        POLYGON 158.580 46.620 158.630 46.620 158.580 46.575 ;
        POLYGON 159.620 46.620 159.620 46.575 159.590 46.575 ;
        RECT 159.620 46.595 160.165 46.620 ;
        POLYGON 160.165 46.660 160.205 46.660 160.165 46.595 ;
        POLYGON 160.715 46.660 160.715 46.655 160.710 46.655 ;
        RECT 160.715 46.655 161.325 46.665 ;
        POLYGON 160.710 46.655 160.710 46.640 160.705 46.640 ;
        RECT 160.710 46.640 161.325 46.655 ;
        POLYGON 160.705 46.640 160.705 46.595 160.680 46.595 ;
        RECT 160.705 46.595 161.325 46.640 ;
        RECT 159.620 46.575 160.145 46.595 ;
        RECT 151.045 46.570 158.380 46.575 ;
        RECT 117.235 46.530 150.075 46.570 ;
        POLYGON 150.075 46.570 150.105 46.530 150.075 46.530 ;
        POLYGON 151.045 46.570 151.075 46.570 151.075 46.540 ;
        RECT 151.075 46.540 158.380 46.570 ;
        POLYGON 151.075 46.540 151.080 46.540 151.080 46.530 ;
        RECT 151.080 46.530 158.380 46.540 ;
        RECT 117.235 46.460 150.105 46.530 ;
        POLYGON 150.105 46.530 150.150 46.460 150.105 46.460 ;
        POLYGON 151.080 46.530 151.125 46.530 151.125 46.480 ;
        RECT 151.125 46.480 158.380 46.530 ;
        POLYGON 151.125 46.480 151.145 46.480 151.145 46.460 ;
        RECT 151.145 46.460 158.380 46.480 ;
        RECT 117.235 46.445 150.150 46.460 ;
        POLYGON 150.150 46.460 150.165 46.445 150.150 46.445 ;
        POLYGON 151.145 46.460 151.160 46.460 151.160 46.445 ;
        RECT 151.160 46.445 158.380 46.460 ;
        RECT 117.235 46.425 150.165 46.445 ;
        POLYGON 150.165 46.445 150.180 46.425 150.165 46.425 ;
        POLYGON 151.160 46.445 151.175 46.445 151.175 46.425 ;
        RECT 151.175 46.425 158.380 46.445 ;
        RECT 117.235 46.415 150.180 46.425 ;
        POLYGON 117.235 46.415 117.245 46.415 117.245 46.005 ;
        RECT 117.245 46.315 150.180 46.415 ;
        POLYGON 150.180 46.425 150.265 46.315 150.180 46.315 ;
        POLYGON 151.175 46.425 151.285 46.425 151.285 46.315 ;
        RECT 151.285 46.375 158.380 46.425 ;
        POLYGON 158.380 46.575 158.580 46.575 158.380 46.375 ;
        POLYGON 159.590 46.575 159.590 46.545 159.570 46.545 ;
        RECT 159.590 46.565 160.145 46.575 ;
        POLYGON 160.145 46.595 160.165 46.595 160.145 46.565 ;
        POLYGON 160.680 46.595 160.680 46.570 160.665 46.570 ;
        RECT 160.680 46.575 161.325 46.595 ;
        POLYGON 161.325 46.840 161.455 46.840 161.325 46.575 ;
        POLYGON 162.115 46.840 162.115 46.800 162.100 46.800 ;
        RECT 162.115 46.800 162.995 46.840 ;
        POLYGON 162.100 46.800 162.100 46.775 162.090 46.775 ;
        RECT 162.100 46.775 162.995 46.800 ;
        POLYGON 162.090 46.775 162.090 46.720 162.065 46.720 ;
        RECT 162.090 46.765 162.995 46.775 ;
        POLYGON 162.995 47.105 163.120 47.105 162.995 46.765 ;
        POLYGON 164.015 47.105 164.015 47.085 164.010 47.085 ;
        RECT 164.015 47.085 165.190 47.105 ;
        POLYGON 164.010 47.085 164.010 47.000 163.985 47.000 ;
        RECT 164.010 47.000 165.190 47.085 ;
        POLYGON 163.985 47.000 163.985 46.790 163.915 46.790 ;
        RECT 163.985 46.790 165.190 47.000 ;
        POLYGON 163.915 46.790 163.915 46.765 163.905 46.765 ;
        RECT 163.915 46.765 165.190 46.790 ;
        RECT 162.090 46.720 162.825 46.765 ;
        POLYGON 162.065 46.720 162.065 46.695 162.055 46.695 ;
        RECT 162.065 46.695 162.825 46.720 ;
        POLYGON 162.055 46.695 162.055 46.640 162.030 46.640 ;
        RECT 162.055 46.640 162.825 46.695 ;
        POLYGON 162.030 46.640 162.030 46.575 162.000 46.575 ;
        RECT 162.030 46.575 162.825 46.640 ;
        RECT 160.680 46.570 161.305 46.575 ;
        RECT 159.590 46.545 160.045 46.565 ;
        POLYGON 159.570 46.545 159.570 46.540 159.565 46.540 ;
        RECT 159.570 46.540 160.045 46.545 ;
        POLYGON 159.565 46.540 159.565 46.530 159.560 46.530 ;
        RECT 159.565 46.530 160.045 46.540 ;
        POLYGON 159.560 46.530 159.560 46.440 159.490 46.440 ;
        RECT 159.560 46.440 160.045 46.530 ;
        POLYGON 159.490 46.440 159.490 46.410 159.465 46.410 ;
        RECT 159.490 46.420 160.045 46.440 ;
        POLYGON 160.045 46.565 160.145 46.565 160.045 46.420 ;
        POLYGON 160.665 46.565 160.665 46.550 160.650 46.550 ;
        RECT 160.665 46.550 161.305 46.570 ;
        POLYGON 160.650 46.550 160.650 46.485 160.610 46.485 ;
        RECT 160.650 46.540 161.305 46.550 ;
        POLYGON 161.305 46.575 161.325 46.575 161.305 46.540 ;
        POLYGON 162.000 46.575 162.000 46.540 161.985 46.540 ;
        RECT 162.000 46.540 162.825 46.575 ;
        RECT 160.650 46.485 161.240 46.540 ;
        POLYGON 160.610 46.485 160.610 46.445 160.585 46.445 ;
        RECT 160.610 46.445 161.240 46.485 ;
        POLYGON 160.585 46.445 160.585 46.420 160.565 46.420 ;
        RECT 160.585 46.420 161.240 46.445 ;
        RECT 159.490 46.410 160.005 46.420 ;
        POLYGON 159.465 46.410 159.465 46.375 159.435 46.375 ;
        RECT 159.465 46.375 160.005 46.410 ;
        RECT 151.285 46.315 158.230 46.375 ;
        RECT 117.245 46.240 150.265 46.315 ;
        POLYGON 150.265 46.315 150.325 46.240 150.265 46.240 ;
        POLYGON 151.285 46.315 151.315 46.315 151.315 46.290 ;
        RECT 151.315 46.290 158.230 46.315 ;
        POLYGON 151.315 46.290 151.365 46.290 151.365 46.240 ;
        RECT 151.365 46.240 158.230 46.290 ;
        RECT 117.245 46.220 150.325 46.240 ;
        POLYGON 150.325 46.240 150.340 46.220 150.325 46.220 ;
        POLYGON 151.365 46.240 151.385 46.240 151.385 46.220 ;
        RECT 151.385 46.235 158.230 46.240 ;
        POLYGON 158.230 46.375 158.380 46.375 158.230 46.235 ;
        POLYGON 159.435 46.375 159.435 46.345 159.415 46.345 ;
        RECT 159.435 46.370 160.005 46.375 ;
        POLYGON 160.005 46.420 160.045 46.420 160.005 46.370 ;
        POLYGON 160.565 46.420 160.565 46.405 160.555 46.405 ;
        RECT 160.565 46.415 161.240 46.420 ;
        POLYGON 161.240 46.540 161.305 46.540 161.240 46.415 ;
        POLYGON 161.985 46.540 161.985 46.415 161.925 46.415 ;
        RECT 161.985 46.415 162.825 46.540 ;
        RECT 160.565 46.405 161.190 46.415 ;
        POLYGON 160.555 46.405 160.555 46.375 160.540 46.375 ;
        RECT 160.555 46.375 161.190 46.405 ;
        RECT 159.435 46.345 159.940 46.370 ;
        POLYGON 159.415 46.345 159.415 46.250 159.335 46.250 ;
        RECT 159.415 46.280 159.940 46.345 ;
        POLYGON 159.940 46.370 160.005 46.370 159.940 46.280 ;
        POLYGON 160.540 46.370 160.540 46.365 160.535 46.365 ;
        RECT 160.540 46.365 161.190 46.375 ;
        POLYGON 160.535 46.365 160.535 46.295 160.490 46.295 ;
        RECT 160.535 46.320 161.190 46.365 ;
        POLYGON 161.190 46.415 161.240 46.415 161.190 46.320 ;
        POLYGON 161.925 46.410 161.925 46.390 161.915 46.390 ;
        RECT 161.925 46.390 162.825 46.415 ;
        POLYGON 161.915 46.390 161.915 46.375 161.905 46.375 ;
        RECT 161.915 46.375 162.825 46.390 ;
        POLYGON 161.905 46.375 161.905 46.325 161.880 46.325 ;
        RECT 161.905 46.355 162.825 46.375 ;
        POLYGON 162.825 46.765 162.995 46.765 162.825 46.360 ;
        POLYGON 163.905 46.760 163.905 46.575 163.845 46.575 ;
        RECT 163.905 46.710 165.190 46.765 ;
        POLYGON 165.190 47.235 165.300 47.235 165.190 46.710 ;
        POLYGON 166.880 47.230 166.880 47.030 166.850 47.030 ;
        RECT 166.880 47.030 168.890 47.235 ;
        POLYGON 166.850 47.030 166.850 46.960 166.840 46.960 ;
        RECT 166.850 46.960 168.890 47.030 ;
        POLYGON 166.840 46.960 166.840 46.860 166.825 46.860 ;
        RECT 166.840 46.870 168.890 46.960 ;
        POLYGON 168.890 47.365 168.965 47.365 168.890 46.870 ;
        POLYGON 171.680 47.360 171.680 47.315 171.675 47.315 ;
        RECT 171.680 47.315 175.685 47.365 ;
        POLYGON 171.675 47.315 171.675 46.870 171.630 46.870 ;
        RECT 171.675 46.870 175.685 47.315 ;
        RECT 166.840 46.860 168.840 46.870 ;
        POLYGON 166.825 46.860 166.825 46.725 166.800 46.725 ;
        RECT 166.825 46.725 168.840 46.860 ;
        RECT 163.905 46.575 165.140 46.710 ;
        POLYGON 163.845 46.575 163.845 46.380 163.775 46.380 ;
        RECT 163.845 46.520 165.140 46.575 ;
        POLYGON 165.140 46.710 165.190 46.710 165.140 46.520 ;
        POLYGON 166.800 46.710 166.800 46.695 166.795 46.695 ;
        RECT 166.800 46.695 168.840 46.725 ;
        POLYGON 166.795 46.695 166.795 46.690 166.790 46.690 ;
        RECT 166.795 46.690 168.840 46.695 ;
        POLYGON 166.790 46.690 166.790 46.530 166.755 46.530 ;
        RECT 166.790 46.620 168.840 46.690 ;
        POLYGON 168.840 46.870 168.890 46.870 168.840 46.620 ;
        POLYGON 171.630 46.870 171.630 46.670 171.610 46.670 ;
        RECT 171.630 46.670 175.685 46.870 ;
        POLYGON 171.610 46.670 171.610 46.625 171.605 46.625 ;
        RECT 171.610 46.625 175.685 46.670 ;
        RECT 166.790 46.530 168.795 46.620 ;
        RECT 163.845 46.455 165.125 46.520 ;
        POLYGON 165.125 46.520 165.140 46.520 165.125 46.455 ;
        POLYGON 166.755 46.520 166.755 46.465 166.740 46.465 ;
        RECT 166.755 46.465 168.795 46.530 ;
        RECT 163.845 46.380 165.090 46.455 ;
        POLYGON 163.775 46.380 163.775 46.365 163.770 46.365 ;
        RECT 163.775 46.365 165.090 46.380 ;
        RECT 161.905 46.325 162.790 46.355 ;
        RECT 160.535 46.295 161.040 46.320 ;
        POLYGON 160.490 46.295 160.490 46.280 160.475 46.280 ;
        RECT 160.490 46.280 161.040 46.295 ;
        RECT 159.415 46.250 159.910 46.280 ;
        POLYGON 159.335 46.250 159.335 46.235 159.325 46.235 ;
        RECT 159.335 46.245 159.910 46.250 ;
        POLYGON 159.910 46.280 159.940 46.280 159.910 46.245 ;
        POLYGON 160.475 46.280 160.475 46.245 160.450 46.245 ;
        RECT 160.475 46.245 161.040 46.280 ;
        RECT 159.335 46.235 159.800 46.245 ;
        RECT 151.385 46.225 158.215 46.235 ;
        POLYGON 158.215 46.235 158.230 46.235 158.215 46.225 ;
        POLYGON 159.325 46.235 159.325 46.225 159.315 46.225 ;
        RECT 159.325 46.225 159.800 46.235 ;
        RECT 151.385 46.220 158.190 46.225 ;
        RECT 117.245 46.205 150.340 46.220 ;
        POLYGON 150.340 46.220 150.355 46.205 150.340 46.205 ;
        POLYGON 151.385 46.220 151.400 46.220 151.400 46.205 ;
        RECT 151.400 46.205 158.190 46.220 ;
        RECT 117.245 46.185 150.355 46.205 ;
        POLYGON 150.355 46.205 150.370 46.185 150.355 46.185 ;
        POLYGON 151.400 46.205 151.425 46.205 151.425 46.185 ;
        RECT 151.425 46.200 158.190 46.205 ;
        POLYGON 158.190 46.225 158.215 46.225 158.190 46.200 ;
        POLYGON 159.315 46.225 159.315 46.200 159.290 46.200 ;
        RECT 159.315 46.200 159.800 46.225 ;
        RECT 151.425 46.185 158.050 46.200 ;
        RECT 117.245 46.115 150.370 46.185 ;
        POLYGON 150.370 46.185 150.430 46.115 150.370 46.115 ;
        POLYGON 151.425 46.185 151.465 46.185 151.465 46.150 ;
        RECT 151.465 46.150 158.050 46.185 ;
        POLYGON 151.465 46.150 151.475 46.150 151.475 46.140 ;
        RECT 151.475 46.140 158.050 46.150 ;
        POLYGON 151.475 46.140 151.500 46.140 151.500 46.115 ;
        RECT 151.500 46.115 158.050 46.140 ;
        RECT 117.245 46.095 150.430 46.115 ;
        POLYGON 150.430 46.115 150.450 46.095 150.430 46.095 ;
        POLYGON 151.500 46.115 151.520 46.115 151.520 46.100 ;
        RECT 151.520 46.100 158.050 46.115 ;
        POLYGON 151.520 46.100 151.525 46.100 151.525 46.095 ;
        RECT 151.525 46.095 158.050 46.100 ;
        RECT 117.245 46.085 150.450 46.095 ;
        RECT 117.245 46.075 149.940 46.085 ;
        POLYGON 149.940 46.085 149.945 46.085 149.945 46.080 ;
        RECT 149.945 46.080 150.450 46.085 ;
        POLYGON 149.940 46.080 149.945 46.075 149.940 46.075 ;
        RECT 117.245 46.055 149.945 46.075 ;
        POLYGON 149.945 46.080 149.955 46.080 149.955 46.070 ;
        RECT 149.955 46.070 150.450 46.080 ;
        POLYGON 149.945 46.070 149.955 46.055 149.945 46.055 ;
        RECT 117.245 46.010 149.955 46.055 ;
        POLYGON 149.955 46.070 149.975 46.070 149.975 46.050 ;
        RECT 149.975 46.055 150.450 46.070 ;
        POLYGON 150.450 46.095 150.485 46.055 150.450 46.055 ;
        POLYGON 151.525 46.095 151.570 46.095 151.570 46.055 ;
        RECT 151.570 46.085 158.050 46.095 ;
        POLYGON 158.050 46.200 158.190 46.200 158.050 46.085 ;
        POLYGON 159.290 46.200 159.290 46.180 159.275 46.180 ;
        RECT 159.290 46.180 159.800 46.200 ;
        POLYGON 159.275 46.180 159.275 46.150 159.250 46.150 ;
        RECT 159.275 46.150 159.800 46.180 ;
        POLYGON 159.250 46.150 159.250 46.085 159.190 46.085 ;
        RECT 159.250 46.110 159.800 46.150 ;
        POLYGON 159.800 46.245 159.910 46.245 159.800 46.110 ;
        POLYGON 160.450 46.245 160.450 46.170 160.400 46.170 ;
        RECT 160.450 46.170 161.040 46.245 ;
        POLYGON 160.400 46.170 160.400 46.145 160.385 46.145 ;
        RECT 160.400 46.145 161.040 46.170 ;
        POLYGON 160.385 46.145 160.385 46.110 160.360 46.110 ;
        RECT 160.385 46.110 161.040 46.145 ;
        RECT 159.250 46.085 159.770 46.110 ;
        RECT 151.570 46.055 157.945 46.085 ;
        RECT 149.975 46.050 150.485 46.055 ;
        POLYGON 149.955 46.050 149.975 46.010 149.955 46.010 ;
        POLYGON 149.975 46.050 150.010 46.050 150.010 46.010 ;
        RECT 150.010 46.030 150.485 46.050 ;
        POLYGON 150.485 46.055 150.505 46.030 150.485 46.030 ;
        POLYGON 151.570 46.055 151.600 46.055 151.600 46.030 ;
        RECT 151.600 46.030 157.945 46.055 ;
        RECT 150.010 46.010 150.505 46.030 ;
        RECT 117.245 45.995 149.975 46.010 ;
        POLYGON 149.975 46.010 149.980 45.995 149.975 45.995 ;
        POLYGON 150.010 46.010 150.020 46.010 150.020 45.995 ;
        RECT 150.020 45.995 150.505 46.010 ;
        RECT 117.245 45.975 149.980 45.995 ;
        POLYGON 149.980 45.995 149.990 45.975 149.980 45.975 ;
        RECT 117.245 45.940 149.990 45.975 ;
        POLYGON 150.020 45.995 150.050 45.995 150.050 45.965 ;
        RECT 150.050 45.980 150.505 45.995 ;
        POLYGON 150.505 46.030 150.555 45.980 150.505 45.980 ;
        POLYGON 151.600 46.030 151.635 46.030 151.635 46.000 ;
        RECT 151.635 46.000 157.945 46.030 ;
        POLYGON 157.945 46.085 158.050 46.085 157.945 46.000 ;
        POLYGON 159.190 46.085 159.190 46.020 159.130 46.020 ;
        RECT 159.190 46.075 159.770 46.085 ;
        POLYGON 159.770 46.110 159.800 46.110 159.770 46.075 ;
        POLYGON 160.360 46.110 160.360 46.090 160.345 46.090 ;
        RECT 160.360 46.090 161.040 46.110 ;
        POLYGON 160.345 46.090 160.345 46.075 160.335 46.075 ;
        RECT 160.345 46.075 161.040 46.090 ;
        RECT 159.190 46.020 159.620 46.075 ;
        POLYGON 159.130 46.020 159.130 46.000 159.115 46.000 ;
        RECT 159.130 46.000 159.620 46.020 ;
        POLYGON 151.640 46.000 151.660 46.000 151.660 45.980 ;
        RECT 151.660 45.980 157.885 46.000 ;
        RECT 150.050 45.965 150.555 45.980 ;
        POLYGON 149.990 45.965 150.005 45.940 149.990 45.940 ;
        RECT 117.245 45.915 150.005 45.940 ;
        POLYGON 150.050 45.965 150.075 45.965 150.075 45.935 ;
        RECT 150.075 45.935 150.555 45.965 ;
        POLYGON 150.005 45.935 150.015 45.915 150.005 45.915 ;
        RECT 117.245 45.840 150.015 45.915 ;
        POLYGON 150.075 45.935 150.095 45.935 150.095 45.910 ;
        RECT 150.095 45.925 150.555 45.935 ;
        POLYGON 150.555 45.980 150.605 45.925 150.555 45.925 ;
        POLYGON 151.660 45.980 151.730 45.980 151.730 45.925 ;
        RECT 151.730 45.950 157.885 45.980 ;
        POLYGON 157.885 46.000 157.945 46.000 157.885 45.950 ;
        POLYGON 159.115 46.000 159.115 45.950 159.065 45.950 ;
        RECT 159.115 45.950 159.620 46.000 ;
        RECT 151.730 45.925 157.780 45.950 ;
        RECT 150.095 45.910 150.605 45.925 ;
        RECT 55.200 45.690 112.885 45.840 ;
        POLYGON 112.885 45.840 112.930 45.690 112.885 45.690 ;
        POLYGON 117.245 45.840 117.250 45.840 117.250 45.735 ;
        RECT 117.250 45.835 150.015 45.840 ;
        POLYGON 150.015 45.910 150.050 45.835 150.015 45.835 ;
        POLYGON 150.095 45.910 150.170 45.910 150.170 45.835 ;
        RECT 150.170 45.875 150.605 45.910 ;
        POLYGON 150.605 45.925 150.655 45.875 150.605 45.875 ;
        POLYGON 151.730 45.925 151.795 45.925 151.795 45.875 ;
        RECT 151.795 45.875 157.780 45.925 ;
        POLYGON 157.780 45.950 157.885 45.950 157.780 45.875 ;
        POLYGON 159.065 45.950 159.065 45.875 158.990 45.875 ;
        RECT 159.065 45.910 159.620 45.950 ;
        POLYGON 159.620 46.075 159.770 46.075 159.620 45.910 ;
        POLYGON 160.335 46.075 160.335 46.050 160.315 46.050 ;
        RECT 160.335 46.070 161.040 46.075 ;
        POLYGON 161.040 46.320 161.190 46.320 161.040 46.070 ;
        POLYGON 161.880 46.320 161.880 46.260 161.850 46.260 ;
        RECT 161.880 46.285 162.790 46.325 ;
        POLYGON 162.790 46.355 162.825 46.355 162.790 46.285 ;
        POLYGON 163.770 46.360 163.770 46.285 163.740 46.285 ;
        RECT 163.770 46.325 165.090 46.365 ;
        POLYGON 165.090 46.455 165.125 46.455 165.090 46.325 ;
        POLYGON 166.740 46.455 166.740 46.440 166.735 46.440 ;
        RECT 166.740 46.440 168.795 46.465 ;
        POLYGON 166.735 46.440 166.735 46.380 166.720 46.380 ;
        RECT 166.735 46.380 168.795 46.440 ;
        POLYGON 166.720 46.380 166.720 46.330 166.705 46.330 ;
        RECT 166.720 46.375 168.795 46.380 ;
        POLYGON 168.795 46.620 168.840 46.620 168.795 46.375 ;
        POLYGON 171.605 46.620 171.605 46.580 171.600 46.580 ;
        RECT 171.605 46.580 175.685 46.625 ;
        POLYGON 171.600 46.580 171.600 46.375 171.570 46.375 ;
        RECT 171.600 46.375 175.685 46.580 ;
        RECT 166.720 46.330 168.685 46.375 ;
        RECT 163.770 46.285 165.055 46.325 ;
        RECT 161.880 46.260 162.630 46.285 ;
        POLYGON 161.850 46.260 161.850 46.110 161.770 46.110 ;
        RECT 161.850 46.110 162.630 46.260 ;
        POLYGON 161.770 46.110 161.770 46.095 161.765 46.095 ;
        RECT 161.770 46.095 162.630 46.110 ;
        POLYGON 161.765 46.095 161.765 46.070 161.750 46.070 ;
        RECT 161.765 46.070 162.630 46.095 ;
        RECT 160.335 46.050 160.975 46.070 ;
        POLYGON 160.315 46.050 160.315 46.005 160.280 46.005 ;
        RECT 160.315 46.005 160.975 46.050 ;
        POLYGON 160.280 46.005 160.280 45.910 160.210 45.910 ;
        RECT 160.280 45.965 160.975 46.005 ;
        POLYGON 160.975 46.070 161.040 46.070 160.975 45.965 ;
        POLYGON 161.750 46.070 161.750 45.965 161.685 45.965 ;
        RECT 161.750 45.965 162.630 46.070 ;
        RECT 160.280 45.910 160.905 45.965 ;
        RECT 159.065 45.875 159.580 45.910 ;
        RECT 150.170 45.835 150.655 45.875 ;
        RECT 117.250 45.720 150.050 45.835 ;
        POLYGON 150.050 45.835 150.100 45.720 150.050 45.720 ;
        POLYGON 150.170 45.835 150.280 45.835 150.280 45.720 ;
        RECT 150.280 45.830 150.655 45.835 ;
        POLYGON 150.655 45.875 150.695 45.830 150.655 45.830 ;
        POLYGON 151.795 45.875 151.805 45.875 151.805 45.870 ;
        RECT 151.805 45.870 157.715 45.875 ;
        POLYGON 151.810 45.870 151.860 45.870 151.860 45.830 ;
        RECT 151.860 45.830 157.715 45.870 ;
        RECT 150.280 45.825 150.695 45.830 ;
        POLYGON 150.695 45.830 150.700 45.825 150.695 45.825 ;
        POLYGON 151.860 45.830 151.865 45.830 151.865 45.825 ;
        RECT 151.865 45.825 157.715 45.830 ;
        POLYGON 157.715 45.875 157.780 45.875 157.715 45.825 ;
        POLYGON 158.990 45.875 158.990 45.825 158.940 45.825 ;
        RECT 158.990 45.865 159.580 45.875 ;
        POLYGON 159.580 45.910 159.620 45.910 159.580 45.865 ;
        POLYGON 160.210 45.910 160.210 45.905 160.205 45.905 ;
        RECT 160.210 45.905 160.905 45.910 ;
        POLYGON 160.205 45.905 160.205 45.870 160.175 45.870 ;
        RECT 160.205 45.870 160.905 45.905 ;
        RECT 158.990 45.825 159.495 45.865 ;
        RECT 150.280 45.795 150.700 45.825 ;
        POLYGON 150.700 45.825 150.735 45.795 150.700 45.795 ;
        POLYGON 151.865 45.825 151.875 45.825 151.875 45.820 ;
        RECT 151.875 45.820 157.665 45.825 ;
        POLYGON 151.875 45.820 151.910 45.820 151.910 45.795 ;
        RECT 151.910 45.795 157.665 45.820 ;
        RECT 150.280 45.765 150.735 45.795 ;
        POLYGON 150.735 45.795 150.765 45.765 150.735 45.765 ;
        POLYGON 151.910 45.795 151.955 45.795 151.955 45.765 ;
        RECT 151.955 45.790 157.665 45.795 ;
        POLYGON 157.665 45.825 157.715 45.825 157.665 45.790 ;
        POLYGON 158.940 45.825 158.940 45.790 158.905 45.790 ;
        RECT 158.940 45.790 159.495 45.825 ;
        RECT 151.955 45.765 157.545 45.790 ;
        RECT 150.280 45.720 150.765 45.765 ;
        RECT 55.200 45.200 112.930 45.690 ;
        POLYGON 55.200 45.200 56.700 45.200 56.700 42.005 ;
        RECT 56.700 43.145 112.930 45.200 ;
        POLYGON 112.930 45.690 113.750 43.145 112.930 43.145 ;
        RECT 117.250 45.685 150.100 45.720 ;
        POLYGON 150.100 45.720 150.115 45.685 150.100 45.685 ;
        RECT 117.250 45.660 150.115 45.685 ;
        POLYGON 150.280 45.720 150.325 45.720 150.325 45.675 ;
        RECT 150.325 45.675 150.765 45.720 ;
        POLYGON 150.115 45.675 150.125 45.660 150.115 45.660 ;
        RECT 117.250 45.640 150.125 45.660 ;
        POLYGON 150.325 45.675 150.340 45.675 150.340 45.655 ;
        RECT 150.340 45.665 150.765 45.675 ;
        POLYGON 150.765 45.765 150.870 45.665 150.765 45.665 ;
        POLYGON 151.955 45.765 152.105 45.765 152.105 45.665 ;
        RECT 152.105 45.710 157.545 45.765 ;
        POLYGON 157.545 45.790 157.665 45.790 157.545 45.710 ;
        POLYGON 158.905 45.790 158.905 45.710 158.825 45.710 ;
        RECT 158.905 45.775 159.495 45.790 ;
        POLYGON 159.495 45.865 159.580 45.865 159.495 45.775 ;
        POLYGON 160.175 45.865 160.175 45.855 160.165 45.855 ;
        RECT 160.175 45.855 160.905 45.870 ;
        POLYGON 160.905 45.965 160.975 45.965 160.905 45.855 ;
        POLYGON 161.685 45.960 161.685 45.945 161.675 45.945 ;
        RECT 161.685 45.950 162.630 45.965 ;
        POLYGON 162.630 46.285 162.790 46.285 162.630 45.950 ;
        POLYGON 163.740 46.285 163.740 46.270 163.735 46.270 ;
        RECT 163.740 46.270 165.055 46.285 ;
        POLYGON 163.735 46.270 163.735 46.155 163.690 46.155 ;
        RECT 163.735 46.210 165.055 46.270 ;
        POLYGON 165.055 46.325 165.090 46.325 165.055 46.210 ;
        POLYGON 166.705 46.325 166.705 46.210 166.670 46.210 ;
        RECT 166.705 46.210 168.685 46.330 ;
        RECT 163.735 46.155 164.980 46.210 ;
        POLYGON 163.690 46.155 163.690 46.090 163.665 46.090 ;
        RECT 163.690 46.090 164.980 46.155 ;
        POLYGON 163.665 46.090 163.665 45.965 163.610 45.965 ;
        RECT 163.665 45.970 164.980 46.090 ;
        POLYGON 164.980 46.210 165.055 46.210 164.980 45.970 ;
        POLYGON 166.670 46.210 166.670 46.195 166.665 46.195 ;
        RECT 166.670 46.195 168.685 46.210 ;
        POLYGON 166.665 46.185 166.665 46.090 166.635 46.090 ;
        RECT 166.665 46.090 168.685 46.195 ;
        POLYGON 166.635 46.090 166.635 45.975 166.595 45.975 ;
        RECT 166.635 45.975 168.685 46.090 ;
        RECT 163.665 45.965 164.895 45.970 ;
        POLYGON 163.610 45.965 163.610 45.955 163.605 45.955 ;
        RECT 163.610 45.955 164.895 45.965 ;
        RECT 161.685 45.945 162.525 45.950 ;
        POLYGON 161.675 45.945 161.675 45.855 161.625 45.855 ;
        RECT 161.675 45.855 162.525 45.945 ;
        POLYGON 160.165 45.855 160.165 45.825 160.145 45.825 ;
        RECT 160.165 45.825 160.880 45.855 ;
        POLYGON 160.145 45.825 160.145 45.805 160.130 45.805 ;
        RECT 160.145 45.820 160.880 45.825 ;
        POLYGON 160.880 45.855 160.905 45.855 160.880 45.820 ;
        POLYGON 161.625 45.855 161.625 45.845 161.620 45.845 ;
        RECT 161.625 45.845 162.525 45.855 ;
        POLYGON 161.620 45.845 161.620 45.820 161.605 45.820 ;
        RECT 161.620 45.820 162.525 45.845 ;
        RECT 160.145 45.805 160.710 45.820 ;
        POLYGON 160.130 45.805 160.130 45.775 160.105 45.775 ;
        RECT 160.130 45.775 160.710 45.805 ;
        RECT 158.905 45.740 159.465 45.775 ;
        POLYGON 159.465 45.775 159.495 45.775 159.465 45.740 ;
        POLYGON 160.105 45.775 160.105 45.740 160.075 45.740 ;
        RECT 160.105 45.740 160.710 45.775 ;
        RECT 158.905 45.710 159.355 45.740 ;
        RECT 152.105 45.665 157.385 45.710 ;
        RECT 150.340 45.655 150.870 45.665 ;
        POLYGON 150.870 45.665 150.880 45.655 150.870 45.655 ;
        POLYGON 152.105 45.665 152.120 45.665 152.120 45.655 ;
        RECT 152.120 45.655 157.385 45.665 ;
        POLYGON 117.250 45.640 117.265 45.640 117.265 44.935 ;
        RECT 117.265 45.625 150.125 45.640 ;
        POLYGON 150.125 45.655 150.140 45.625 150.125 45.625 ;
        RECT 117.265 45.545 150.140 45.625 ;
        POLYGON 150.340 45.655 150.375 45.655 150.375 45.620 ;
        RECT 150.375 45.635 150.880 45.655 ;
        POLYGON 150.880 45.655 150.905 45.635 150.880 45.635 ;
        POLYGON 152.120 45.655 152.150 45.655 152.150 45.635 ;
        RECT 152.150 45.635 157.385 45.655 ;
        RECT 150.375 45.620 150.905 45.635 ;
        POLYGON 150.140 45.620 150.175 45.545 150.140 45.545 ;
        RECT 117.265 45.520 150.175 45.545 ;
        POLYGON 150.375 45.620 150.460 45.620 150.460 45.540 ;
        RECT 150.460 45.555 150.905 45.620 ;
        POLYGON 150.905 45.635 151.000 45.555 150.905 45.555 ;
        POLYGON 152.150 45.635 152.160 45.635 152.160 45.630 ;
        RECT 152.160 45.630 157.385 45.635 ;
        POLYGON 152.165 45.630 152.260 45.630 152.260 45.570 ;
        RECT 152.260 45.610 157.385 45.630 ;
        POLYGON 157.385 45.710 157.545 45.710 157.385 45.610 ;
        POLYGON 158.825 45.710 158.825 45.675 158.790 45.675 ;
        RECT 158.825 45.675 159.355 45.710 ;
        POLYGON 158.790 45.675 158.790 45.610 158.720 45.610 ;
        RECT 158.790 45.635 159.355 45.675 ;
        POLYGON 159.355 45.740 159.465 45.740 159.355 45.635 ;
        POLYGON 160.075 45.740 160.075 45.705 160.045 45.705 ;
        RECT 160.075 45.705 160.710 45.740 ;
        POLYGON 160.045 45.705 160.045 45.660 160.005 45.660 ;
        RECT 160.045 45.660 160.710 45.705 ;
        POLYGON 160.005 45.660 160.005 45.635 159.985 45.635 ;
        RECT 160.005 45.635 160.710 45.660 ;
        RECT 158.790 45.610 159.300 45.635 ;
        RECT 152.260 45.600 157.370 45.610 ;
        POLYGON 157.370 45.610 157.385 45.610 157.370 45.600 ;
        POLYGON 158.720 45.610 158.720 45.600 158.710 45.600 ;
        RECT 158.720 45.600 159.300 45.610 ;
        RECT 152.260 45.595 157.365 45.600 ;
        POLYGON 157.365 45.600 157.370 45.600 157.365 45.595 ;
        POLYGON 158.710 45.600 158.710 45.595 158.705 45.595 ;
        RECT 158.710 45.595 159.300 45.600 ;
        RECT 152.260 45.570 157.195 45.595 ;
        POLYGON 152.260 45.570 152.280 45.570 152.280 45.555 ;
        RECT 152.280 45.555 157.195 45.570 ;
        RECT 150.460 45.545 151.000 45.555 ;
        POLYGON 151.000 45.555 151.010 45.545 151.000 45.545 ;
        POLYGON 152.280 45.555 152.300 45.555 152.300 45.545 ;
        RECT 152.300 45.545 157.195 45.555 ;
        RECT 150.460 45.540 151.010 45.545 ;
        POLYGON 150.175 45.540 150.185 45.520 150.175 45.520 ;
        RECT 117.265 45.475 150.185 45.520 ;
        POLYGON 150.460 45.540 150.490 45.540 150.490 45.515 ;
        RECT 150.490 45.515 151.010 45.540 ;
        POLYGON 150.185 45.515 150.205 45.475 150.185 45.475 ;
        RECT 117.265 45.465 150.205 45.475 ;
        POLYGON 150.490 45.515 150.540 45.515 150.540 45.470 ;
        RECT 150.540 45.490 151.010 45.515 ;
        POLYGON 151.010 45.545 151.075 45.490 151.010 45.490 ;
        POLYGON 152.300 45.545 152.350 45.545 152.350 45.520 ;
        RECT 152.350 45.520 157.195 45.545 ;
        POLYGON 152.350 45.520 152.395 45.520 152.395 45.490 ;
        RECT 152.395 45.500 157.195 45.520 ;
        POLYGON 157.195 45.595 157.365 45.595 157.195 45.500 ;
        POLYGON 158.705 45.595 158.705 45.545 158.650 45.545 ;
        RECT 158.705 45.580 159.300 45.595 ;
        POLYGON 159.300 45.635 159.355 45.635 159.300 45.580 ;
        POLYGON 159.985 45.635 159.985 45.580 159.940 45.580 ;
        RECT 159.985 45.580 160.710 45.635 ;
        POLYGON 160.710 45.820 160.880 45.820 160.710 45.580 ;
        POLYGON 161.605 45.820 161.605 45.760 161.570 45.760 ;
        RECT 161.605 45.760 162.525 45.820 ;
        POLYGON 162.525 45.950 162.630 45.950 162.525 45.760 ;
        POLYGON 163.605 45.950 163.605 45.820 163.545 45.820 ;
        RECT 163.605 45.820 164.895 45.955 ;
        POLYGON 163.545 45.820 163.545 45.800 163.540 45.800 ;
        RECT 163.545 45.800 164.895 45.820 ;
        POLYGON 163.540 45.800 163.540 45.760 163.520 45.760 ;
        RECT 163.540 45.760 164.895 45.800 ;
        POLYGON 161.570 45.760 161.570 45.735 161.555 45.735 ;
        RECT 161.570 45.735 162.440 45.760 ;
        POLYGON 161.555 45.735 161.555 45.705 161.540 45.705 ;
        RECT 161.555 45.705 162.440 45.735 ;
        POLYGON 161.540 45.705 161.540 45.585 161.460 45.585 ;
        RECT 161.540 45.605 162.440 45.705 ;
        POLYGON 162.440 45.760 162.525 45.760 162.440 45.605 ;
        POLYGON 163.520 45.760 163.520 45.730 163.505 45.730 ;
        RECT 163.520 45.740 164.895 45.760 ;
        POLYGON 164.895 45.970 164.980 45.970 164.895 45.740 ;
        POLYGON 166.595 45.970 166.595 45.930 166.580 45.930 ;
        RECT 166.595 45.930 168.685 45.975 ;
        POLYGON 166.580 45.930 166.580 45.800 166.535 45.800 ;
        RECT 166.580 45.885 168.685 45.930 ;
        POLYGON 168.685 46.375 168.795 46.375 168.685 45.885 ;
        POLYGON 171.570 46.375 171.570 45.935 171.505 45.935 ;
        RECT 171.570 45.935 175.685 46.375 ;
        POLYGON 171.505 45.935 171.505 45.885 171.495 45.885 ;
        RECT 171.505 45.885 175.685 45.935 ;
        RECT 166.580 45.800 168.555 45.885 ;
        POLYGON 166.535 45.800 166.535 45.750 166.515 45.750 ;
        RECT 166.535 45.750 168.555 45.800 ;
        POLYGON 166.515 45.750 166.515 45.740 166.510 45.740 ;
        RECT 166.515 45.740 168.555 45.750 ;
        RECT 163.520 45.730 164.795 45.740 ;
        POLYGON 163.505 45.730 163.505 45.610 163.450 45.610 ;
        RECT 163.505 45.610 164.795 45.730 ;
        RECT 161.540 45.585 162.410 45.605 ;
        RECT 158.705 45.545 159.260 45.580 ;
        POLYGON 159.260 45.580 159.300 45.580 159.260 45.545 ;
        POLYGON 159.940 45.580 159.940 45.565 159.930 45.565 ;
        RECT 159.940 45.565 160.615 45.580 ;
        POLYGON 159.930 45.565 159.930 45.550 159.910 45.550 ;
        RECT 159.930 45.550 160.615 45.565 ;
        POLYGON 159.910 45.550 159.910 45.545 159.905 45.545 ;
        RECT 159.910 45.545 160.615 45.550 ;
        POLYGON 158.650 45.545 158.650 45.525 158.630 45.525 ;
        RECT 158.650 45.525 159.130 45.545 ;
        POLYGON 158.630 45.525 158.630 45.500 158.600 45.500 ;
        RECT 158.630 45.500 159.130 45.525 ;
        RECT 152.395 45.490 157.150 45.500 ;
        RECT 150.540 45.470 151.075 45.490 ;
        POLYGON 150.205 45.470 150.210 45.465 150.205 45.465 ;
        RECT 117.265 45.430 150.210 45.465 ;
        POLYGON 150.540 45.470 150.555 45.470 150.555 45.455 ;
        RECT 150.555 45.455 151.075 45.470 ;
        POLYGON 151.075 45.490 151.120 45.455 151.075 45.455 ;
        POLYGON 152.395 45.490 152.415 45.490 152.415 45.480 ;
        RECT 152.415 45.480 157.150 45.490 ;
        POLYGON 152.415 45.480 152.460 45.480 152.460 45.455 ;
        RECT 152.460 45.475 157.150 45.480 ;
        POLYGON 157.150 45.500 157.195 45.500 157.150 45.475 ;
        POLYGON 158.600 45.500 158.600 45.485 158.580 45.485 ;
        RECT 158.600 45.485 159.130 45.500 ;
        POLYGON 158.580 45.485 158.580 45.475 158.570 45.475 ;
        RECT 158.580 45.475 159.130 45.485 ;
        RECT 152.460 45.455 157.110 45.475 ;
        POLYGON 157.110 45.475 157.150 45.475 157.110 45.455 ;
        POLYGON 158.570 45.475 158.570 45.455 158.545 45.455 ;
        RECT 158.570 45.455 159.130 45.475 ;
        POLYGON 150.210 45.455 150.225 45.430 150.210 45.430 ;
        RECT 117.265 45.405 150.225 45.430 ;
        POLYGON 150.555 45.455 150.590 45.455 150.590 45.420 ;
        RECT 150.590 45.450 151.120 45.455 ;
        POLYGON 151.120 45.455 151.125 45.450 151.120 45.450 ;
        POLYGON 152.460 45.455 152.470 45.455 152.470 45.450 ;
        RECT 152.470 45.450 157.020 45.455 ;
        RECT 150.590 45.425 151.125 45.450 ;
        POLYGON 151.125 45.450 151.160 45.425 151.125 45.425 ;
        POLYGON 152.470 45.450 152.500 45.450 152.500 45.435 ;
        RECT 152.500 45.435 157.020 45.450 ;
        POLYGON 152.505 45.435 152.520 45.435 152.520 45.425 ;
        RECT 152.520 45.425 157.020 45.435 ;
        RECT 150.590 45.420 151.160 45.425 ;
        POLYGON 150.225 45.420 150.235 45.405 150.225 45.405 ;
        RECT 117.265 45.360 150.235 45.405 ;
        POLYGON 150.590 45.420 150.615 45.420 150.615 45.400 ;
        RECT 150.615 45.400 151.160 45.420 ;
        POLYGON 150.235 45.400 150.255 45.360 150.235 45.360 ;
        POLYGON 150.615 45.400 150.655 45.400 150.655 45.360 ;
        RECT 150.655 45.360 151.160 45.400 ;
        RECT 117.265 45.290 150.255 45.360 ;
        POLYGON 150.255 45.360 150.285 45.290 150.255 45.290 ;
        POLYGON 150.655 45.360 150.695 45.360 150.695 45.325 ;
        RECT 150.695 45.355 151.160 45.360 ;
        POLYGON 151.160 45.425 151.250 45.355 151.160 45.355 ;
        POLYGON 152.520 45.425 152.535 45.425 152.535 45.415 ;
        RECT 152.535 45.415 157.020 45.425 ;
        POLYGON 152.535 45.415 152.575 45.415 152.575 45.395 ;
        RECT 152.575 45.405 157.020 45.415 ;
        POLYGON 157.020 45.455 157.110 45.455 157.020 45.405 ;
        POLYGON 158.545 45.455 158.545 45.425 158.510 45.425 ;
        RECT 158.545 45.425 159.130 45.455 ;
        POLYGON 158.510 45.425 158.510 45.405 158.490 45.405 ;
        RECT 158.510 45.420 159.130 45.425 ;
        POLYGON 159.130 45.545 159.260 45.545 159.130 45.420 ;
        POLYGON 159.905 45.545 159.905 45.425 159.800 45.425 ;
        RECT 159.905 45.455 160.615 45.545 ;
        POLYGON 160.615 45.580 160.710 45.580 160.615 45.455 ;
        POLYGON 161.460 45.580 161.460 45.575 161.455 45.575 ;
        RECT 161.460 45.575 162.410 45.585 ;
        POLYGON 161.455 45.575 161.455 45.455 161.375 45.455 ;
        RECT 161.455 45.555 162.410 45.575 ;
        POLYGON 162.410 45.605 162.440 45.605 162.410 45.555 ;
        POLYGON 163.450 45.605 163.450 45.590 163.440 45.590 ;
        RECT 163.450 45.590 164.795 45.610 ;
        POLYGON 163.440 45.590 163.440 45.560 163.425 45.560 ;
        RECT 163.440 45.560 164.795 45.590 ;
        RECT 161.455 45.455 162.210 45.555 ;
        RECT 159.905 45.425 160.540 45.455 ;
        POLYGON 159.800 45.425 159.800 45.420 159.795 45.420 ;
        RECT 159.800 45.420 160.540 45.425 ;
        RECT 158.510 45.405 159.015 45.420 ;
        RECT 152.575 45.395 156.975 45.405 ;
        POLYGON 152.575 45.395 152.660 45.395 152.660 45.355 ;
        RECT 152.660 45.385 156.975 45.395 ;
        POLYGON 156.975 45.405 157.020 45.405 156.975 45.385 ;
        POLYGON 158.490 45.405 158.490 45.385 158.465 45.385 ;
        RECT 158.490 45.385 159.015 45.405 ;
        RECT 152.660 45.370 156.940 45.385 ;
        POLYGON 156.940 45.385 156.975 45.385 156.940 45.370 ;
        POLYGON 158.465 45.385 158.465 45.370 158.450 45.370 ;
        RECT 158.465 45.370 159.015 45.385 ;
        RECT 152.660 45.355 156.845 45.370 ;
        RECT 150.695 45.325 151.250 45.355 ;
        RECT 117.265 45.265 150.285 45.290 ;
        POLYGON 150.695 45.325 150.740 45.325 150.740 45.285 ;
        RECT 150.740 45.305 151.250 45.325 ;
        POLYGON 151.250 45.355 151.310 45.305 151.250 45.305 ;
        POLYGON 152.660 45.355 152.715 45.355 152.715 45.330 ;
        RECT 152.715 45.330 156.845 45.355 ;
        POLYGON 152.715 45.330 152.730 45.330 152.730 45.325 ;
        RECT 152.730 45.325 156.845 45.330 ;
        POLYGON 152.730 45.325 152.770 45.325 152.770 45.305 ;
        RECT 152.770 45.320 156.845 45.325 ;
        POLYGON 156.845 45.370 156.940 45.370 156.845 45.320 ;
        POLYGON 158.450 45.370 158.450 45.345 158.420 45.345 ;
        RECT 158.450 45.345 159.015 45.370 ;
        POLYGON 158.420 45.345 158.420 45.320 158.385 45.320 ;
        RECT 158.420 45.325 159.015 45.345 ;
        POLYGON 159.015 45.420 159.125 45.420 159.015 45.325 ;
        POLYGON 159.795 45.420 159.795 45.395 159.770 45.395 ;
        RECT 159.795 45.395 160.540 45.420 ;
        POLYGON 159.770 45.395 159.770 45.345 159.725 45.345 ;
        RECT 159.770 45.360 160.540 45.395 ;
        POLYGON 160.540 45.455 160.615 45.455 160.540 45.360 ;
        POLYGON 161.375 45.450 161.375 45.360 161.315 45.360 ;
        RECT 161.375 45.360 162.210 45.455 ;
        RECT 159.770 45.350 160.535 45.360 ;
        POLYGON 160.535 45.360 160.540 45.360 160.535 45.350 ;
        POLYGON 161.315 45.360 161.315 45.350 161.310 45.350 ;
        RECT 161.315 45.350 162.210 45.360 ;
        RECT 159.770 45.345 160.345 45.350 ;
        POLYGON 159.725 45.345 159.725 45.325 159.705 45.325 ;
        RECT 159.725 45.325 160.345 45.345 ;
        RECT 158.420 45.320 158.950 45.325 ;
        RECT 152.770 45.305 156.725 45.320 ;
        RECT 150.740 45.285 151.315 45.305 ;
        POLYGON 151.315 45.305 151.340 45.285 151.315 45.285 ;
        POLYGON 152.770 45.305 152.815 45.305 152.815 45.285 ;
        RECT 152.815 45.285 156.725 45.305 ;
        POLYGON 150.285 45.285 150.295 45.265 150.285 45.265 ;
        RECT 117.265 45.175 150.295 45.265 ;
        POLYGON 150.740 45.285 150.770 45.285 150.770 45.260 ;
        RECT 150.770 45.260 151.340 45.285 ;
        POLYGON 150.295 45.260 150.335 45.175 150.295 45.175 ;
        RECT 117.265 45.150 150.335 45.175 ;
        POLYGON 150.770 45.260 150.880 45.260 150.880 45.165 ;
        RECT 150.880 45.255 151.340 45.260 ;
        POLYGON 151.340 45.285 151.385 45.255 151.340 45.255 ;
        POLYGON 152.815 45.285 152.880 45.285 152.880 45.255 ;
        RECT 152.880 45.270 156.725 45.285 ;
        POLYGON 156.725 45.320 156.840 45.320 156.725 45.270 ;
        POLYGON 158.385 45.320 158.385 45.315 158.380 45.315 ;
        RECT 158.385 45.315 158.950 45.320 ;
        POLYGON 158.380 45.315 158.380 45.270 158.325 45.270 ;
        RECT 158.380 45.270 158.950 45.315 ;
        RECT 152.880 45.265 156.715 45.270 ;
        POLYGON 156.715 45.270 156.725 45.270 156.715 45.265 ;
        POLYGON 158.325 45.270 158.325 45.265 158.320 45.265 ;
        RECT 158.325 45.265 158.950 45.270 ;
        POLYGON 158.950 45.325 159.015 45.325 158.950 45.265 ;
        POLYGON 159.705 45.325 159.705 45.265 159.645 45.265 ;
        RECT 159.705 45.265 160.345 45.325 ;
        RECT 152.880 45.255 156.590 45.265 ;
        RECT 150.880 45.200 151.385 45.255 ;
        POLYGON 151.385 45.255 151.465 45.200 151.385 45.200 ;
        POLYGON 152.880 45.255 152.905 45.255 152.905 45.245 ;
        RECT 152.905 45.245 156.590 45.255 ;
        POLYGON 152.905 45.245 152.925 45.245 152.925 45.240 ;
        RECT 152.925 45.240 156.590 45.245 ;
        POLYGON 152.925 45.240 152.930 45.240 152.930 45.235 ;
        RECT 152.930 45.235 156.590 45.240 ;
        POLYGON 152.930 45.235 153.015 45.235 153.015 45.200 ;
        RECT 153.015 45.215 156.590 45.235 ;
        POLYGON 156.590 45.265 156.715 45.265 156.590 45.215 ;
        POLYGON 158.320 45.265 158.320 45.215 158.255 45.215 ;
        RECT 158.320 45.215 158.885 45.265 ;
        POLYGON 158.885 45.265 158.950 45.265 158.885 45.215 ;
        POLYGON 159.645 45.265 159.645 45.215 159.595 45.215 ;
        RECT 159.645 45.215 160.345 45.265 ;
        RECT 153.015 45.200 156.510 45.215 ;
        RECT 150.880 45.195 151.465 45.200 ;
        POLYGON 151.465 45.200 151.470 45.195 151.465 45.195 ;
        POLYGON 153.015 45.200 153.030 45.200 153.030 45.195 ;
        RECT 153.030 45.195 156.510 45.200 ;
        RECT 150.880 45.165 151.475 45.195 ;
        POLYGON 150.335 45.165 150.345 45.150 150.335 45.150 ;
        RECT 117.265 45.140 150.345 45.150 ;
        POLYGON 150.880 45.165 150.905 45.165 150.905 45.145 ;
        RECT 150.905 45.160 151.475 45.165 ;
        POLYGON 151.475 45.195 151.520 45.160 151.475 45.160 ;
        POLYGON 153.030 45.195 153.070 45.195 153.070 45.180 ;
        RECT 153.070 45.185 156.510 45.195 ;
        POLYGON 156.510 45.215 156.590 45.215 156.510 45.185 ;
        POLYGON 158.255 45.215 158.255 45.195 158.230 45.195 ;
        RECT 158.255 45.195 158.765 45.215 ;
        POLYGON 158.230 45.195 158.230 45.185 158.215 45.185 ;
        RECT 158.230 45.185 158.765 45.195 ;
        RECT 153.070 45.180 156.480 45.185 ;
        POLYGON 153.070 45.180 153.120 45.180 153.120 45.165 ;
        RECT 153.120 45.175 156.480 45.180 ;
        POLYGON 156.480 45.185 156.510 45.185 156.480 45.175 ;
        POLYGON 158.215 45.185 158.215 45.175 158.205 45.175 ;
        RECT 158.215 45.175 158.765 45.185 ;
        RECT 153.120 45.165 156.440 45.175 ;
        POLYGON 153.125 45.165 153.135 45.165 153.135 45.160 ;
        RECT 153.135 45.160 156.440 45.165 ;
        POLYGON 156.440 45.175 156.480 45.175 156.440 45.160 ;
        POLYGON 158.205 45.175 158.205 45.165 158.190 45.165 ;
        RECT 158.205 45.165 158.765 45.175 ;
        RECT 150.905 45.145 151.520 45.160 ;
        POLYGON 150.345 45.145 150.350 45.140 150.345 45.140 ;
        RECT 117.265 45.070 150.350 45.140 ;
        POLYGON 150.905 45.145 150.920 45.145 150.920 45.135 ;
        RECT 150.920 45.135 151.520 45.145 ;
        POLYGON 150.350 45.135 150.380 45.070 150.350 45.070 ;
        RECT 117.265 45.020 150.380 45.070 ;
        POLYGON 150.920 45.135 151.010 45.135 151.010 45.065 ;
        RECT 151.010 45.125 151.520 45.135 ;
        POLYGON 151.520 45.160 151.575 45.125 151.520 45.125 ;
        POLYGON 153.135 45.160 153.145 45.160 153.145 45.155 ;
        RECT 153.145 45.155 156.300 45.160 ;
        POLYGON 153.145 45.155 153.225 45.155 153.225 45.125 ;
        RECT 153.225 45.125 156.300 45.155 ;
        RECT 151.010 45.085 151.575 45.125 ;
        POLYGON 151.575 45.125 151.635 45.085 151.575 45.085 ;
        POLYGON 153.225 45.125 153.240 45.125 153.240 45.120 ;
        RECT 153.240 45.120 156.300 45.125 ;
        POLYGON 153.240 45.120 153.325 45.120 153.325 45.095 ;
        RECT 153.325 45.110 156.300 45.120 ;
        POLYGON 156.300 45.160 156.440 45.160 156.300 45.110 ;
        POLYGON 158.190 45.160 158.190 45.110 158.115 45.110 ;
        RECT 158.190 45.120 158.765 45.165 ;
        POLYGON 158.765 45.215 158.885 45.215 158.765 45.120 ;
        POLYGON 159.595 45.215 159.595 45.200 159.580 45.200 ;
        RECT 159.595 45.200 160.345 45.215 ;
        POLYGON 159.580 45.200 159.580 45.135 159.520 45.135 ;
        RECT 159.580 45.135 160.345 45.200 ;
        POLYGON 159.520 45.135 159.520 45.120 159.505 45.120 ;
        RECT 159.520 45.120 160.345 45.135 ;
        POLYGON 160.345 45.350 160.535 45.350 160.345 45.120 ;
        POLYGON 161.310 45.350 161.310 45.340 161.305 45.340 ;
        RECT 161.310 45.340 162.210 45.350 ;
        POLYGON 161.305 45.335 161.305 45.250 161.240 45.250 ;
        RECT 161.305 45.250 162.210 45.340 ;
        POLYGON 161.240 45.250 161.240 45.175 161.190 45.175 ;
        RECT 161.240 45.235 162.210 45.250 ;
        POLYGON 162.210 45.555 162.410 45.555 162.210 45.235 ;
        POLYGON 163.425 45.555 163.425 45.500 163.395 45.500 ;
        RECT 163.425 45.500 164.795 45.560 ;
        POLYGON 163.395 45.500 163.395 45.450 163.370 45.450 ;
        RECT 163.395 45.490 164.795 45.500 ;
        POLYGON 164.795 45.740 164.895 45.740 164.795 45.490 ;
        POLYGON 166.510 45.735 166.510 45.660 166.485 45.660 ;
        RECT 166.510 45.660 168.555 45.740 ;
        POLYGON 166.485 45.660 166.485 45.515 166.425 45.515 ;
        RECT 166.485 45.515 168.555 45.660 ;
        POLYGON 166.425 45.515 166.425 45.490 166.415 45.490 ;
        RECT 166.425 45.490 168.555 45.515 ;
        RECT 163.395 45.450 164.705 45.490 ;
        POLYGON 163.370 45.450 163.370 45.335 163.315 45.335 ;
        RECT 163.370 45.335 164.705 45.450 ;
        POLYGON 163.315 45.335 163.315 45.250 163.270 45.250 ;
        RECT 163.315 45.270 164.705 45.335 ;
        POLYGON 164.705 45.490 164.795 45.490 164.705 45.270 ;
        POLYGON 166.415 45.490 166.415 45.430 166.390 45.430 ;
        RECT 166.415 45.430 168.555 45.490 ;
        POLYGON 166.390 45.430 166.390 45.275 166.325 45.275 ;
        RECT 166.390 45.395 168.555 45.430 ;
        POLYGON 168.555 45.885 168.685 45.885 168.555 45.395 ;
        POLYGON 171.495 45.880 171.495 45.850 171.490 45.850 ;
        RECT 171.495 45.850 175.685 45.885 ;
        POLYGON 171.490 45.850 171.490 45.580 171.435 45.580 ;
        RECT 171.490 45.765 175.685 45.850 ;
        POLYGON 175.685 48.380 175.700 48.380 175.685 45.765 ;
        POLYGON 182.900 48.705 182.935 48.705 182.935 47.185 ;
        POLYGON 182.935 47.185 182.935 45.765 182.900 45.765 ;
        RECT 182.935 46.970 197.600 48.705 ;
        POLYGON 197.600 48.720 197.810 46.970 197.600 46.970 ;
        POLYGON 207.210 48.720 207.230 48.720 207.230 48.615 ;
        RECT 207.230 48.655 222.255 48.720 ;
        POLYGON 222.255 50.495 222.360 48.655 222.255 48.655 ;
        POLYGON 229.225 50.495 229.250 50.495 229.250 49.985 ;
        RECT 229.250 50.270 233.200 50.495 ;
        POLYGON 233.200 51.175 233.220 50.270 233.200 50.270 ;
        POLYGON 235.985 51.390 235.985 50.605 235.975 50.605 ;
        RECT 235.985 51.370 237.985 51.390 ;
        POLYGON 237.985 51.765 238.020 51.765 237.985 51.370 ;
        POLYGON 239.650 51.765 239.650 51.380 239.620 51.380 ;
        RECT 239.650 51.575 240.700 51.765 ;
        POLYGON 240.700 51.865 240.735 51.865 240.700 51.575 ;
        POLYGON 241.700 51.865 241.700 51.710 241.670 51.710 ;
        RECT 241.700 51.855 242.525 51.870 ;
        POLYGON 242.525 51.970 242.550 51.970 242.525 51.855 ;
        POLYGON 243.190 51.980 243.190 51.910 243.170 51.910 ;
        RECT 243.190 51.955 243.675 51.990 ;
        POLYGON 243.675 52.150 243.735 52.150 243.675 51.960 ;
        POLYGON 244.330 52.150 244.330 52.125 244.320 52.125 ;
        RECT 244.330 52.125 245.090 52.150 ;
        POLYGON 244.320 52.125 244.320 52.040 244.295 52.040 ;
        RECT 244.320 52.090 245.090 52.125 ;
        POLYGON 245.090 52.150 245.115 52.150 245.090 52.090 ;
        POLYGON 254.505 52.150 254.525 52.150 254.525 52.120 ;
        RECT 254.525 52.120 255.175 52.150 ;
        POLYGON 254.525 52.120 254.540 52.120 254.540 52.090 ;
        RECT 254.540 52.110 255.175 52.120 ;
        POLYGON 255.175 52.190 255.210 52.110 255.175 52.110 ;
        POLYGON 255.680 52.190 255.705 52.190 255.705 52.120 ;
        RECT 255.705 52.110 256.080 52.190 ;
        RECT 254.540 52.090 255.210 52.110 ;
        RECT 244.320 52.040 245.045 52.090 ;
        POLYGON 244.295 52.040 244.295 51.965 244.275 51.965 ;
        RECT 244.295 51.985 245.045 52.040 ;
        POLYGON 245.045 52.090 245.090 52.090 245.045 51.985 ;
        POLYGON 254.540 52.090 254.570 52.090 254.570 52.035 ;
        RECT 254.570 52.060 255.210 52.090 ;
        POLYGON 255.210 52.110 255.235 52.060 255.210 52.060 ;
        POLYGON 255.705 52.110 255.725 52.110 255.725 52.060 ;
        RECT 255.725 52.085 256.080 52.110 ;
        POLYGON 256.080 52.310 256.175 52.085 256.080 52.085 ;
        POLYGON 256.665 52.310 256.710 52.310 256.710 52.180 ;
        RECT 256.710 52.235 257.235 52.310 ;
        POLYGON 257.235 52.435 257.305 52.235 257.235 52.235 ;
        POLYGON 258.050 52.435 258.085 52.435 258.085 52.350 ;
        RECT 258.085 52.350 258.940 52.435 ;
        POLYGON 258.940 52.590 259.020 52.350 258.940 52.350 ;
        POLYGON 260.150 52.590 260.210 52.590 260.210 52.350 ;
        RECT 260.210 52.420 261.590 52.590 ;
        POLYGON 261.590 52.590 261.635 52.420 261.590 52.420 ;
        POLYGON 263.650 52.590 263.665 52.590 263.665 52.535 ;
        RECT 263.665 52.535 266.340 52.590 ;
        POLYGON 263.665 52.535 263.690 52.535 263.690 52.420 ;
        RECT 263.690 52.495 266.340 52.535 ;
        POLYGON 266.340 52.590 266.365 52.495 266.340 52.495 ;
        POLYGON 270.555 52.590 270.560 52.590 270.560 52.520 ;
        RECT 270.560 52.495 277.425 52.590 ;
        RECT 263.690 52.430 266.365 52.495 ;
        POLYGON 266.365 52.495 266.380 52.430 266.365 52.430 ;
        POLYGON 270.560 52.495 270.565 52.495 270.565 52.450 ;
        RECT 270.565 52.455 277.425 52.495 ;
        POLYGON 277.425 52.590 277.455 52.455 277.425 52.455 ;
        RECT 270.565 52.430 277.455 52.455 ;
        RECT 263.690 52.420 266.380 52.430 ;
        RECT 260.210 52.350 261.635 52.420 ;
        POLYGON 258.085 52.350 258.120 52.350 258.120 52.240 ;
        RECT 258.120 52.315 259.020 52.350 ;
        POLYGON 259.020 52.350 259.030 52.315 259.020 52.315 ;
        POLYGON 260.210 52.350 260.215 52.350 260.215 52.330 ;
        RECT 260.215 52.315 261.635 52.350 ;
        RECT 258.120 52.235 259.030 52.315 ;
        RECT 256.710 52.180 257.305 52.235 ;
        POLYGON 256.710 52.180 256.715 52.180 256.715 52.160 ;
        RECT 256.715 52.160 257.305 52.180 ;
        POLYGON 256.715 52.160 256.735 52.160 256.735 52.105 ;
        RECT 256.735 52.150 257.305 52.160 ;
        POLYGON 257.305 52.235 257.330 52.150 257.305 52.150 ;
        POLYGON 258.120 52.235 258.140 52.235 258.140 52.180 ;
        RECT 258.140 52.180 259.030 52.235 ;
        POLYGON 258.140 52.180 258.145 52.180 258.145 52.160 ;
        RECT 258.145 52.150 259.030 52.180 ;
        RECT 256.735 52.105 257.330 52.150 ;
        POLYGON 256.735 52.105 256.740 52.105 256.740 52.085 ;
        RECT 256.740 52.085 257.330 52.105 ;
        RECT 255.725 52.060 256.175 52.085 ;
        RECT 254.570 52.035 255.235 52.060 ;
        POLYGON 254.570 52.035 254.590 52.035 254.590 51.990 ;
        RECT 254.590 52.010 255.235 52.035 ;
        POLYGON 255.235 52.060 255.255 52.010 255.235 52.010 ;
        POLYGON 255.725 52.060 255.735 52.060 255.735 52.020 ;
        RECT 255.735 52.045 256.175 52.060 ;
        POLYGON 256.175 52.085 256.190 52.045 256.175 52.045 ;
        POLYGON 256.740 52.085 256.750 52.085 256.750 52.055 ;
        RECT 256.750 52.045 257.330 52.085 ;
        RECT 255.735 52.025 256.190 52.045 ;
        POLYGON 256.190 52.045 256.195 52.025 256.190 52.025 ;
        POLYGON 256.750 52.045 256.755 52.045 256.755 52.035 ;
        RECT 256.755 52.025 257.330 52.045 ;
        RECT 255.735 52.010 256.195 52.025 ;
        RECT 254.590 51.985 255.255 52.010 ;
        RECT 244.295 51.965 245.025 51.985 ;
        RECT 243.190 51.910 243.655 51.955 ;
        POLYGON 243.170 51.910 243.170 51.855 243.155 51.855 ;
        RECT 243.170 51.885 243.655 51.910 ;
        POLYGON 243.655 51.955 243.675 51.955 243.655 51.885 ;
        POLYGON 244.275 51.960 244.275 51.925 244.265 51.925 ;
        RECT 244.275 51.940 245.025 51.965 ;
        POLYGON 245.025 51.985 245.045 51.985 245.025 51.940 ;
        POLYGON 254.590 51.985 254.615 51.985 254.615 51.940 ;
        RECT 254.615 51.940 255.255 51.985 ;
        RECT 244.275 51.925 245.010 51.940 ;
        POLYGON 244.265 51.925 244.265 51.885 244.255 51.885 ;
        RECT 244.265 51.900 245.010 51.925 ;
        POLYGON 245.010 51.940 245.025 51.940 245.010 51.900 ;
        POLYGON 254.615 51.940 254.635 51.940 254.635 51.900 ;
        RECT 254.635 51.900 255.255 51.940 ;
        RECT 244.265 51.890 245.005 51.900 ;
        POLYGON 245.005 51.900 245.010 51.900 245.005 51.890 ;
        POLYGON 254.635 51.900 254.640 51.900 254.640 51.890 ;
        RECT 254.640 51.895 255.255 51.900 ;
        POLYGON 255.255 52.010 255.300 51.895 255.255 51.895 ;
        POLYGON 255.735 52.010 255.765 52.010 255.765 51.900 ;
        RECT 255.765 51.895 256.195 52.010 ;
        RECT 254.640 51.890 255.300 51.895 ;
        RECT 244.265 51.885 244.980 51.890 ;
        RECT 243.170 51.855 243.630 51.885 ;
        RECT 241.700 51.710 242.490 51.855 ;
        POLYGON 241.670 51.710 241.670 51.595 241.645 51.595 ;
        RECT 241.670 51.695 242.490 51.710 ;
        POLYGON 242.490 51.855 242.525 51.855 242.490 51.700 ;
        POLYGON 243.155 51.845 243.155 51.700 243.120 51.700 ;
        RECT 243.155 51.805 243.630 51.855 ;
        POLYGON 243.630 51.885 243.655 51.885 243.630 51.805 ;
        POLYGON 244.255 51.885 244.255 51.820 244.240 51.820 ;
        RECT 244.255 51.820 244.980 51.885 ;
        POLYGON 244.980 51.890 245.005 51.890 244.980 51.820 ;
        POLYGON 254.640 51.890 254.645 51.890 254.645 51.885 ;
        RECT 254.645 51.885 255.300 51.890 ;
        POLYGON 254.645 51.885 254.670 51.885 254.670 51.825 ;
        RECT 254.670 51.830 255.300 51.885 ;
        POLYGON 255.300 51.895 255.325 51.830 255.300 51.830 ;
        POLYGON 255.765 51.895 255.780 51.895 255.780 51.840 ;
        RECT 255.780 51.830 256.195 51.895 ;
        RECT 254.670 51.820 255.325 51.830 ;
        POLYGON 244.240 51.820 244.240 51.805 244.235 51.805 ;
        RECT 244.240 51.805 244.935 51.820 ;
        RECT 243.155 51.705 243.600 51.805 ;
        POLYGON 243.600 51.805 243.630 51.805 243.600 51.705 ;
        POLYGON 244.235 51.800 244.235 51.740 244.220 51.740 ;
        RECT 244.235 51.740 244.935 51.805 ;
        POLYGON 244.220 51.740 244.220 51.705 244.210 51.705 ;
        RECT 244.220 51.705 244.935 51.740 ;
        POLYGON 244.935 51.820 244.980 51.820 244.935 51.705 ;
        POLYGON 254.670 51.820 254.710 51.820 254.710 51.735 ;
        RECT 254.710 51.770 255.325 51.820 ;
        POLYGON 255.325 51.830 255.345 51.770 255.325 51.770 ;
        POLYGON 255.780 51.830 255.795 51.830 255.795 51.780 ;
        RECT 255.795 51.815 256.195 51.830 ;
        POLYGON 256.195 52.025 256.270 51.815 256.195 51.815 ;
        POLYGON 256.755 52.025 256.800 52.025 256.800 51.890 ;
        RECT 256.800 51.940 257.330 52.025 ;
        POLYGON 257.330 52.150 257.390 51.940 257.330 51.940 ;
        POLYGON 258.145 52.150 258.155 52.150 258.155 52.130 ;
        RECT 258.155 52.130 259.030 52.150 ;
        POLYGON 258.155 52.130 258.200 52.130 258.200 51.990 ;
        RECT 258.200 52.050 259.030 52.130 ;
        POLYGON 259.030 52.315 259.105 52.050 259.030 52.050 ;
        POLYGON 260.215 52.315 260.225 52.315 260.225 52.290 ;
        RECT 260.225 52.290 261.635 52.315 ;
        RECT 258.200 52.015 259.105 52.050 ;
        POLYGON 260.225 52.290 260.270 52.290 260.270 52.040 ;
        RECT 260.270 52.270 261.635 52.290 ;
        POLYGON 261.635 52.420 261.665 52.270 261.635 52.270 ;
        POLYGON 263.690 52.420 263.720 52.420 263.720 52.285 ;
        RECT 263.720 52.270 266.380 52.420 ;
        RECT 260.270 52.040 261.665 52.270 ;
        POLYGON 259.105 52.040 259.110 52.015 259.105 52.015 ;
        POLYGON 260.270 52.040 260.275 52.040 260.275 52.015 ;
        RECT 260.275 52.015 261.665 52.040 ;
        RECT 258.200 51.990 259.110 52.015 ;
        POLYGON 258.200 51.990 258.210 51.990 258.210 51.950 ;
        RECT 258.210 51.940 259.110 51.990 ;
        RECT 256.800 51.890 257.390 51.940 ;
        POLYGON 256.800 51.890 256.820 51.890 256.820 51.820 ;
        RECT 256.820 51.815 257.390 51.890 ;
        RECT 255.795 51.790 256.270 51.815 ;
        POLYGON 256.270 51.815 256.280 51.790 256.270 51.790 ;
        POLYGON 256.820 51.815 256.825 51.815 256.825 51.805 ;
        RECT 256.825 51.805 257.390 51.815 ;
        POLYGON 257.390 51.940 257.425 51.805 257.390 51.805 ;
        POLYGON 258.210 51.940 258.245 51.940 258.245 51.815 ;
        RECT 258.245 51.825 259.110 51.940 ;
        POLYGON 259.110 52.015 259.160 51.825 259.110 51.825 ;
        POLYGON 260.275 52.015 260.290 52.015 260.290 51.935 ;
        RECT 260.290 52.005 261.665 52.015 ;
        POLYGON 261.665 52.270 261.720 52.005 261.665 52.005 ;
        POLYGON 263.720 52.270 263.780 52.270 263.780 52.015 ;
        RECT 263.780 52.005 266.380 52.270 ;
        RECT 260.290 51.935 261.720 52.005 ;
        POLYGON 260.290 51.935 260.310 51.935 260.310 51.835 ;
        RECT 260.310 51.915 261.720 51.935 ;
        POLYGON 261.720 52.005 261.735 51.915 261.720 51.915 ;
        POLYGON 263.780 52.005 263.795 52.005 263.795 51.935 ;
        RECT 263.795 51.930 266.380 52.005 ;
        POLYGON 266.380 52.430 266.470 51.930 266.380 51.930 ;
        POLYGON 270.565 52.430 270.585 52.430 270.585 52.160 ;
        RECT 270.585 52.270 277.455 52.430 ;
        POLYGON 277.455 52.455 277.490 52.270 277.455 52.270 ;
        RECT 270.585 52.160 277.490 52.270 ;
        POLYGON 270.585 52.160 270.595 52.160 270.595 52.000 ;
        RECT 270.595 51.930 277.490 52.160 ;
        RECT 263.795 51.915 266.470 51.930 ;
        RECT 260.310 51.825 261.735 51.915 ;
        RECT 258.245 51.805 259.160 51.825 ;
        RECT 256.825 51.790 257.425 51.805 ;
        RECT 255.795 51.775 256.280 51.790 ;
        POLYGON 256.280 51.790 256.285 51.775 256.280 51.775 ;
        POLYGON 256.825 51.790 256.830 51.790 256.830 51.785 ;
        RECT 256.830 51.775 257.425 51.790 ;
        RECT 255.795 51.770 256.285 51.775 ;
        RECT 254.710 51.735 255.345 51.770 ;
        POLYGON 254.710 51.735 254.720 51.735 254.720 51.705 ;
        RECT 254.720 51.730 255.345 51.735 ;
        POLYGON 255.345 51.770 255.360 51.730 255.345 51.730 ;
        POLYGON 255.795 51.770 255.800 51.770 255.800 51.765 ;
        RECT 255.800 51.765 256.285 51.770 ;
        POLYGON 255.800 51.765 255.805 51.765 255.805 51.750 ;
        RECT 255.805 51.730 256.285 51.765 ;
        RECT 254.720 51.705 255.360 51.730 ;
        RECT 243.155 51.700 243.595 51.705 ;
        RECT 241.670 51.595 242.440 51.695 ;
        POLYGON 241.645 51.595 241.645 51.575 241.640 51.575 ;
        RECT 241.645 51.575 242.440 51.595 ;
        RECT 239.650 51.380 240.675 51.575 ;
        RECT 235.985 51.210 237.975 51.370 ;
        POLYGON 237.975 51.370 237.985 51.370 237.975 51.210 ;
        POLYGON 239.620 51.370 239.620 51.210 239.605 51.210 ;
        RECT 239.620 51.335 240.675 51.380 ;
        POLYGON 240.675 51.575 240.700 51.575 240.675 51.335 ;
        POLYGON 241.640 51.565 241.640 51.410 241.615 51.410 ;
        RECT 241.640 51.415 242.440 51.575 ;
        POLYGON 242.440 51.695 242.490 51.695 242.440 51.415 ;
        POLYGON 243.120 51.700 243.120 51.680 243.115 51.680 ;
        RECT 243.120 51.680 243.595 51.700 ;
        POLYGON 243.115 51.680 243.115 51.665 243.110 51.665 ;
        RECT 243.115 51.670 243.595 51.680 ;
        POLYGON 243.595 51.705 243.600 51.705 243.595 51.670 ;
        POLYGON 244.210 51.695 244.210 51.675 244.205 51.675 ;
        RECT 244.210 51.675 244.920 51.705 ;
        RECT 243.115 51.665 243.555 51.670 ;
        POLYGON 243.110 51.665 243.110 51.605 243.100 51.605 ;
        RECT 243.110 51.605 243.555 51.665 ;
        POLYGON 243.100 51.605 243.100 51.450 243.065 51.450 ;
        RECT 243.100 51.505 243.555 51.605 ;
        POLYGON 243.555 51.670 243.595 51.670 243.555 51.505 ;
        POLYGON 244.205 51.670 244.205 51.605 244.190 51.605 ;
        RECT 244.205 51.655 244.920 51.675 ;
        POLYGON 244.920 51.705 244.935 51.705 244.920 51.655 ;
        POLYGON 254.720 51.705 254.725 51.705 254.725 51.690 ;
        RECT 254.725 51.690 255.360 51.705 ;
        POLYGON 254.725 51.690 254.730 51.690 254.730 51.680 ;
        RECT 254.730 51.680 255.360 51.690 ;
        POLYGON 254.730 51.680 254.735 51.680 254.735 51.665 ;
        RECT 254.735 51.665 255.360 51.680 ;
        POLYGON 255.360 51.730 255.385 51.665 255.360 51.665 ;
        POLYGON 255.805 51.730 255.820 51.730 255.820 51.670 ;
        RECT 255.820 51.710 256.285 51.730 ;
        POLYGON 256.285 51.775 256.305 51.710 256.285 51.710 ;
        POLYGON 256.830 51.775 256.850 51.775 256.850 51.720 ;
        RECT 256.850 51.755 257.425 51.775 ;
        POLYGON 257.425 51.805 257.440 51.755 257.425 51.755 ;
        POLYGON 258.245 51.805 258.260 51.805 258.260 51.755 ;
        RECT 258.260 51.755 259.160 51.805 ;
        RECT 256.850 51.720 257.440 51.755 ;
        POLYGON 257.440 51.755 257.445 51.720 257.440 51.720 ;
        POLYGON 258.260 51.755 258.270 51.755 258.270 51.720 ;
        RECT 258.270 51.750 259.160 51.755 ;
        POLYGON 259.160 51.825 259.175 51.750 259.160 51.750 ;
        POLYGON 260.310 51.825 260.325 51.825 260.325 51.760 ;
        RECT 260.325 51.755 261.735 51.825 ;
        POLYGON 261.735 51.915 261.760 51.755 261.735 51.755 ;
        POLYGON 263.795 51.915 263.820 51.915 263.820 51.805 ;
        RECT 263.820 51.905 266.470 51.915 ;
        POLYGON 266.470 51.930 266.475 51.905 266.470 51.905 ;
        POLYGON 270.595 51.930 270.600 51.930 270.600 51.920 ;
        RECT 270.600 51.905 277.490 51.930 ;
        RECT 263.820 51.840 266.475 51.905 ;
        POLYGON 266.475 51.905 266.490 51.840 266.475 51.840 ;
        POLYGON 270.600 51.905 270.605 51.905 270.605 51.840 ;
        RECT 270.605 51.840 277.490 51.905 ;
        RECT 263.820 51.805 266.490 51.840 ;
        POLYGON 263.820 51.805 263.825 51.805 263.825 51.775 ;
        RECT 263.825 51.755 266.490 51.805 ;
        RECT 260.325 51.750 261.760 51.755 ;
        RECT 258.270 51.720 259.175 51.750 ;
        RECT 256.850 51.710 257.445 51.720 ;
        RECT 254.735 51.655 255.385 51.665 ;
        RECT 244.205 51.605 244.875 51.655 ;
        POLYGON 244.190 51.605 244.190 51.505 244.170 51.505 ;
        RECT 244.190 51.520 244.875 51.605 ;
        POLYGON 244.875 51.655 244.920 51.655 244.875 51.520 ;
        POLYGON 254.735 51.655 254.765 51.655 254.765 51.585 ;
        RECT 254.765 51.650 255.385 51.655 ;
        POLYGON 255.385 51.665 255.390 51.650 255.385 51.650 ;
        RECT 255.820 51.650 256.305 51.710 ;
        RECT 254.765 51.585 255.390 51.650 ;
        POLYGON 254.765 51.585 254.785 51.585 254.785 51.525 ;
        RECT 254.785 51.520 255.390 51.585 ;
        RECT 244.190 51.510 244.870 51.520 ;
        POLYGON 244.870 51.520 244.875 51.520 244.870 51.510 ;
        POLYGON 254.785 51.520 254.790 51.520 254.790 51.510 ;
        RECT 254.790 51.510 255.390 51.520 ;
        RECT 244.190 51.505 244.865 51.510 ;
        RECT 243.100 51.450 243.540 51.505 ;
        POLYGON 243.540 51.505 243.555 51.505 243.540 51.450 ;
        POLYGON 244.170 51.505 244.170 51.455 244.160 51.455 ;
        RECT 244.170 51.495 244.865 51.505 ;
        POLYGON 244.865 51.510 244.870 51.510 244.865 51.495 ;
        POLYGON 254.790 51.510 254.795 51.510 254.795 51.495 ;
        RECT 254.795 51.495 255.390 51.510 ;
        RECT 244.170 51.460 244.855 51.495 ;
        POLYGON 244.855 51.495 244.865 51.495 244.855 51.460 ;
        POLYGON 254.795 51.495 254.805 51.495 254.805 51.465 ;
        RECT 254.805 51.465 255.390 51.495 ;
        POLYGON 255.390 51.650 255.445 51.465 255.390 51.465 ;
        POLYGON 255.820 51.650 255.825 51.650 255.825 51.645 ;
        RECT 255.825 51.645 256.305 51.650 ;
        POLYGON 255.825 51.645 255.860 51.645 255.860 51.470 ;
        RECT 255.860 51.540 256.305 51.645 ;
        POLYGON 256.305 51.710 256.355 51.540 256.305 51.540 ;
        POLYGON 256.850 51.710 256.855 51.710 256.855 51.705 ;
        RECT 256.855 51.705 257.445 51.710 ;
        POLYGON 256.855 51.705 256.860 51.705 256.860 51.675 ;
        RECT 256.860 51.675 257.445 51.705 ;
        POLYGON 256.860 51.675 256.890 51.675 256.890 51.545 ;
        RECT 256.890 51.630 257.445 51.675 ;
        POLYGON 257.445 51.720 257.465 51.630 257.445 51.630 ;
        POLYGON 258.270 51.720 258.290 51.720 258.290 51.640 ;
        RECT 258.290 51.710 259.175 51.720 ;
        POLYGON 259.175 51.750 259.185 51.710 259.175 51.710 ;
        POLYGON 260.325 51.750 260.330 51.750 260.330 51.720 ;
        RECT 260.330 51.710 261.760 51.750 ;
        RECT 258.290 51.630 259.185 51.710 ;
        RECT 256.890 51.540 257.465 51.630 ;
        RECT 255.860 51.500 256.355 51.540 ;
        POLYGON 256.355 51.540 256.365 51.500 256.355 51.500 ;
        POLYGON 256.890 51.540 256.895 51.540 256.895 51.525 ;
        RECT 256.895 51.525 257.465 51.540 ;
        POLYGON 256.895 51.525 256.900 51.525 256.900 51.500 ;
        RECT 256.900 51.500 257.465 51.525 ;
        RECT 255.860 51.465 256.365 51.500 ;
        RECT 254.805 51.460 255.445 51.465 ;
        RECT 244.170 51.455 244.820 51.460 ;
        POLYGON 243.065 51.450 243.065 51.420 243.060 51.420 ;
        RECT 243.065 51.420 243.530 51.450 ;
        RECT 241.640 51.410 242.435 51.415 ;
        POLYGON 242.435 51.415 242.440 51.415 242.435 51.410 ;
        POLYGON 241.615 51.410 241.615 51.335 241.600 51.335 ;
        RECT 241.615 51.335 242.400 51.410 ;
        RECT 239.620 51.210 240.655 51.335 ;
        POLYGON 235.975 50.605 235.985 50.605 235.985 50.270 ;
        RECT 229.250 50.180 233.220 50.270 ;
        POLYGON 233.220 50.270 233.225 50.180 233.220 50.180 ;
        RECT 235.985 50.180 237.955 51.210 ;
        POLYGON 237.955 51.210 237.975 51.210 237.955 50.830 ;
        POLYGON 239.605 51.190 239.605 50.995 239.590 50.995 ;
        RECT 239.605 51.015 240.655 51.210 ;
        POLYGON 240.655 51.335 240.675 51.335 240.655 51.015 ;
        POLYGON 241.600 51.325 241.600 51.270 241.590 51.270 ;
        RECT 241.600 51.270 242.400 51.335 ;
        POLYGON 241.590 51.270 241.590 51.020 241.560 51.020 ;
        RECT 241.590 51.140 242.400 51.270 ;
        POLYGON 242.400 51.410 242.435 51.410 242.400 51.140 ;
        POLYGON 243.060 51.410 243.060 51.290 243.040 51.290 ;
        RECT 243.060 51.390 243.530 51.420 ;
        POLYGON 243.530 51.450 243.540 51.450 243.530 51.400 ;
        POLYGON 244.160 51.450 244.160 51.430 244.155 51.430 ;
        RECT 244.160 51.430 244.820 51.455 ;
        POLYGON 244.155 51.430 244.155 51.400 244.150 51.400 ;
        RECT 244.155 51.400 244.820 51.430 ;
        RECT 243.060 51.290 243.490 51.390 ;
        POLYGON 243.040 51.290 243.040 51.220 243.030 51.220 ;
        RECT 243.040 51.220 243.490 51.290 ;
        POLYGON 243.030 51.220 243.030 51.155 243.020 51.155 ;
        RECT 243.030 51.185 243.490 51.220 ;
        POLYGON 243.490 51.390 243.530 51.390 243.490 51.185 ;
        POLYGON 244.150 51.395 244.150 51.260 244.130 51.260 ;
        RECT 244.150 51.330 244.820 51.400 ;
        POLYGON 244.820 51.460 244.855 51.460 244.820 51.330 ;
        POLYGON 254.805 51.460 254.815 51.460 254.815 51.435 ;
        RECT 254.815 51.435 255.445 51.460 ;
        POLYGON 254.815 51.435 254.840 51.435 254.840 51.340 ;
        RECT 254.840 51.415 255.445 51.435 ;
        POLYGON 255.445 51.465 255.460 51.415 255.445 51.415 ;
        POLYGON 255.860 51.465 255.865 51.465 255.865 51.450 ;
        RECT 255.865 51.450 256.365 51.465 ;
        POLYGON 255.865 51.450 255.870 51.450 255.870 51.415 ;
        RECT 254.840 51.390 255.460 51.415 ;
        POLYGON 255.460 51.415 255.470 51.390 255.460 51.390 ;
        RECT 255.870 51.390 256.365 51.450 ;
        RECT 254.840 51.330 255.470 51.390 ;
        RECT 244.150 51.315 244.815 51.330 ;
        POLYGON 244.815 51.330 244.820 51.330 244.815 51.315 ;
        POLYGON 254.840 51.330 254.845 51.330 254.845 51.320 ;
        RECT 254.845 51.315 255.470 51.330 ;
        RECT 244.150 51.260 244.780 51.315 ;
        POLYGON 244.130 51.260 244.130 51.185 244.115 51.185 ;
        RECT 244.130 51.185 244.780 51.260 ;
        RECT 243.030 51.155 243.480 51.185 ;
        RECT 241.590 51.120 242.395 51.140 ;
        POLYGON 242.395 51.140 242.400 51.140 242.395 51.120 ;
        POLYGON 243.020 51.140 243.020 51.120 243.015 51.120 ;
        RECT 243.020 51.120 243.480 51.155 ;
        RECT 241.590 51.020 242.385 51.120 ;
        RECT 239.605 50.995 240.640 51.015 ;
        POLYGON 239.590 50.995 239.590 50.880 239.585 50.880 ;
        RECT 239.590 50.880 240.640 50.995 ;
        POLYGON 239.585 50.830 239.585 50.310 239.560 50.310 ;
        RECT 239.585 50.795 240.640 50.880 ;
        POLYGON 240.640 51.015 240.655 51.015 240.640 50.795 ;
        POLYGON 241.560 51.015 241.560 50.945 241.550 50.945 ;
        RECT 241.560 51.000 242.385 51.020 ;
        POLYGON 242.385 51.120 242.395 51.120 242.385 51.000 ;
        POLYGON 243.015 51.120 243.015 51.000 242.995 51.000 ;
        RECT 243.015 51.110 243.480 51.120 ;
        POLYGON 243.480 51.185 243.490 51.185 243.480 51.110 ;
        POLYGON 244.115 51.175 244.115 51.115 244.105 51.115 ;
        RECT 244.115 51.160 244.780 51.185 ;
        POLYGON 244.780 51.315 244.815 51.315 244.780 51.160 ;
        POLYGON 254.845 51.315 254.855 51.315 254.855 51.285 ;
        RECT 254.855 51.285 255.470 51.315 ;
        POLYGON 255.470 51.390 255.500 51.285 255.470 51.285 ;
        POLYGON 255.870 51.390 255.885 51.390 255.885 51.315 ;
        RECT 255.885 51.355 256.365 51.390 ;
        POLYGON 256.365 51.500 256.405 51.355 256.365 51.355 ;
        POLYGON 256.900 51.500 256.930 51.500 256.930 51.370 ;
        RECT 256.930 51.355 257.465 51.500 ;
        POLYGON 257.465 51.630 257.525 51.355 257.465 51.355 ;
        POLYGON 258.290 51.630 258.295 51.630 258.295 51.625 ;
        RECT 258.295 51.620 259.185 51.630 ;
        POLYGON 258.295 51.620 258.310 51.620 258.310 51.545 ;
        RECT 258.310 51.545 259.185 51.620 ;
        POLYGON 258.310 51.545 258.350 51.545 258.350 51.355 ;
        RECT 258.350 51.445 259.185 51.545 ;
        POLYGON 259.185 51.710 259.240 51.445 259.185 51.445 ;
        POLYGON 260.330 51.710 260.365 51.710 260.365 51.460 ;
        RECT 260.365 51.580 261.760 51.710 ;
        POLYGON 261.760 51.755 261.790 51.580 261.760 51.580 ;
        RECT 260.365 51.555 261.790 51.580 ;
        POLYGON 263.825 51.755 263.860 51.755 263.860 51.575 ;
        POLYGON 261.790 51.575 261.795 51.555 261.790 51.555 ;
        RECT 263.860 51.555 266.490 51.755 ;
        RECT 260.365 51.445 261.795 51.555 ;
        RECT 258.350 51.405 259.240 51.445 ;
        POLYGON 259.240 51.445 259.245 51.405 259.240 51.405 ;
        POLYGON 260.365 51.445 260.370 51.445 260.370 51.425 ;
        RECT 260.370 51.405 261.795 51.445 ;
        RECT 258.350 51.355 259.245 51.405 ;
        RECT 255.885 51.285 256.405 51.355 ;
        POLYGON 254.855 51.285 254.880 51.285 254.880 51.175 ;
        RECT 254.880 51.220 255.500 51.285 ;
        POLYGON 255.500 51.285 255.515 51.220 255.500 51.220 ;
        POLYGON 255.885 51.285 255.895 51.285 255.895 51.245 ;
        RECT 255.895 51.265 256.405 51.285 ;
        POLYGON 256.405 51.355 256.425 51.265 256.405 51.265 ;
        POLYGON 256.930 51.355 256.955 51.355 256.955 51.265 ;
        RECT 256.955 51.265 257.525 51.355 ;
        RECT 255.895 51.225 256.425 51.265 ;
        POLYGON 256.425 51.265 256.435 51.225 256.425 51.225 ;
        POLYGON 256.955 51.265 256.960 51.265 256.960 51.245 ;
        RECT 256.960 51.225 257.525 51.265 ;
        RECT 255.895 51.220 256.435 51.225 ;
        RECT 254.880 51.160 255.515 51.220 ;
        RECT 244.115 51.120 244.770 51.160 ;
        POLYGON 244.770 51.160 244.780 51.160 244.770 51.120 ;
        POLYGON 254.880 51.160 254.890 51.160 254.890 51.135 ;
        RECT 254.890 51.145 255.515 51.160 ;
        POLYGON 255.515 51.220 255.530 51.145 255.515 51.145 ;
        POLYGON 255.895 51.220 255.910 51.220 255.910 51.145 ;
        RECT 255.910 51.145 256.435 51.220 ;
        RECT 254.890 51.120 255.530 51.145 ;
        RECT 244.115 51.115 244.745 51.120 ;
        RECT 243.015 51.000 243.460 51.110 ;
        RECT 241.560 50.945 242.370 51.000 ;
        POLYGON 241.550 50.945 241.550 50.815 241.540 50.815 ;
        RECT 241.550 50.860 242.370 50.945 ;
        POLYGON 242.370 51.000 242.385 51.000 242.370 50.895 ;
        RECT 242.995 50.985 243.460 51.000 ;
        POLYGON 243.460 51.110 243.480 51.110 243.460 50.985 ;
        POLYGON 244.105 51.110 244.105 51.090 244.100 51.090 ;
        RECT 244.105 51.090 244.745 51.115 ;
        POLYGON 244.100 51.090 244.100 50.990 244.090 50.990 ;
        RECT 244.100 50.995 244.745 51.090 ;
        POLYGON 244.745 51.120 244.770 51.120 244.745 50.995 ;
        POLYGON 254.890 51.120 254.900 51.120 254.900 51.070 ;
        RECT 254.900 51.100 255.530 51.120 ;
        POLYGON 255.530 51.145 255.540 51.100 255.530 51.100 ;
        POLYGON 255.910 51.145 255.915 51.145 255.915 51.115 ;
        RECT 255.915 51.100 256.435 51.145 ;
        RECT 254.900 51.070 255.540 51.100 ;
        POLYGON 254.900 51.070 254.910 51.070 254.910 51.010 ;
        RECT 254.910 51.045 255.540 51.070 ;
        POLYGON 255.540 51.100 255.555 51.045 255.540 51.045 ;
        POLYGON 255.915 51.100 255.920 51.100 255.920 51.060 ;
        RECT 255.920 51.045 256.435 51.100 ;
        RECT 254.910 50.995 255.555 51.045 ;
        RECT 244.100 50.990 244.735 50.995 ;
        POLYGON 242.995 50.985 242.995 50.925 242.990 50.925 ;
        RECT 242.995 50.925 243.450 50.985 ;
        RECT 242.990 50.920 243.450 50.925 ;
        POLYGON 243.450 50.985 243.460 50.985 243.450 50.920 ;
        POLYGON 244.090 50.985 244.090 50.945 244.085 50.945 ;
        RECT 244.090 50.945 244.735 50.990 ;
        RECT 244.085 50.925 244.735 50.945 ;
        POLYGON 244.735 50.995 244.745 50.995 244.735 50.925 ;
        POLYGON 254.910 50.995 254.920 50.995 254.920 50.955 ;
        RECT 254.920 50.925 255.555 50.995 ;
        POLYGON 242.990 50.895 242.990 50.860 242.985 50.860 ;
        RECT 242.990 50.860 243.445 50.920 ;
        RECT 241.550 50.820 242.365 50.860 ;
        POLYGON 242.365 50.860 242.370 50.860 242.365 50.820 ;
        POLYGON 242.985 50.860 242.985 50.820 242.980 50.820 ;
        RECT 242.985 50.835 243.445 50.860 ;
        POLYGON 243.445 50.920 243.450 50.920 243.445 50.835 ;
        POLYGON 244.085 50.920 244.085 50.845 244.075 50.845 ;
        RECT 244.085 50.845 244.720 50.925 ;
        RECT 242.985 50.820 243.440 50.835 ;
        RECT 241.550 50.815 242.345 50.820 ;
        RECT 239.585 50.310 240.635 50.795 ;
        RECT 229.250 49.985 233.225 50.180 ;
        POLYGON 229.250 49.985 229.305 49.985 229.305 49.475 ;
        RECT 229.305 49.475 233.225 49.985 ;
        POLYGON 229.305 49.475 229.390 49.475 229.390 48.665 ;
        RECT 229.390 49.360 233.225 49.475 ;
        POLYGON 233.225 50.180 233.290 49.360 233.225 49.360 ;
        POLYGON 235.985 50.180 236.005 50.180 236.005 49.825 ;
        RECT 236.005 49.825 237.955 50.180 ;
        POLYGON 236.005 49.825 236.045 49.825 236.045 49.395 ;
        RECT 236.045 49.765 237.955 49.825 ;
        POLYGON 237.955 50.225 237.975 49.765 237.955 49.765 ;
        POLYGON 239.560 50.225 239.560 49.765 239.550 49.765 ;
        RECT 239.560 50.065 240.635 50.310 ;
        POLYGON 240.635 50.795 240.640 50.795 240.635 50.255 ;
        POLYGON 241.540 50.795 241.540 50.620 241.525 50.620 ;
        RECT 241.540 50.620 242.345 50.815 ;
        POLYGON 240.635 50.255 240.640 50.065 240.635 50.065 ;
        POLYGON 241.525 50.620 241.525 50.295 241.510 50.295 ;
        RECT 241.525 50.525 242.345 50.620 ;
        POLYGON 242.345 50.820 242.365 50.820 242.345 50.575 ;
        RECT 242.980 50.815 243.440 50.820 ;
        POLYGON 243.440 50.835 243.445 50.835 243.440 50.815 ;
        POLYGON 244.075 50.835 244.075 50.815 244.070 50.815 ;
        RECT 244.075 50.815 244.720 50.845 ;
        POLYGON 244.720 50.925 244.735 50.925 244.720 50.825 ;
        POLYGON 254.920 50.925 254.935 50.925 254.935 50.850 ;
        RECT 254.935 50.915 255.555 50.925 ;
        POLYGON 255.555 51.045 255.580 50.915 255.555 50.915 ;
        POLYGON 255.920 51.045 255.930 51.045 255.930 50.960 ;
        RECT 255.930 50.985 256.435 51.045 ;
        POLYGON 256.435 51.225 256.485 50.985 256.435 50.985 ;
        POLYGON 256.960 51.225 256.980 51.225 256.980 51.100 ;
        RECT 256.980 51.100 257.525 51.225 ;
        POLYGON 256.980 51.100 256.995 51.100 256.995 51.010 ;
        RECT 256.995 50.995 257.525 51.100 ;
        POLYGON 257.525 51.355 257.585 50.995 257.525 50.995 ;
        POLYGON 258.350 51.355 258.370 51.355 258.370 51.265 ;
        RECT 258.370 51.265 259.245 51.355 ;
        POLYGON 258.370 51.265 258.410 51.265 258.410 51.020 ;
        RECT 258.410 51.135 259.245 51.265 ;
        POLYGON 259.245 51.405 259.290 51.135 259.245 51.135 ;
        POLYGON 260.370 51.405 260.400 51.405 260.400 51.205 ;
        RECT 260.400 51.225 261.795 51.405 ;
        POLYGON 261.795 51.555 261.840 51.225 261.795 51.225 ;
        POLYGON 263.860 51.555 263.875 51.555 263.875 51.495 ;
        RECT 263.875 51.495 266.490 51.555 ;
        POLYGON 263.875 51.495 263.910 51.495 263.910 51.230 ;
        RECT 263.910 51.310 266.490 51.495 ;
        POLYGON 266.490 51.840 266.570 51.310 266.490 51.310 ;
        POLYGON 270.605 51.840 270.635 51.840 270.635 51.365 ;
        RECT 270.635 51.310 277.490 51.840 ;
        RECT 263.910 51.245 266.570 51.310 ;
        POLYGON 266.570 51.310 266.580 51.245 266.570 51.245 ;
        POLYGON 270.635 51.310 270.640 51.310 270.640 51.285 ;
        RECT 270.640 51.245 277.490 51.310 ;
        RECT 263.910 51.225 266.580 51.245 ;
        RECT 260.400 51.205 261.840 51.225 ;
        POLYGON 260.400 51.205 260.405 51.205 260.405 51.155 ;
        RECT 260.405 51.150 261.840 51.205 ;
        POLYGON 261.840 51.225 261.850 51.150 261.840 51.150 ;
        POLYGON 263.910 51.225 263.920 51.225 263.920 51.150 ;
        RECT 263.920 51.150 266.580 51.225 ;
        RECT 260.405 51.135 261.850 51.150 ;
        RECT 258.410 51.100 259.290 51.135 ;
        POLYGON 259.290 51.135 259.300 51.100 259.290 51.100 ;
        POLYGON 260.405 51.135 260.410 51.135 260.410 51.105 ;
        RECT 260.410 51.100 261.850 51.135 ;
        RECT 258.410 50.995 259.300 51.100 ;
        RECT 256.995 50.985 257.585 50.995 ;
        RECT 255.930 50.950 256.485 50.985 ;
        POLYGON 256.485 50.985 256.490 50.950 256.485 50.950 ;
        POLYGON 256.995 50.985 257.005 50.985 257.005 50.950 ;
        RECT 257.005 50.950 257.585 50.985 ;
        RECT 255.930 50.920 256.490 50.950 ;
        POLYGON 256.490 50.950 256.495 50.920 256.490 50.920 ;
        POLYGON 257.005 50.950 257.010 50.950 257.010 50.920 ;
        RECT 257.010 50.940 257.585 50.950 ;
        POLYGON 257.585 50.995 257.590 50.940 257.585 50.940 ;
        POLYGON 258.410 50.995 258.420 50.995 258.420 50.960 ;
        RECT 258.420 50.940 259.300 50.995 ;
        RECT 257.010 50.920 257.590 50.940 ;
        RECT 255.930 50.915 256.495 50.920 ;
        RECT 254.935 50.890 255.580 50.915 ;
        POLYGON 255.580 50.915 255.585 50.890 255.580 50.890 ;
        POLYGON 255.930 50.915 255.935 50.915 255.935 50.910 ;
        RECT 254.935 50.870 255.585 50.890 ;
        POLYGON 255.585 50.890 255.590 50.870 255.585 50.870 ;
        RECT 255.935 50.875 256.495 50.915 ;
        POLYGON 256.495 50.920 256.505 50.875 256.495 50.875 ;
        POLYGON 257.010 50.920 257.015 50.920 257.015 50.890 ;
        RECT 257.015 50.875 257.590 50.920 ;
        RECT 255.935 50.870 256.505 50.875 ;
        RECT 254.935 50.825 255.590 50.870 ;
        POLYGON 242.980 50.810 242.980 50.755 242.975 50.755 ;
        RECT 242.980 50.755 243.425 50.815 ;
        POLYGON 242.975 50.755 242.975 50.580 242.960 50.580 ;
        RECT 242.975 50.655 243.425 50.755 ;
        POLYGON 243.425 50.815 243.440 50.815 243.425 50.655 ;
        RECT 244.070 50.810 244.720 50.815 ;
        POLYGON 244.070 50.795 244.070 50.765 244.065 50.765 ;
        RECT 244.070 50.765 244.705 50.810 ;
        POLYGON 244.065 50.765 244.065 50.690 244.060 50.690 ;
        RECT 244.065 50.725 244.705 50.765 ;
        POLYGON 244.705 50.810 244.720 50.810 244.705 50.725 ;
        POLYGON 254.935 50.825 254.945 50.825 254.945 50.780 ;
        RECT 254.945 50.780 255.590 50.825 ;
        POLYGON 254.945 50.780 254.950 50.780 254.950 50.735 ;
        RECT 254.950 50.730 255.590 50.780 ;
        POLYGON 255.590 50.870 255.610 50.730 255.590 50.730 ;
        POLYGON 255.935 50.870 255.940 50.870 255.940 50.860 ;
        RECT 255.940 50.860 256.505 50.870 ;
        POLYGON 255.940 50.860 255.950 50.860 255.950 50.760 ;
        RECT 255.950 50.730 256.505 50.860 ;
        RECT 254.950 50.725 255.610 50.730 ;
        RECT 244.065 50.690 244.700 50.725 ;
        RECT 244.060 50.655 244.700 50.690 ;
        POLYGON 244.700 50.725 244.705 50.725 244.700 50.655 ;
        POLYGON 254.950 50.725 254.955 50.725 254.955 50.690 ;
        RECT 254.955 50.685 255.610 50.725 ;
        POLYGON 255.610 50.730 255.615 50.685 255.610 50.685 ;
        POLYGON 255.950 50.730 255.955 50.730 255.955 50.690 ;
        RECT 255.955 50.710 256.505 50.730 ;
        POLYGON 256.505 50.875 256.530 50.710 256.505 50.710 ;
        POLYGON 257.015 50.875 257.030 50.875 257.030 50.805 ;
        RECT 257.030 50.805 257.590 50.875 ;
        POLYGON 257.030 50.805 257.035 50.805 257.035 50.750 ;
        RECT 257.035 50.710 257.590 50.805 ;
        RECT 255.955 50.685 256.530 50.710 ;
        RECT 254.955 50.655 255.615 50.685 ;
        RECT 242.975 50.580 243.420 50.655 ;
        RECT 241.525 50.295 242.335 50.525 ;
        POLYGON 242.335 50.525 242.345 50.525 242.335 50.295 ;
        POLYGON 242.960 50.575 242.960 50.520 242.955 50.520 ;
        RECT 242.960 50.540 243.420 50.580 ;
        POLYGON 243.420 50.655 243.425 50.655 243.420 50.540 ;
        POLYGON 244.060 50.655 244.060 50.540 244.050 50.540 ;
        RECT 244.060 50.540 244.690 50.655 ;
        RECT 242.960 50.520 243.410 50.540 ;
        POLYGON 242.955 50.520 242.955 50.295 242.950 50.295 ;
        RECT 242.955 50.295 243.410 50.520 ;
        POLYGON 243.410 50.540 243.420 50.540 243.410 50.385 ;
        POLYGON 244.050 50.540 244.050 50.465 244.045 50.465 ;
        RECT 244.050 50.490 244.690 50.540 ;
        POLYGON 244.690 50.655 244.700 50.655 244.690 50.530 ;
        POLYGON 254.955 50.655 254.970 50.655 254.970 50.560 ;
        RECT 254.970 50.560 255.615 50.655 ;
        POLYGON 255.615 50.685 255.635 50.560 255.615 50.560 ;
        POLYGON 255.955 50.685 255.960 50.685 255.960 50.620 ;
        RECT 255.960 50.620 256.530 50.685 ;
        RECT 254.970 50.530 255.635 50.560 ;
        POLYGON 255.960 50.620 255.965 50.620 255.965 50.545 ;
        RECT 244.050 50.465 244.685 50.490 ;
        RECT 241.510 50.065 242.335 50.295 ;
        RECT 239.560 49.765 240.640 50.065 ;
        RECT 236.045 49.670 237.975 49.765 ;
        POLYGON 237.975 49.765 237.985 49.670 237.975 49.670 ;
        RECT 239.550 49.715 240.640 49.765 ;
        POLYGON 240.640 50.065 240.655 49.715 240.640 49.715 ;
        POLYGON 241.510 50.065 241.515 50.065 241.515 49.965 ;
        RECT 241.515 49.965 242.335 50.065 ;
        POLYGON 242.950 50.285 242.950 50.055 242.945 50.055 ;
        POLYGON 242.945 50.055 242.950 50.055 242.950 50.020 ;
        RECT 242.950 50.015 243.410 50.295 ;
        POLYGON 244.045 50.385 244.045 50.130 244.040 50.130 ;
        RECT 244.045 50.130 244.685 50.465 ;
        POLYGON 244.685 50.490 244.690 50.490 244.685 50.335 ;
        POLYGON 254.970 50.530 254.985 50.530 254.985 50.435 ;
        RECT 254.985 50.510 255.635 50.530 ;
        POLYGON 255.635 50.545 255.640 50.510 255.635 50.510 ;
        RECT 255.965 50.510 256.530 50.620 ;
        RECT 254.985 50.435 255.640 50.510 ;
        RECT 244.040 50.115 244.685 50.130 ;
        POLYGON 244.685 50.335 244.690 50.115 244.685 50.115 ;
        POLYGON 254.985 50.435 255.000 50.435 255.000 50.170 ;
        RECT 255.000 50.360 255.640 50.435 ;
        POLYGON 255.640 50.510 255.655 50.360 255.640 50.360 ;
        POLYGON 255.965 50.510 255.975 50.510 255.975 50.395 ;
        RECT 255.975 50.430 256.530 50.510 ;
        POLYGON 256.530 50.710 256.565 50.430 256.530 50.430 ;
        POLYGON 257.035 50.710 257.060 50.710 257.060 50.480 ;
        RECT 257.060 50.665 257.590 50.710 ;
        POLYGON 257.590 50.940 257.625 50.665 257.590 50.665 ;
        POLYGON 258.420 50.940 258.430 50.940 258.430 50.900 ;
        RECT 258.430 50.900 259.300 50.940 ;
        POLYGON 258.430 50.900 258.445 50.900 258.445 50.785 ;
        RECT 258.445 50.820 259.300 50.900 ;
        POLYGON 259.300 51.100 259.335 50.820 259.300 50.820 ;
        POLYGON 260.410 51.100 260.420 51.100 260.420 51.005 ;
        RECT 260.420 51.005 261.850 51.100 ;
        POLYGON 260.420 51.005 260.440 51.005 260.440 50.820 ;
        RECT 260.440 50.845 261.850 51.005 ;
        POLYGON 261.850 51.150 261.880 50.845 261.850 50.845 ;
        POLYGON 263.920 51.150 263.945 51.150 263.945 50.965 ;
        RECT 263.945 50.965 266.580 51.150 ;
        POLYGON 263.945 50.965 263.955 50.965 263.955 50.865 ;
        RECT 263.955 50.845 266.580 50.965 ;
        RECT 258.445 50.790 259.335 50.820 ;
        POLYGON 259.335 50.820 259.340 50.790 259.335 50.790 ;
        RECT 260.440 50.790 261.880 50.845 ;
        RECT 258.445 50.785 259.340 50.790 ;
        RECT 257.060 50.555 257.625 50.665 ;
        POLYGON 258.445 50.785 258.460 50.785 258.460 50.655 ;
        RECT 258.460 50.655 259.340 50.785 ;
        POLYGON 257.625 50.655 257.635 50.555 257.625 50.555 ;
        POLYGON 258.460 50.655 258.465 50.655 258.465 50.595 ;
        RECT 258.465 50.555 259.340 50.655 ;
        RECT 257.060 50.510 257.635 50.555 ;
        POLYGON 257.635 50.555 257.640 50.510 257.635 50.510 ;
        POLYGON 258.465 50.555 258.470 50.555 258.470 50.535 ;
        RECT 258.470 50.510 259.340 50.555 ;
        POLYGON 259.340 50.790 259.365 50.510 259.340 50.510 ;
        POLYGON 260.440 50.790 260.460 50.790 260.460 50.640 ;
        RECT 260.460 50.640 261.880 50.790 ;
        POLYGON 260.460 50.640 260.465 50.640 260.465 50.545 ;
        RECT 260.465 50.520 261.880 50.640 ;
        POLYGON 261.880 50.845 261.910 50.520 261.880 50.520 ;
        POLYGON 263.955 50.845 263.990 50.845 263.990 50.530 ;
        RECT 263.990 50.710 266.580 50.845 ;
        POLYGON 266.580 51.245 266.645 50.710 266.580 50.710 ;
        POLYGON 270.640 51.245 270.660 51.245 270.660 50.970 ;
        RECT 270.660 51.220 277.490 51.245 ;
        POLYGON 277.490 52.270 277.650 51.220 277.490 51.220 ;
        POLYGON 287.935 52.270 287.935 51.515 287.930 51.515 ;
        RECT 287.935 51.515 303.120 58.190 ;
        RECT 270.660 51.210 277.650 51.220 ;
        POLYGON 277.650 51.220 277.655 51.210 277.650 51.210 ;
        RECT 270.660 51.070 277.655 51.210 ;
        POLYGON 277.655 51.210 277.670 51.070 277.655 51.070 ;
        RECT 270.660 50.710 277.670 51.070 ;
        RECT 263.990 50.520 266.645 50.710 ;
        RECT 257.060 50.480 257.640 50.510 ;
        RECT 255.000 50.175 255.655 50.360 ;
        POLYGON 255.655 50.330 255.665 50.175 255.655 50.175 ;
        POLYGON 241.515 49.965 241.525 49.965 241.525 49.730 ;
        RECT 241.525 49.730 242.335 49.965 ;
        POLYGON 242.335 50.015 242.345 49.730 242.335 49.730 ;
        POLYGON 242.950 50.015 242.955 50.015 242.955 49.820 ;
        RECT 242.955 49.835 243.410 50.015 ;
        POLYGON 243.410 50.035 243.420 49.835 243.410 49.835 ;
        RECT 244.040 49.890 244.690 50.115 ;
        RECT 255.000 50.125 255.665 50.175 ;
        POLYGON 255.665 50.175 255.670 50.125 255.665 50.125 ;
        RECT 255.975 50.140 256.565 50.430 ;
        POLYGON 257.060 50.480 257.065 50.480 257.065 50.420 ;
        RECT 257.065 50.390 257.640 50.480 ;
        POLYGON 256.565 50.390 256.585 50.140 256.565 50.140 ;
        POLYGON 257.065 50.390 257.070 50.390 257.070 50.365 ;
        RECT 257.070 50.365 257.640 50.390 ;
        POLYGON 257.070 50.365 257.075 50.365 257.075 50.215 ;
        RECT 257.075 50.300 257.640 50.365 ;
        POLYGON 257.640 50.510 257.655 50.300 257.640 50.300 ;
        POLYGON 258.470 50.510 258.485 50.510 258.485 50.315 ;
        RECT 258.485 50.500 259.365 50.510 ;
        POLYGON 259.365 50.510 259.370 50.500 259.365 50.500 ;
        RECT 258.485 50.300 259.370 50.500 ;
        RECT 260.465 50.480 261.910 50.520 ;
        RECT 255.975 50.125 256.585 50.140 ;
        POLYGON 244.690 50.095 244.700 49.890 244.690 49.890 ;
        RECT 255.000 49.995 255.670 50.125 ;
        POLYGON 255.670 50.125 255.675 49.995 255.670 49.995 ;
        POLYGON 255.975 50.125 255.980 50.125 255.980 50.025 ;
        RECT 244.040 49.835 244.700 49.890 ;
        RECT 241.525 49.715 242.345 49.730 ;
        RECT 239.550 49.670 240.655 49.715 ;
        RECT 236.045 49.360 237.985 49.670 ;
        RECT 229.390 49.270 233.290 49.360 ;
        POLYGON 233.290 49.360 233.305 49.270 233.290 49.270 ;
        POLYGON 236.045 49.360 236.055 49.360 236.055 49.280 ;
        RECT 236.055 49.270 237.985 49.360 ;
        RECT 207.230 48.615 222.360 48.655 ;
        RECT 229.390 48.635 233.305 49.270 ;
        POLYGON 207.230 48.615 207.310 48.615 207.310 48.300 ;
        RECT 207.310 48.300 222.360 48.615 ;
        POLYGON 207.310 48.300 207.630 48.300 207.630 47.030 ;
        RECT 207.630 47.875 222.360 48.300 ;
        POLYGON 222.360 48.635 222.455 47.875 222.360 47.875 ;
        POLYGON 229.390 48.635 229.395 48.635 229.395 48.620 ;
        RECT 229.395 48.620 233.305 48.635 ;
        POLYGON 229.395 48.620 229.485 48.620 229.485 48.090 ;
        RECT 229.485 48.445 233.305 48.620 ;
        POLYGON 233.305 49.270 233.415 48.445 233.305 48.445 ;
        POLYGON 236.055 49.270 236.075 49.270 236.075 49.050 ;
        RECT 236.075 49.235 237.985 49.270 ;
        POLYGON 237.985 49.670 238.020 49.235 237.985 49.235 ;
        POLYGON 239.550 49.670 239.560 49.670 239.560 49.510 ;
        RECT 239.560 49.510 240.655 49.670 ;
        POLYGON 239.560 49.510 239.565 49.510 239.565 49.335 ;
        RECT 239.565 49.495 240.655 49.510 ;
        POLYGON 240.655 49.715 240.675 49.495 240.655 49.495 ;
        POLYGON 241.525 49.715 241.530 49.715 241.530 49.645 ;
        RECT 241.530 49.645 242.345 49.715 ;
        RECT 242.955 49.770 243.420 49.835 ;
        POLYGON 242.955 49.770 242.960 49.770 242.960 49.705 ;
        RECT 242.960 49.765 243.420 49.770 ;
        POLYGON 243.420 49.835 243.425 49.765 243.420 49.765 ;
        POLYGON 244.040 49.835 244.045 49.835 244.045 49.805 ;
        RECT 244.045 49.825 244.700 49.835 ;
        POLYGON 244.700 49.890 244.705 49.825 244.700 49.825 ;
        RECT 244.045 49.765 244.705 49.825 ;
        RECT 242.960 49.705 243.425 49.765 ;
        POLYGON 241.530 49.645 241.540 49.645 241.540 49.525 ;
        RECT 241.540 49.495 242.345 49.645 ;
        RECT 239.565 49.235 240.675 49.495 ;
        RECT 236.075 49.125 238.020 49.235 ;
        POLYGON 238.020 49.235 238.035 49.125 238.020 49.125 ;
        POLYGON 239.565 49.235 239.570 49.235 239.570 49.165 ;
        RECT 239.570 49.180 240.675 49.235 ;
        POLYGON 240.675 49.495 240.700 49.180 240.675 49.180 ;
        POLYGON 241.540 49.495 241.550 49.495 241.550 49.405 ;
        RECT 241.550 49.450 242.345 49.495 ;
        POLYGON 242.345 49.705 242.365 49.450 242.345 49.450 ;
        POLYGON 242.960 49.705 242.970 49.705 242.970 49.585 ;
        RECT 242.970 49.585 243.425 49.705 ;
        POLYGON 242.970 49.585 242.975 49.585 242.975 49.535 ;
        RECT 242.975 49.580 243.425 49.585 ;
        POLYGON 243.425 49.765 243.440 49.580 243.425 49.580 ;
        POLYGON 244.045 49.765 244.060 49.765 244.060 49.610 ;
        RECT 244.060 49.700 244.705 49.765 ;
        POLYGON 244.705 49.825 244.720 49.700 244.705 49.700 ;
        RECT 255.000 49.810 255.675 49.995 ;
        RECT 242.975 49.555 243.440 49.580 ;
        POLYGON 243.440 49.580 243.445 49.555 243.440 49.555 ;
        RECT 244.060 49.570 244.720 49.700 ;
        POLYGON 255.000 49.725 255.000 49.675 254.995 49.675 ;
        RECT 255.000 49.675 255.670 49.810 ;
        POLYGON 244.720 49.675 244.735 49.570 244.720 49.570 ;
        POLYGON 254.995 49.665 254.995 49.605 254.990 49.605 ;
        RECT 254.995 49.625 255.670 49.675 ;
        POLYGON 255.670 49.810 255.675 49.810 255.670 49.625 ;
        RECT 254.995 49.605 255.655 49.625 ;
        RECT 244.060 49.555 244.735 49.570 ;
        RECT 242.975 49.535 243.445 49.555 ;
        POLYGON 242.975 49.535 242.980 49.535 242.980 49.475 ;
        RECT 242.980 49.490 243.445 49.535 ;
        POLYGON 243.445 49.555 243.450 49.490 243.445 49.490 ;
        POLYGON 244.060 49.555 244.065 49.555 244.065 49.545 ;
        RECT 244.065 49.490 244.735 49.555 ;
        RECT 242.980 49.450 243.450 49.490 ;
        RECT 241.550 49.420 242.365 49.450 ;
        POLYGON 242.365 49.450 242.370 49.420 242.365 49.420 ;
        RECT 241.550 49.405 242.370 49.420 ;
        POLYGON 242.980 49.450 242.985 49.450 242.985 49.415 ;
        POLYGON 241.550 49.405 241.560 49.405 241.560 49.320 ;
        RECT 241.560 49.315 242.370 49.405 ;
        RECT 242.985 49.385 243.450 49.450 ;
        POLYGON 241.560 49.315 241.575 49.315 241.575 49.210 ;
        RECT 241.575 49.285 242.370 49.315 ;
        POLYGON 242.370 49.385 242.385 49.285 242.370 49.285 ;
        POLYGON 242.985 49.385 242.990 49.385 242.990 49.355 ;
        RECT 242.990 49.355 243.450 49.385 ;
        POLYGON 242.990 49.355 242.995 49.355 242.995 49.300 ;
        RECT 242.995 49.285 243.450 49.355 ;
        RECT 241.575 49.180 242.385 49.285 ;
        RECT 239.570 49.125 240.700 49.180 ;
        RECT 236.075 49.050 238.035 49.125 ;
        POLYGON 236.075 49.050 236.145 49.050 236.145 48.600 ;
        RECT 236.145 48.710 238.035 49.050 ;
        POLYGON 238.035 49.125 238.090 48.710 238.035 48.710 ;
        POLYGON 239.570 49.125 239.590 49.125 239.590 48.975 ;
        RECT 239.590 48.975 240.700 49.125 ;
        POLYGON 239.590 48.975 239.610 48.975 239.610 48.730 ;
        RECT 239.610 48.940 240.700 48.975 ;
        POLYGON 240.700 49.180 240.735 48.940 240.700 48.940 ;
        POLYGON 241.575 49.180 241.590 49.180 241.590 49.105 ;
        RECT 241.590 49.170 242.385 49.180 ;
        POLYGON 242.385 49.285 242.395 49.170 242.385 49.170 ;
        POLYGON 242.995 49.285 243.010 49.285 243.010 49.195 ;
        RECT 243.010 49.280 243.450 49.285 ;
        POLYGON 243.450 49.490 243.480 49.280 243.450 49.280 ;
        POLYGON 244.065 49.490 244.070 49.490 244.070 49.485 ;
        RECT 244.070 49.475 244.735 49.490 ;
        POLYGON 244.070 49.475 244.085 49.475 244.085 49.325 ;
        RECT 244.085 49.460 244.735 49.475 ;
        POLYGON 244.735 49.570 244.745 49.460 244.735 49.460 ;
        POLYGON 254.990 49.570 254.990 49.460 254.980 49.460 ;
        RECT 254.990 49.460 255.655 49.605 ;
        RECT 244.085 49.315 244.745 49.460 ;
        POLYGON 244.745 49.460 244.770 49.315 244.745 49.315 ;
        POLYGON 254.980 49.445 254.980 49.330 254.965 49.330 ;
        RECT 254.980 49.435 255.655 49.460 ;
        POLYGON 255.655 49.625 255.670 49.625 255.655 49.445 ;
        POLYGON 255.980 49.625 255.980 49.550 255.975 49.550 ;
        RECT 255.980 49.550 256.585 50.125 ;
        RECT 257.075 50.110 257.655 50.300 ;
        POLYGON 256.585 50.110 256.590 49.830 256.585 49.830 ;
        POLYGON 255.975 49.550 255.975 49.460 255.970 49.460 ;
        RECT 255.975 49.545 256.585 49.550 ;
        POLYGON 256.585 49.830 256.590 49.830 256.585 49.545 ;
        POLYGON 257.075 50.110 257.085 50.110 257.085 49.925 ;
        RECT 257.085 50.070 257.655 50.110 ;
        POLYGON 257.655 50.300 257.670 50.070 257.655 50.070 ;
        POLYGON 258.485 50.300 258.495 50.300 258.495 50.170 ;
        RECT 258.495 50.265 259.370 50.300 ;
        POLYGON 259.370 50.480 259.385 50.265 259.370 50.265 ;
        POLYGON 260.465 50.480 260.475 50.480 260.475 50.355 ;
        RECT 260.475 50.280 261.910 50.480 ;
        POLYGON 261.910 50.520 261.930 50.280 261.910 50.280 ;
        POLYGON 263.990 50.520 264.000 50.520 264.000 50.435 ;
        RECT 264.000 50.435 266.645 50.520 ;
        POLYGON 264.000 50.435 264.010 50.435 264.010 50.280 ;
        RECT 260.475 50.265 261.930 50.280 ;
        RECT 264.010 50.265 266.645 50.435 ;
        RECT 258.495 50.200 259.385 50.265 ;
        POLYGON 259.385 50.265 259.390 50.200 259.385 50.200 ;
        POLYGON 260.475 50.265 260.480 50.265 260.480 50.260 ;
        RECT 258.495 50.170 259.390 50.200 ;
        RECT 260.480 50.170 261.930 50.265 ;
        POLYGON 257.085 49.925 257.085 49.545 257.075 49.545 ;
        RECT 257.085 49.545 257.670 50.070 ;
        POLYGON 258.495 50.170 258.500 50.170 258.500 49.985 ;
        RECT 258.500 49.920 259.390 50.170 ;
        POLYGON 257.670 49.920 257.680 49.620 257.670 49.620 ;
        POLYGON 258.500 49.920 258.505 49.920 258.505 49.805 ;
        RECT 258.505 49.890 259.390 49.920 ;
        POLYGON 259.390 50.170 259.400 49.890 259.390 49.890 ;
        POLYGON 260.480 50.170 260.490 50.170 260.490 50.070 ;
        RECT 255.975 49.460 256.565 49.545 ;
        RECT 254.980 49.330 255.640 49.435 ;
        RECT 244.085 49.280 244.770 49.315 ;
        RECT 243.010 49.220 243.480 49.280 ;
        POLYGON 243.480 49.280 243.490 49.220 243.480 49.220 ;
        POLYGON 244.085 49.280 244.095 49.280 244.095 49.225 ;
        RECT 244.095 49.250 244.770 49.280 ;
        POLYGON 244.770 49.315 244.780 49.250 244.770 49.250 ;
        POLYGON 254.965 49.315 254.965 49.290 254.960 49.290 ;
        RECT 254.965 49.290 255.640 49.330 ;
        POLYGON 254.960 49.290 254.960 49.260 254.955 49.260 ;
        RECT 254.960 49.265 255.640 49.290 ;
        POLYGON 255.640 49.435 255.655 49.435 255.640 49.265 ;
        POLYGON 255.970 49.445 255.970 49.275 255.960 49.275 ;
        RECT 255.970 49.275 256.565 49.460 ;
        RECT 255.960 49.265 256.565 49.275 ;
        POLYGON 256.565 49.545 256.585 49.545 256.565 49.265 ;
        POLYGON 257.075 49.480 257.075 49.410 257.070 49.410 ;
        RECT 257.075 49.410 257.670 49.545 ;
        POLYGON 257.070 49.410 257.070 49.285 257.060 49.285 ;
        RECT 257.070 49.320 257.670 49.410 ;
        POLYGON 257.670 49.620 257.680 49.620 257.670 49.320 ;
        POLYGON 258.505 49.805 258.505 49.480 258.495 49.480 ;
        RECT 258.505 49.545 259.400 49.890 ;
        RECT 258.505 49.480 259.390 49.545 ;
        POLYGON 258.495 49.440 258.495 49.320 258.485 49.320 ;
        RECT 258.495 49.320 259.390 49.480 ;
        RECT 257.070 49.285 257.655 49.320 ;
        RECT 254.960 49.260 255.590 49.265 ;
        RECT 244.095 49.220 244.780 49.250 ;
        RECT 243.010 49.170 243.490 49.220 ;
        RECT 241.590 49.155 242.395 49.170 ;
        POLYGON 242.395 49.170 242.400 49.155 242.395 49.155 ;
        POLYGON 243.010 49.170 243.015 49.170 243.015 49.160 ;
        RECT 243.015 49.155 243.490 49.170 ;
        RECT 241.590 49.105 242.400 49.155 ;
        POLYGON 241.590 49.105 241.610 49.105 241.610 48.970 ;
        RECT 241.610 48.940 242.400 49.105 ;
        RECT 239.610 48.795 240.735 48.940 ;
        POLYGON 240.735 48.940 240.755 48.795 240.735 48.795 ;
        POLYGON 241.610 48.940 241.630 48.940 241.630 48.835 ;
        RECT 241.630 48.890 242.400 48.940 ;
        POLYGON 242.400 49.155 242.435 48.890 242.400 48.890 ;
        POLYGON 243.015 49.155 243.020 49.155 243.020 49.125 ;
        RECT 243.020 49.125 243.490 49.155 ;
        POLYGON 243.020 49.125 243.030 49.125 243.030 49.075 ;
        RECT 243.030 49.075 243.490 49.125 ;
        POLYGON 243.030 49.075 243.055 49.075 243.055 48.895 ;
        RECT 243.055 48.995 243.490 49.075 ;
        POLYGON 243.490 49.220 243.530 48.995 243.490 48.995 ;
        POLYGON 244.095 49.220 244.100 49.220 244.100 49.180 ;
        RECT 244.100 49.180 244.780 49.220 ;
        POLYGON 244.100 49.180 244.105 49.180 244.105 49.170 ;
        RECT 243.055 48.890 243.530 48.995 ;
        RECT 244.105 49.155 244.780 49.180 ;
        POLYGON 244.105 49.155 244.130 49.155 244.130 48.990 ;
        RECT 244.130 49.070 244.780 49.155 ;
        POLYGON 244.780 49.250 244.815 49.070 244.780 49.070 ;
        POLYGON 254.955 49.250 254.955 49.200 254.945 49.200 ;
        RECT 254.955 49.200 255.590 49.260 ;
        POLYGON 254.945 49.200 254.945 49.070 254.925 49.070 ;
        RECT 254.945 49.070 255.590 49.200 ;
        RECT 244.130 49.045 244.815 49.070 ;
        POLYGON 244.815 49.070 244.820 49.045 244.815 49.045 ;
        POLYGON 254.925 49.070 254.925 49.045 254.920 49.045 ;
        RECT 254.925 49.045 255.590 49.070 ;
        RECT 244.130 48.990 244.820 49.045 ;
        POLYGON 243.530 48.990 243.555 48.890 243.530 48.890 ;
        POLYGON 244.130 48.990 244.145 48.990 244.145 48.895 ;
        RECT 244.145 48.890 244.820 48.990 ;
        POLYGON 244.820 49.045 244.855 48.890 244.820 48.890 ;
        POLYGON 254.920 49.035 254.920 48.980 254.910 48.980 ;
        RECT 254.920 48.980 255.590 49.045 ;
        POLYGON 254.910 48.980 254.910 48.940 254.900 48.940 ;
        RECT 254.910 48.940 255.590 48.980 ;
        POLYGON 254.900 48.940 254.900 48.890 254.890 48.890 ;
        RECT 254.900 48.905 255.590 48.940 ;
        POLYGON 255.590 49.265 255.640 49.265 255.590 48.905 ;
        POLYGON 255.960 49.265 255.960 49.170 255.950 49.170 ;
        RECT 255.960 49.170 256.530 49.265 ;
        POLYGON 255.950 49.170 255.950 49.050 255.940 49.050 ;
        RECT 255.950 49.050 256.530 49.170 ;
        POLYGON 255.940 49.050 255.940 48.910 255.930 48.910 ;
        RECT 255.940 48.985 256.530 49.050 ;
        POLYGON 256.530 49.265 256.565 49.265 256.530 48.985 ;
        POLYGON 257.060 49.265 257.060 49.040 257.040 49.040 ;
        RECT 257.060 49.040 257.655 49.285 ;
        POLYGON 257.040 49.040 257.040 49.005 257.035 49.005 ;
        RECT 257.040 49.020 257.655 49.040 ;
        POLYGON 257.655 49.320 257.670 49.320 257.655 49.020 ;
        POLYGON 258.485 49.300 258.485 49.095 258.470 49.095 ;
        RECT 258.485 49.235 259.390 49.320 ;
        POLYGON 259.390 49.545 259.400 49.545 259.390 49.235 ;
        RECT 260.490 50.005 261.930 50.170 ;
        POLYGON 260.490 50.005 260.500 50.005 260.500 49.490 ;
        RECT 260.500 49.515 261.930 50.005 ;
        POLYGON 261.930 50.265 261.955 49.515 261.930 49.515 ;
        POLYGON 264.010 50.265 264.035 50.265 264.035 49.900 ;
        RECT 264.035 50.050 266.645 50.265 ;
        POLYGON 266.645 50.710 266.700 50.050 266.645 50.050 ;
        POLYGON 270.660 50.710 270.670 50.710 270.670 50.230 ;
        RECT 270.670 50.125 277.670 50.710 ;
        POLYGON 277.670 51.070 277.775 50.125 277.670 50.125 ;
        RECT 270.670 50.050 277.775 50.125 ;
        RECT 264.035 49.900 266.700 50.050 ;
        POLYGON 264.035 49.900 264.045 49.900 264.045 49.540 ;
        RECT 264.045 49.515 266.700 49.900 ;
        POLYGON 260.500 49.490 260.500 49.235 260.490 49.235 ;
        RECT 260.500 49.235 261.955 49.515 ;
        POLYGON 261.955 49.515 261.960 49.355 261.955 49.355 ;
        RECT 258.485 49.095 259.370 49.235 ;
        POLYGON 258.470 49.080 258.470 49.025 258.465 49.025 ;
        RECT 258.470 49.025 259.370 49.095 ;
        RECT 257.040 49.005 257.625 49.020 ;
        RECT 255.940 48.910 256.505 48.985 ;
        RECT 254.900 48.890 255.555 48.905 ;
        RECT 241.630 48.885 242.435 48.890 ;
        POLYGON 242.435 48.890 242.440 48.885 242.435 48.885 ;
        RECT 243.055 48.885 243.555 48.890 ;
        RECT 241.630 48.835 242.440 48.885 ;
        RECT 239.610 48.710 240.755 48.795 ;
        POLYGON 241.630 48.835 241.640 48.835 241.640 48.790 ;
        RECT 241.640 48.780 242.440 48.835 ;
        RECT 236.145 48.600 238.090 48.710 ;
        POLYGON 236.145 48.600 236.165 48.600 236.165 48.470 ;
        RECT 236.165 48.585 238.090 48.600 ;
        POLYGON 238.090 48.710 238.110 48.585 238.090 48.585 ;
        POLYGON 239.610 48.710 239.615 48.710 239.615 48.670 ;
        RECT 239.615 48.670 240.755 48.710 ;
        POLYGON 239.615 48.670 239.625 48.670 239.625 48.600 ;
        RECT 239.625 48.650 240.755 48.670 ;
        POLYGON 240.755 48.780 240.775 48.650 240.755 48.650 ;
        POLYGON 241.640 48.780 241.645 48.780 241.645 48.770 ;
        RECT 241.645 48.770 242.440 48.780 ;
        POLYGON 241.645 48.770 241.665 48.770 241.665 48.670 ;
        RECT 241.665 48.650 242.440 48.770 ;
        RECT 239.625 48.585 240.775 48.650 ;
        RECT 236.165 48.445 238.110 48.585 ;
        POLYGON 238.110 48.585 238.135 48.445 238.110 48.445 ;
        POLYGON 239.625 48.585 239.645 48.585 239.645 48.465 ;
        RECT 239.645 48.445 240.775 48.585 ;
        RECT 229.485 48.375 233.415 48.445 ;
        POLYGON 233.415 48.445 233.430 48.375 233.415 48.375 ;
        POLYGON 236.165 48.445 236.180 48.445 236.180 48.375 ;
        RECT 236.180 48.375 238.135 48.445 ;
        RECT 229.485 48.140 233.430 48.375 ;
        POLYGON 233.430 48.375 233.475 48.140 233.430 48.140 ;
        POLYGON 236.180 48.375 236.195 48.375 236.195 48.280 ;
        RECT 236.195 48.280 238.135 48.375 ;
        POLYGON 236.195 48.280 236.220 48.280 236.220 48.160 ;
        RECT 236.220 48.190 238.135 48.280 ;
        POLYGON 238.135 48.445 238.180 48.190 238.135 48.190 ;
        POLYGON 239.645 48.445 239.650 48.445 239.650 48.435 ;
        RECT 239.650 48.435 240.775 48.445 ;
        POLYGON 239.650 48.435 239.655 48.435 239.655 48.430 ;
        RECT 239.655 48.415 240.775 48.435 ;
        POLYGON 240.775 48.650 240.820 48.415 240.775 48.415 ;
        POLYGON 241.665 48.650 241.710 48.650 241.710 48.450 ;
        RECT 241.710 48.615 242.440 48.650 ;
        POLYGON 242.440 48.885 242.490 48.615 242.440 48.615 ;
        POLYGON 243.055 48.885 243.065 48.885 243.065 48.845 ;
        RECT 243.065 48.845 243.555 48.885 ;
        POLYGON 243.065 48.845 243.100 48.845 243.100 48.665 ;
        RECT 243.100 48.715 243.555 48.845 ;
        POLYGON 243.555 48.890 243.595 48.715 243.555 48.715 ;
        POLYGON 244.145 48.890 244.150 48.890 244.150 48.865 ;
        RECT 244.150 48.865 244.855 48.890 ;
        POLYGON 244.150 48.865 244.155 48.865 244.155 48.850 ;
        RECT 244.155 48.850 244.855 48.865 ;
        POLYGON 244.155 48.850 244.180 48.850 244.180 48.730 ;
        RECT 244.180 48.845 244.855 48.850 ;
        POLYGON 244.855 48.890 244.865 48.845 244.855 48.845 ;
        POLYGON 254.890 48.890 254.890 48.850 254.880 48.850 ;
        RECT 254.890 48.850 255.555 48.890 ;
        RECT 244.180 48.830 244.865 48.845 ;
        POLYGON 244.865 48.845 244.870 48.830 244.865 48.830 ;
        POLYGON 254.880 48.845 254.880 48.830 254.875 48.830 ;
        RECT 254.880 48.830 255.555 48.850 ;
        RECT 244.180 48.820 244.870 48.830 ;
        POLYGON 244.870 48.830 244.875 48.820 244.870 48.820 ;
        POLYGON 254.875 48.830 254.875 48.820 254.870 48.820 ;
        RECT 254.875 48.820 255.555 48.830 ;
        RECT 244.180 48.715 244.875 48.820 ;
        RECT 243.100 48.685 243.595 48.715 ;
        POLYGON 243.595 48.715 243.600 48.685 243.595 48.685 ;
        POLYGON 244.180 48.715 244.185 48.715 244.185 48.705 ;
        RECT 244.185 48.685 244.875 48.715 ;
        RECT 243.100 48.665 243.600 48.685 ;
        POLYGON 243.100 48.665 243.110 48.665 243.110 48.625 ;
        RECT 243.110 48.625 243.600 48.665 ;
        POLYGON 243.110 48.625 243.115 48.625 243.115 48.615 ;
        RECT 241.710 48.455 242.490 48.615 ;
        RECT 243.115 48.610 243.600 48.625 ;
        POLYGON 242.490 48.610 242.525 48.455 242.490 48.455 ;
        POLYGON 243.115 48.610 243.150 48.610 243.150 48.460 ;
        RECT 243.150 48.580 243.600 48.610 ;
        POLYGON 243.600 48.685 243.630 48.580 243.600 48.580 ;
        POLYGON 244.185 48.685 244.210 48.685 244.210 48.585 ;
        RECT 244.210 48.650 244.875 48.685 ;
        POLYGON 244.875 48.820 244.920 48.650 244.875 48.650 ;
        POLYGON 254.870 48.815 254.870 48.760 254.855 48.760 ;
        RECT 254.870 48.760 255.555 48.820 ;
        POLYGON 254.855 48.760 254.855 48.680 254.835 48.680 ;
        RECT 254.855 48.725 255.555 48.760 ;
        POLYGON 255.555 48.905 255.590 48.905 255.555 48.725 ;
        POLYGON 255.930 48.905 255.930 48.730 255.905 48.730 ;
        RECT 255.930 48.825 256.505 48.910 ;
        POLYGON 256.505 48.985 256.530 48.985 256.505 48.825 ;
        POLYGON 257.035 48.985 257.035 48.965 257.030 48.965 ;
        RECT 257.035 48.965 257.625 49.005 ;
        POLYGON 257.030 48.965 257.030 48.835 257.010 48.835 ;
        RECT 257.030 48.835 257.625 48.965 ;
        RECT 255.930 48.730 256.485 48.825 ;
        RECT 254.855 48.680 255.520 48.725 ;
        POLYGON 254.835 48.680 254.835 48.650 254.825 48.650 ;
        RECT 254.835 48.650 255.520 48.680 ;
        RECT 244.210 48.595 244.920 48.650 ;
        POLYGON 244.920 48.650 244.935 48.595 244.920 48.595 ;
        POLYGON 254.825 48.650 254.825 48.615 254.815 48.615 ;
        RECT 254.825 48.615 255.520 48.650 ;
        POLYGON 254.815 48.610 254.815 48.595 254.810 48.595 ;
        RECT 254.815 48.595 255.520 48.615 ;
        RECT 244.210 48.580 244.935 48.595 ;
        RECT 243.150 48.500 243.630 48.580 ;
        POLYGON 243.630 48.580 243.655 48.500 243.630 48.500 ;
        POLYGON 244.210 48.580 244.220 48.580 244.220 48.550 ;
        RECT 244.220 48.550 244.935 48.580 ;
        POLYGON 244.220 48.550 244.230 48.550 244.230 48.510 ;
        RECT 244.230 48.500 244.935 48.550 ;
        RECT 243.150 48.455 243.655 48.500 ;
        RECT 241.710 48.450 242.525 48.455 ;
        POLYGON 241.710 48.450 241.715 48.450 241.715 48.425 ;
        RECT 241.715 48.415 242.525 48.450 ;
        RECT 239.655 48.410 240.820 48.415 ;
        POLYGON 239.655 48.410 239.695 48.410 239.695 48.195 ;
        RECT 239.695 48.190 240.820 48.410 ;
        RECT 236.220 48.155 238.180 48.190 ;
        POLYGON 238.180 48.190 238.190 48.155 238.180 48.155 ;
        POLYGON 239.695 48.190 239.700 48.190 239.700 48.170 ;
        RECT 239.700 48.155 240.820 48.190 ;
        RECT 236.220 48.140 238.190 48.155 ;
        RECT 229.485 48.090 233.475 48.140 ;
        POLYGON 229.485 48.090 229.520 48.090 229.520 47.875 ;
        RECT 207.630 47.150 222.455 47.875 ;
        RECT 229.520 47.865 233.475 48.090 ;
        POLYGON 222.455 47.865 222.585 47.150 222.455 47.150 ;
        POLYGON 229.520 47.865 229.620 47.865 229.620 47.275 ;
        RECT 229.620 47.535 233.475 47.865 ;
        POLYGON 233.475 48.140 233.590 47.535 233.475 47.535 ;
        POLYGON 236.220 48.140 236.295 48.140 236.295 47.810 ;
        RECT 236.295 48.045 238.190 48.140 ;
        POLYGON 238.190 48.155 238.215 48.045 238.190 48.045 ;
        POLYGON 239.700 48.155 239.725 48.155 239.725 48.050 ;
        RECT 239.725 48.135 240.820 48.155 ;
        POLYGON 240.820 48.415 240.870 48.135 240.820 48.135 ;
        POLYGON 241.715 48.415 241.730 48.415 241.730 48.365 ;
        RECT 241.730 48.365 242.525 48.415 ;
        POLYGON 241.730 48.365 241.790 48.365 241.790 48.140 ;
        RECT 241.790 48.345 242.525 48.365 ;
        POLYGON 242.525 48.455 242.550 48.345 242.525 48.345 ;
        POLYGON 243.150 48.455 243.155 48.455 243.155 48.440 ;
        RECT 243.155 48.440 243.655 48.455 ;
        POLYGON 243.155 48.440 243.170 48.440 243.170 48.385 ;
        RECT 243.170 48.430 243.655 48.440 ;
        POLYGON 243.655 48.500 243.675 48.430 243.655 48.430 ;
        POLYGON 244.230 48.500 244.240 48.500 244.240 48.470 ;
        RECT 244.240 48.470 244.935 48.500 ;
        POLYGON 244.240 48.470 244.250 48.470 244.250 48.430 ;
        RECT 244.250 48.455 244.935 48.470 ;
        POLYGON 244.935 48.595 244.980 48.455 244.935 48.455 ;
        POLYGON 254.810 48.595 254.810 48.530 254.790 48.530 ;
        RECT 254.810 48.575 255.520 48.595 ;
        POLYGON 255.520 48.725 255.555 48.725 255.520 48.575 ;
        POLYGON 255.905 48.725 255.905 48.590 255.885 48.590 ;
        RECT 255.905 48.705 256.485 48.730 ;
        POLYGON 256.485 48.825 256.505 48.825 256.485 48.705 ;
        POLYGON 257.010 48.825 257.010 48.705 256.990 48.705 ;
        RECT 257.010 48.720 257.625 48.835 ;
        POLYGON 257.625 49.020 257.655 49.020 257.625 48.725 ;
        POLYGON 258.465 49.020 258.465 48.965 258.460 48.965 ;
        RECT 258.465 48.965 259.370 49.025 ;
        POLYGON 258.460 48.965 258.460 48.830 258.445 48.830 ;
        RECT 258.460 48.940 259.370 48.965 ;
        POLYGON 259.370 49.235 259.390 49.235 259.370 48.940 ;
        POLYGON 260.490 49.120 260.490 48.940 260.485 48.940 ;
        RECT 260.490 48.940 261.955 49.235 ;
        RECT 258.460 48.925 259.365 48.940 ;
        POLYGON 259.365 48.940 259.370 48.940 259.365 48.925 ;
        RECT 258.460 48.830 259.335 48.925 ;
        POLYGON 258.445 48.830 258.445 48.725 258.430 48.725 ;
        RECT 258.445 48.725 259.335 48.830 ;
        RECT 257.010 48.705 257.610 48.720 ;
        RECT 255.905 48.590 256.425 48.705 ;
        RECT 254.810 48.550 255.515 48.575 ;
        POLYGON 255.515 48.575 255.520 48.575 255.515 48.550 ;
        POLYGON 255.885 48.575 255.885 48.555 255.880 48.555 ;
        RECT 255.885 48.555 256.425 48.590 ;
        RECT 254.810 48.530 255.495 48.550 ;
        POLYGON 254.790 48.530 254.790 48.455 254.765 48.455 ;
        RECT 254.790 48.475 255.495 48.530 ;
        POLYGON 255.495 48.550 255.515 48.550 255.495 48.475 ;
        POLYGON 255.880 48.550 255.880 48.485 255.870 48.485 ;
        RECT 255.880 48.485 256.425 48.555 ;
        RECT 254.790 48.455 255.470 48.475 ;
        RECT 243.170 48.385 243.675 48.430 ;
        RECT 244.250 48.425 244.980 48.455 ;
        POLYGON 243.170 48.385 243.180 48.385 243.180 48.345 ;
        RECT 241.790 48.135 242.550 48.345 ;
        RECT 243.180 48.330 243.675 48.385 ;
        RECT 239.725 48.045 240.870 48.135 ;
        RECT 236.295 47.810 238.215 48.045 ;
        POLYGON 236.295 47.810 236.350 47.810 236.350 47.540 ;
        RECT 236.350 47.675 238.215 47.810 ;
        POLYGON 238.215 48.045 238.295 47.675 238.215 47.675 ;
        POLYGON 239.725 48.045 239.745 48.045 239.745 47.960 ;
        RECT 239.745 47.960 240.870 48.045 ;
        POLYGON 239.745 47.960 239.760 47.960 239.760 47.915 ;
        RECT 239.760 47.915 240.870 47.960 ;
        POLYGON 239.760 47.915 239.805 47.915 239.805 47.725 ;
        RECT 239.805 47.895 240.870 47.915 ;
        POLYGON 240.870 48.135 240.930 47.895 240.870 47.895 ;
        POLYGON 241.790 48.135 241.855 48.135 241.855 47.900 ;
        RECT 241.855 48.130 242.550 48.135 ;
        POLYGON 242.550 48.330 242.605 48.130 242.550 48.130 ;
        POLYGON 243.180 48.330 243.215 48.330 243.215 48.215 ;
        RECT 243.215 48.235 243.675 48.330 ;
        POLYGON 243.675 48.425 243.735 48.235 243.675 48.235 ;
        POLYGON 244.250 48.425 244.290 48.425 244.290 48.275 ;
        RECT 244.290 48.380 244.980 48.425 ;
        POLYGON 244.980 48.455 245.005 48.380 244.980 48.380 ;
        POLYGON 254.765 48.455 254.765 48.385 254.740 48.385 ;
        RECT 254.765 48.385 255.470 48.455 ;
        RECT 244.290 48.375 245.005 48.380 ;
        POLYGON 245.005 48.380 245.010 48.375 245.005 48.375 ;
        POLYGON 254.740 48.380 254.740 48.375 254.735 48.375 ;
        RECT 254.740 48.375 255.470 48.385 ;
        POLYGON 255.470 48.475 255.495 48.475 255.470 48.375 ;
        POLYGON 255.870 48.475 255.870 48.375 255.850 48.375 ;
        RECT 255.870 48.430 256.425 48.485 ;
        POLYGON 256.425 48.705 256.485 48.705 256.425 48.430 ;
        POLYGON 256.990 48.700 256.990 48.635 256.980 48.635 ;
        RECT 256.990 48.635 257.610 48.705 ;
        POLYGON 256.980 48.635 256.980 48.600 256.975 48.600 ;
        RECT 256.980 48.610 257.610 48.635 ;
        POLYGON 257.610 48.720 257.625 48.720 257.610 48.610 ;
        POLYGON 258.430 48.715 258.430 48.620 258.415 48.620 ;
        RECT 258.430 48.620 259.335 48.725 ;
        RECT 258.415 48.615 259.335 48.620 ;
        POLYGON 259.335 48.925 259.365 48.925 259.335 48.615 ;
        POLYGON 260.485 48.915 260.485 48.615 260.465 48.615 ;
        RECT 260.485 48.615 261.955 48.940 ;
        RECT 256.980 48.600 257.585 48.610 ;
        POLYGON 256.975 48.600 256.975 48.515 256.960 48.515 ;
        RECT 256.975 48.515 257.585 48.600 ;
        POLYGON 256.960 48.515 256.960 48.430 256.940 48.430 ;
        RECT 256.960 48.435 257.585 48.515 ;
        POLYGON 257.585 48.610 257.610 48.610 257.585 48.435 ;
        POLYGON 258.415 48.610 258.415 48.435 258.385 48.435 ;
        RECT 258.415 48.435 259.290 48.615 ;
        RECT 256.960 48.430 257.530 48.435 ;
        RECT 255.870 48.375 256.410 48.430 ;
        POLYGON 256.410 48.430 256.425 48.430 256.410 48.375 ;
        POLYGON 256.940 48.420 256.940 48.375 256.930 48.375 ;
        RECT 256.940 48.375 257.530 48.430 ;
        RECT 244.290 48.320 245.010 48.375 ;
        POLYGON 245.010 48.375 245.025 48.320 245.010 48.320 ;
        POLYGON 254.735 48.370 254.735 48.355 254.730 48.355 ;
        RECT 254.735 48.355 255.360 48.375 ;
        POLYGON 254.730 48.355 254.730 48.345 254.725 48.345 ;
        RECT 254.730 48.345 255.360 48.355 ;
        POLYGON 254.725 48.345 254.725 48.330 254.720 48.330 ;
        RECT 254.725 48.330 255.360 48.345 ;
        RECT 244.290 48.275 245.025 48.320 ;
        POLYGON 244.290 48.275 244.300 48.275 244.300 48.235 ;
        RECT 244.300 48.265 245.025 48.275 ;
        POLYGON 245.025 48.320 245.045 48.265 245.025 48.265 ;
        POLYGON 254.720 48.320 254.720 48.270 254.700 48.270 ;
        RECT 254.720 48.270 255.360 48.330 ;
        RECT 244.300 48.235 245.045 48.265 ;
        RECT 243.215 48.215 243.735 48.235 ;
        POLYGON 243.215 48.215 243.230 48.215 243.230 48.165 ;
        RECT 243.230 48.165 243.735 48.215 ;
        POLYGON 243.230 48.165 243.240 48.165 243.240 48.130 ;
        RECT 243.240 48.145 243.735 48.165 ;
        POLYGON 243.735 48.235 243.765 48.145 243.735 48.145 ;
        POLYGON 244.300 48.235 244.330 48.235 244.330 48.145 ;
        RECT 244.330 48.150 245.045 48.235 ;
        POLYGON 245.045 48.265 245.090 48.150 245.045 48.150 ;
        POLYGON 254.700 48.265 254.700 48.240 254.690 48.240 ;
        RECT 254.700 48.240 255.360 48.270 ;
        POLYGON 254.690 48.240 254.690 48.155 254.655 48.155 ;
        RECT 254.690 48.155 255.360 48.240 ;
        RECT 244.330 48.145 245.090 48.150 ;
        RECT 243.240 48.130 243.765 48.145 ;
        RECT 241.855 48.085 242.605 48.130 ;
        POLYGON 242.605 48.130 242.615 48.085 242.605 48.085 ;
        POLYGON 243.240 48.130 243.255 48.130 243.255 48.085 ;
        RECT 243.255 48.085 243.765 48.130 ;
        RECT 241.855 48.055 242.615 48.085 ;
        POLYGON 242.615 48.085 242.625 48.055 242.615 48.055 ;
        POLYGON 243.255 48.085 243.260 48.085 243.260 48.065 ;
        RECT 243.260 48.055 243.765 48.085 ;
        RECT 241.855 47.895 242.625 48.055 ;
        RECT 239.805 47.725 240.930 47.895 ;
        POLYGON 239.805 47.725 239.820 47.725 239.820 47.680 ;
        RECT 239.820 47.675 240.930 47.725 ;
        RECT 236.350 47.535 238.295 47.675 ;
        RECT 229.620 47.400 233.590 47.535 ;
        POLYGON 233.590 47.535 233.620 47.400 233.590 47.400 ;
        POLYGON 236.350 47.535 236.355 47.535 236.355 47.520 ;
        RECT 236.355 47.520 238.295 47.535 ;
        POLYGON 236.355 47.520 236.385 47.520 236.385 47.405 ;
        RECT 236.385 47.510 238.295 47.520 ;
        POLYGON 238.295 47.675 238.340 47.510 238.295 47.510 ;
        POLYGON 239.820 47.675 239.830 47.675 239.830 47.655 ;
        RECT 239.830 47.655 240.930 47.675 ;
        POLYGON 239.830 47.655 239.870 47.655 239.870 47.515 ;
        RECT 239.870 47.630 240.930 47.655 ;
        POLYGON 240.930 47.895 240.995 47.630 240.930 47.630 ;
        POLYGON 241.855 47.895 241.865 47.895 241.865 47.875 ;
        RECT 241.865 47.875 242.625 47.895 ;
        POLYGON 241.865 47.875 241.885 47.875 241.885 47.825 ;
        RECT 241.885 47.860 242.625 47.875 ;
        POLYGON 242.625 48.055 242.685 47.860 242.625 47.860 ;
        POLYGON 243.260 48.055 243.285 48.055 243.285 47.990 ;
        RECT 243.285 47.990 243.765 48.055 ;
        POLYGON 243.285 47.990 243.300 47.990 243.300 47.940 ;
        RECT 243.300 47.940 243.765 47.990 ;
        POLYGON 243.300 47.940 243.325 47.940 243.325 47.865 ;
        RECT 243.325 47.915 243.765 47.940 ;
        POLYGON 243.765 48.145 243.850 47.915 243.765 47.915 ;
        POLYGON 244.330 48.145 244.380 48.145 244.380 47.990 ;
        RECT 244.380 48.080 245.090 48.145 ;
        POLYGON 245.090 48.150 245.115 48.080 245.090 48.080 ;
        POLYGON 254.655 48.150 254.655 48.130 254.645 48.130 ;
        RECT 254.655 48.130 255.360 48.155 ;
        POLYGON 254.645 48.130 254.645 48.105 254.630 48.105 ;
        RECT 254.645 48.105 255.360 48.130 ;
        POLYGON 254.630 48.095 254.630 48.085 254.625 48.085 ;
        RECT 254.630 48.085 255.360 48.105 ;
        RECT 244.380 47.990 245.115 48.080 ;
        POLYGON 244.380 47.990 244.385 47.990 244.385 47.975 ;
        RECT 244.385 47.970 245.115 47.990 ;
        POLYGON 245.115 48.080 245.165 47.970 245.115 47.970 ;
        POLYGON 254.625 48.080 254.625 47.970 254.570 47.970 ;
        RECT 254.625 48.030 255.360 48.085 ;
        POLYGON 255.360 48.375 255.470 48.375 255.360 48.030 ;
        POLYGON 255.850 48.365 255.850 48.225 255.825 48.225 ;
        RECT 255.850 48.225 256.355 48.375 ;
        POLYGON 255.825 48.210 255.825 48.125 255.805 48.125 ;
        RECT 255.825 48.155 256.355 48.225 ;
        POLYGON 256.355 48.375 256.410 48.375 256.355 48.155 ;
        POLYGON 256.930 48.375 256.930 48.210 256.895 48.210 ;
        RECT 256.930 48.210 257.530 48.375 ;
        POLYGON 256.895 48.210 256.895 48.165 256.885 48.165 ;
        RECT 256.895 48.165 257.530 48.210 ;
        POLYGON 256.885 48.165 256.885 48.155 256.880 48.155 ;
        RECT 256.885 48.155 257.530 48.165 ;
        RECT 255.825 48.125 256.280 48.155 ;
        POLYGON 255.805 48.125 255.805 48.115 255.800 48.115 ;
        RECT 255.805 48.115 256.280 48.125 ;
        POLYGON 255.800 48.115 255.800 48.030 255.780 48.030 ;
        RECT 255.800 48.030 256.280 48.115 ;
        RECT 254.625 47.990 255.345 48.030 ;
        POLYGON 255.345 48.030 255.360 48.030 255.345 47.990 ;
        POLYGON 255.780 48.025 255.780 47.990 255.770 47.990 ;
        RECT 255.780 47.990 256.280 48.030 ;
        RECT 254.625 47.970 255.320 47.990 ;
        POLYGON 244.385 47.970 244.405 47.970 244.405 47.915 ;
        RECT 244.405 47.935 245.165 47.970 ;
        POLYGON 245.165 47.970 245.180 47.935 245.165 47.935 ;
        POLYGON 254.570 47.970 254.570 47.955 254.565 47.955 ;
        RECT 254.570 47.955 255.320 47.970 ;
        POLYGON 254.565 47.955 254.565 47.935 254.555 47.935 ;
        RECT 254.565 47.935 255.320 47.955 ;
        RECT 244.405 47.915 245.180 47.935 ;
        RECT 243.325 47.860 243.850 47.915 ;
        RECT 241.885 47.830 242.685 47.860 ;
        POLYGON 242.685 47.860 242.695 47.830 242.685 47.830 ;
        POLYGON 243.325 47.860 243.335 47.860 243.335 47.840 ;
        RECT 243.335 47.855 243.850 47.860 ;
        POLYGON 243.850 47.915 243.875 47.855 243.850 47.855 ;
        POLYGON 244.405 47.915 244.425 47.915 244.425 47.860 ;
        RECT 244.425 47.910 245.180 47.915 ;
        POLYGON 245.180 47.935 245.190 47.910 245.180 47.910 ;
        POLYGON 254.555 47.935 254.555 47.915 254.545 47.915 ;
        RECT 254.555 47.920 255.320 47.935 ;
        POLYGON 255.320 47.990 255.345 47.990 255.320 47.920 ;
        POLYGON 255.770 47.980 255.770 47.920 255.755 47.920 ;
        RECT 255.770 47.920 256.280 47.990 ;
        RECT 254.555 47.915 255.235 47.920 ;
        RECT 244.425 47.900 245.190 47.910 ;
        POLYGON 245.190 47.910 245.195 47.900 245.190 47.900 ;
        POLYGON 254.545 47.910 254.545 47.905 254.540 47.905 ;
        RECT 254.545 47.905 255.235 47.915 ;
        RECT 243.335 47.830 243.875 47.855 ;
        RECT 244.425 47.850 245.195 47.900 ;
        RECT 241.885 47.825 242.695 47.830 ;
        POLYGON 241.885 47.825 241.950 47.825 241.950 47.630 ;
        RECT 241.950 47.780 242.695 47.825 ;
        POLYGON 242.695 47.830 242.710 47.780 242.695 47.780 ;
        POLYGON 243.335 47.830 243.355 47.830 243.355 47.780 ;
        RECT 243.355 47.780 243.875 47.830 ;
        RECT 241.950 47.630 242.710 47.780 ;
        RECT 239.870 47.610 240.995 47.630 ;
        POLYGON 240.995 47.630 241.005 47.610 240.995 47.610 ;
        POLYGON 241.950 47.630 241.955 47.630 241.955 47.615 ;
        RECT 241.955 47.610 242.710 47.630 ;
        RECT 239.870 47.510 241.005 47.610 ;
        RECT 236.385 47.400 238.340 47.510 ;
        RECT 229.620 47.275 233.620 47.400 ;
        POLYGON 229.620 47.275 229.645 47.275 229.645 47.160 ;
        RECT 207.630 47.030 222.585 47.150 ;
        RECT 229.645 47.140 233.620 47.275 ;
        POLYGON 222.585 47.140 222.610 47.030 222.585 47.030 ;
        POLYGON 229.645 47.140 229.670 47.140 229.670 47.045 ;
        RECT 229.670 47.040 233.620 47.140 ;
        POLYGON 233.620 47.400 233.710 47.040 233.620 47.040 ;
        POLYGON 236.385 47.400 236.390 47.400 236.390 47.390 ;
        RECT 236.390 47.390 238.340 47.400 ;
        RECT 229.670 47.030 233.710 47.040 ;
        POLYGON 236.390 47.390 236.485 47.390 236.485 47.035 ;
        RECT 236.485 47.170 238.340 47.390 ;
        POLYGON 238.340 47.510 238.435 47.170 238.340 47.170 ;
        POLYGON 239.870 47.510 239.905 47.510 239.905 47.395 ;
        RECT 239.905 47.400 241.005 47.510 ;
        POLYGON 241.005 47.610 241.070 47.400 241.005 47.400 ;
        POLYGON 241.955 47.610 241.990 47.610 241.990 47.510 ;
        RECT 241.990 47.575 242.710 47.610 ;
        POLYGON 242.710 47.780 242.780 47.575 242.710 47.575 ;
        POLYGON 243.355 47.780 243.360 47.780 243.360 47.770 ;
        RECT 243.360 47.770 243.875 47.780 ;
        POLYGON 243.360 47.770 243.375 47.770 243.375 47.720 ;
        RECT 243.375 47.720 243.875 47.770 ;
        POLYGON 243.375 47.720 243.395 47.720 243.395 47.670 ;
        RECT 243.395 47.670 243.875 47.720 ;
        POLYGON 243.395 47.670 243.430 47.670 243.430 47.575 ;
        RECT 243.430 47.625 243.875 47.670 ;
        POLYGON 243.875 47.850 243.975 47.625 243.875 47.625 ;
        POLYGON 244.425 47.850 244.480 47.850 244.480 47.715 ;
        RECT 244.480 47.725 245.195 47.850 ;
        POLYGON 245.195 47.900 245.280 47.725 245.195 47.725 ;
        POLYGON 254.540 47.900 254.540 47.885 254.530 47.885 ;
        RECT 254.540 47.885 255.235 47.905 ;
        POLYGON 254.530 47.885 254.530 47.880 254.525 47.880 ;
        RECT 254.530 47.880 255.235 47.885 ;
        POLYGON 254.525 47.880 254.525 47.815 254.495 47.815 ;
        RECT 254.525 47.815 255.235 47.880 ;
        POLYGON 254.495 47.815 254.495 47.810 254.490 47.810 ;
        RECT 254.495 47.810 255.235 47.815 ;
        POLYGON 254.490 47.810 254.490 47.725 254.445 47.725 ;
        RECT 254.490 47.725 255.235 47.810 ;
        RECT 244.480 47.715 245.280 47.725 ;
        POLYGON 244.480 47.715 244.490 47.715 244.490 47.690 ;
        RECT 244.490 47.690 245.280 47.715 ;
        POLYGON 244.490 47.690 244.515 47.690 244.515 47.625 ;
        RECT 244.515 47.625 245.280 47.690 ;
        RECT 243.430 47.575 243.975 47.625 ;
        RECT 241.990 47.510 242.780 47.575 ;
        POLYGON 242.780 47.575 242.805 47.510 242.780 47.510 ;
        POLYGON 243.430 47.575 243.440 47.575 243.440 47.550 ;
        RECT 243.440 47.570 243.975 47.575 ;
        POLYGON 243.975 47.625 243.995 47.570 243.975 47.570 ;
        POLYGON 244.515 47.625 244.535 47.625 244.535 47.580 ;
        RECT 244.535 47.615 245.280 47.625 ;
        POLYGON 245.280 47.725 245.335 47.615 245.280 47.615 ;
        POLYGON 254.445 47.725 254.445 47.680 254.420 47.680 ;
        RECT 254.445 47.690 255.235 47.725 ;
        POLYGON 255.235 47.920 255.320 47.920 255.235 47.690 ;
        POLYGON 255.755 47.915 255.755 47.890 255.750 47.890 ;
        RECT 255.755 47.910 256.280 47.920 ;
        POLYGON 256.280 48.155 256.355 48.155 256.280 47.910 ;
        RECT 256.880 48.145 257.530 48.155 ;
        POLYGON 257.530 48.435 257.585 48.435 257.530 48.145 ;
        POLYGON 258.385 48.430 258.385 48.365 258.375 48.365 ;
        RECT 258.385 48.365 259.290 48.435 ;
        POLYGON 258.375 48.365 258.375 48.345 258.370 48.345 ;
        RECT 258.375 48.345 259.290 48.365 ;
        POLYGON 258.370 48.345 258.370 48.150 258.330 48.150 ;
        RECT 258.370 48.305 259.290 48.345 ;
        POLYGON 259.290 48.615 259.335 48.615 259.290 48.305 ;
        POLYGON 260.465 48.590 260.465 48.510 260.460 48.510 ;
        RECT 260.465 48.525 261.955 48.615 ;
        POLYGON 261.955 49.355 261.960 49.355 261.955 48.525 ;
        POLYGON 264.045 49.515 264.050 49.515 264.050 49.365 ;
        RECT 264.050 49.510 266.700 49.515 ;
        POLYGON 266.700 50.050 266.725 49.510 266.700 49.510 ;
        POLYGON 270.670 50.050 270.675 50.050 270.675 49.860 ;
        RECT 270.675 49.910 277.775 50.050 ;
        POLYGON 277.775 50.125 277.795 49.910 277.775 49.910 ;
        RECT 270.675 49.510 277.795 49.910 ;
        RECT 264.050 49.450 266.725 49.510 ;
        POLYGON 266.725 49.510 266.730 49.450 266.725 49.450 ;
        POLYGON 270.675 49.510 270.680 49.510 270.680 49.490 ;
        RECT 270.680 49.450 277.795 49.510 ;
        POLYGON 264.050 49.365 264.050 48.830 264.045 48.830 ;
        RECT 264.050 48.845 266.730 49.450 ;
        POLYGON 266.730 49.450 266.740 48.845 266.730 48.845 ;
        RECT 264.050 48.830 266.725 48.845 ;
        POLYGON 264.045 48.830 264.045 48.580 264.035 48.580 ;
        RECT 264.045 48.580 266.725 48.830 ;
        RECT 260.465 48.510 261.950 48.525 ;
        POLYGON 260.460 48.510 260.460 48.345 260.445 48.345 ;
        RECT 260.460 48.465 261.950 48.510 ;
        POLYGON 261.950 48.525 261.955 48.525 261.950 48.465 ;
        POLYGON 264.035 48.525 264.035 48.465 264.030 48.465 ;
        RECT 264.035 48.465 266.725 48.580 ;
        RECT 260.460 48.345 261.930 48.465 ;
        POLYGON 260.445 48.345 260.445 48.305 260.440 48.305 ;
        RECT 260.445 48.305 261.930 48.345 ;
        RECT 258.370 48.150 259.240 48.305 ;
        POLYGON 256.880 48.145 256.880 48.075 256.860 48.075 ;
        RECT 256.880 48.075 257.465 48.145 ;
        POLYGON 256.860 48.075 256.860 48.045 256.855 48.045 ;
        RECT 256.860 48.045 257.465 48.075 ;
        POLYGON 256.855 48.045 256.855 47.910 256.815 47.910 ;
        RECT 256.855 47.910 257.465 48.045 ;
        RECT 255.755 47.890 256.270 47.910 ;
        POLYGON 255.750 47.890 255.750 47.795 255.725 47.795 ;
        RECT 255.750 47.880 256.270 47.890 ;
        POLYGON 256.270 47.910 256.280 47.910 256.270 47.880 ;
        POLYGON 256.815 47.905 256.815 47.880 256.805 47.880 ;
        RECT 256.815 47.880 257.465 47.910 ;
        RECT 255.750 47.810 256.245 47.880 ;
        POLYGON 256.245 47.880 256.270 47.880 256.245 47.810 ;
        POLYGON 256.805 47.870 256.805 47.855 256.800 47.855 ;
        RECT 256.805 47.855 257.465 47.880 ;
        POLYGON 257.465 48.145 257.530 48.145 257.465 47.855 ;
        POLYGON 258.330 48.145 258.330 48.050 258.310 48.050 ;
        RECT 258.330 48.050 259.240 48.150 ;
        POLYGON 258.310 48.050 258.310 48.010 258.305 48.010 ;
        RECT 258.310 48.010 259.240 48.050 ;
        POLYGON 258.305 48.010 258.305 47.985 258.295 47.985 ;
        RECT 258.305 47.995 259.240 48.010 ;
        POLYGON 259.240 48.305 259.290 48.305 259.240 47.995 ;
        POLYGON 260.440 48.300 260.440 48.120 260.420 48.120 ;
        RECT 260.440 48.120 261.930 48.305 ;
        POLYGON 260.420 48.120 260.420 47.995 260.405 47.995 ;
        RECT 260.420 47.995 261.930 48.120 ;
        RECT 258.305 47.985 259.175 47.995 ;
        POLYGON 258.295 47.975 258.295 47.855 258.265 47.855 ;
        RECT 258.295 47.855 259.175 47.985 ;
        POLYGON 256.800 47.855 256.800 47.815 256.790 47.815 ;
        RECT 256.800 47.815 257.425 47.855 ;
        RECT 255.750 47.795 256.175 47.810 ;
        POLYGON 255.725 47.795 255.725 47.735 255.710 47.735 ;
        RECT 255.725 47.735 256.175 47.795 ;
        POLYGON 255.710 47.735 255.710 47.690 255.695 47.690 ;
        RECT 255.710 47.690 256.175 47.735 ;
        RECT 254.445 47.680 255.160 47.690 ;
        POLYGON 254.420 47.680 254.420 47.655 254.405 47.655 ;
        RECT 254.420 47.655 255.160 47.680 ;
        POLYGON 254.405 47.655 254.405 47.615 254.380 47.615 ;
        RECT 254.405 47.615 255.160 47.655 ;
        RECT 244.535 47.570 245.335 47.615 ;
        RECT 243.440 47.565 243.995 47.570 ;
        POLYGON 243.995 47.570 244.000 47.565 243.995 47.565 ;
        POLYGON 244.535 47.570 244.540 47.570 244.540 47.565 ;
        RECT 244.540 47.565 245.335 47.570 ;
        RECT 243.440 47.550 244.000 47.565 ;
        POLYGON 243.440 47.550 243.455 47.550 243.455 47.515 ;
        RECT 243.455 47.510 244.000 47.550 ;
        POLYGON 241.990 47.510 242.010 47.510 242.010 47.450 ;
        RECT 242.010 47.450 242.805 47.510 ;
        POLYGON 242.010 47.450 242.030 47.450 242.030 47.400 ;
        RECT 242.030 47.400 242.805 47.450 ;
        POLYGON 242.805 47.510 242.850 47.400 242.805 47.400 ;
        POLYGON 243.455 47.510 243.460 47.510 243.460 47.505 ;
        RECT 243.460 47.505 244.000 47.510 ;
        POLYGON 243.460 47.505 243.500 47.505 243.500 47.405 ;
        RECT 243.500 47.480 244.000 47.505 ;
        POLYGON 244.000 47.565 244.040 47.480 244.000 47.480 ;
        POLYGON 244.540 47.565 244.575 47.565 244.575 47.490 ;
        RECT 244.575 47.560 245.335 47.565 ;
        POLYGON 245.335 47.615 245.365 47.560 245.335 47.560 ;
        POLYGON 254.380 47.610 254.380 47.560 254.350 47.560 ;
        RECT 254.380 47.560 255.160 47.615 ;
        RECT 244.575 47.555 245.365 47.560 ;
        POLYGON 245.365 47.560 245.370 47.555 245.365 47.555 ;
        RECT 244.575 47.525 245.370 47.555 ;
        POLYGON 245.370 47.555 245.385 47.525 245.370 47.525 ;
        POLYGON 254.350 47.555 254.350 47.525 254.330 47.525 ;
        RECT 254.350 47.535 255.160 47.560 ;
        POLYGON 255.160 47.690 255.235 47.690 255.160 47.535 ;
        POLYGON 255.695 47.690 255.695 47.645 255.680 47.645 ;
        RECT 255.695 47.645 256.175 47.690 ;
        POLYGON 255.680 47.640 255.680 47.610 255.670 47.610 ;
        RECT 255.680 47.610 256.175 47.645 ;
        POLYGON 256.175 47.810 256.245 47.810 256.175 47.610 ;
        POLYGON 256.790 47.810 256.790 47.740 256.770 47.740 ;
        RECT 256.790 47.740 257.425 47.815 ;
        POLYGON 256.770 47.740 256.770 47.635 256.735 47.635 ;
        RECT 256.770 47.705 257.425 47.740 ;
        POLYGON 257.425 47.855 257.465 47.855 257.425 47.705 ;
        POLYGON 258.265 47.855 258.265 47.715 258.230 47.715 ;
        RECT 258.265 47.715 259.175 47.855 ;
        RECT 256.770 47.650 257.410 47.705 ;
        POLYGON 257.410 47.705 257.425 47.705 257.410 47.650 ;
        POLYGON 258.230 47.705 258.230 47.655 258.215 47.655 ;
        RECT 258.230 47.685 259.175 47.715 ;
        POLYGON 259.175 47.995 259.240 47.995 259.175 47.685 ;
        POLYGON 260.405 47.985 260.405 47.940 260.400 47.940 ;
        RECT 260.405 47.940 261.930 47.995 ;
        POLYGON 260.400 47.940 260.400 47.785 260.385 47.785 ;
        RECT 260.400 47.830 261.930 47.940 ;
        POLYGON 261.930 48.465 261.950 48.465 261.930 47.830 ;
        POLYGON 264.030 48.435 264.030 48.290 264.025 48.290 ;
        RECT 264.030 48.290 266.725 48.465 ;
        POLYGON 264.025 48.290 264.025 48.020 264.000 48.020 ;
        RECT 264.025 48.245 266.725 48.290 ;
        POLYGON 266.725 48.845 266.740 48.845 266.725 48.245 ;
        POLYGON 270.680 49.450 270.695 49.450 270.695 48.380 ;
        RECT 270.695 49.030 277.795 49.450 ;
        POLYGON 277.795 49.910 277.860 49.030 277.795 49.030 ;
        RECT 270.695 48.520 277.860 49.030 ;
        POLYGON 277.860 49.030 277.885 48.520 277.860 48.520 ;
        RECT 264.025 48.020 266.695 48.245 ;
        POLYGON 264.000 48.020 264.000 47.830 263.985 47.830 ;
        RECT 264.000 47.830 266.695 48.020 ;
        RECT 260.400 47.785 261.910 47.830 ;
        POLYGON 260.385 47.785 260.385 47.690 260.370 47.690 ;
        RECT 260.385 47.690 261.910 47.785 ;
        RECT 258.230 47.655 259.150 47.685 ;
        RECT 256.770 47.635 257.390 47.650 ;
        POLYGON 256.735 47.635 256.735 47.610 256.725 47.610 ;
        RECT 256.735 47.610 257.390 47.635 ;
        POLYGON 255.670 47.610 255.670 47.590 255.665 47.590 ;
        RECT 255.670 47.590 256.070 47.610 ;
        POLYGON 255.665 47.590 255.665 47.570 255.655 47.570 ;
        RECT 255.665 47.570 256.070 47.590 ;
        POLYGON 255.655 47.570 255.655 47.535 255.645 47.535 ;
        RECT 255.655 47.535 256.070 47.570 ;
        RECT 254.350 47.525 255.135 47.535 ;
        RECT 244.575 47.480 245.385 47.525 ;
        RECT 243.500 47.465 244.040 47.480 ;
        POLYGON 244.040 47.480 244.045 47.465 244.040 47.465 ;
        POLYGON 244.575 47.480 244.585 47.480 244.585 47.465 ;
        RECT 244.585 47.465 245.385 47.480 ;
        RECT 243.500 47.420 244.045 47.465 ;
        POLYGON 244.045 47.465 244.070 47.420 244.045 47.420 ;
        POLYGON 244.585 47.465 244.605 47.465 244.605 47.425 ;
        RECT 244.605 47.420 245.385 47.465 ;
        RECT 243.500 47.400 244.070 47.420 ;
        RECT 239.905 47.395 241.070 47.400 ;
        POLYGON 239.905 47.395 239.955 47.395 239.955 47.240 ;
        RECT 239.955 47.340 241.070 47.395 ;
        POLYGON 241.070 47.400 241.090 47.340 241.070 47.340 ;
        POLYGON 242.030 47.400 242.050 47.400 242.050 47.350 ;
        RECT 242.050 47.340 242.850 47.400 ;
        RECT 239.955 47.240 241.090 47.340 ;
        POLYGON 239.955 47.240 239.975 47.240 239.975 47.180 ;
        RECT 239.975 47.170 241.090 47.240 ;
        RECT 236.485 47.030 238.435 47.170 ;
        POLYGON 238.435 47.170 238.480 47.030 238.435 47.030 ;
        POLYGON 239.975 47.170 239.995 47.170 239.995 47.120 ;
        RECT 239.995 47.150 241.090 47.170 ;
        POLYGON 241.090 47.340 241.150 47.150 241.090 47.150 ;
        POLYGON 242.050 47.340 242.105 47.340 242.105 47.215 ;
        RECT 242.105 47.325 242.850 47.340 ;
        POLYGON 242.850 47.400 242.880 47.325 242.850 47.325 ;
        POLYGON 243.500 47.400 243.530 47.400 243.530 47.335 ;
        RECT 243.530 47.365 244.070 47.400 ;
        POLYGON 244.070 47.420 244.095 47.365 244.070 47.365 ;
        POLYGON 244.605 47.420 244.630 47.420 244.630 47.370 ;
        RECT 244.630 47.385 245.385 47.420 ;
        POLYGON 245.385 47.525 245.465 47.385 245.385 47.385 ;
        POLYGON 254.330 47.525 254.330 47.500 254.315 47.500 ;
        RECT 254.330 47.500 255.135 47.525 ;
        POLYGON 254.310 47.500 254.310 47.485 254.305 47.485 ;
        RECT 254.310 47.485 255.135 47.500 ;
        POLYGON 254.305 47.485 254.305 47.405 254.255 47.405 ;
        RECT 254.305 47.470 255.135 47.485 ;
        POLYGON 255.135 47.535 255.160 47.535 255.135 47.470 ;
        POLYGON 255.645 47.535 255.645 47.520 255.640 47.520 ;
        RECT 255.645 47.520 256.070 47.535 ;
        POLYGON 255.640 47.520 255.640 47.470 255.620 47.470 ;
        RECT 255.640 47.470 256.070 47.520 ;
        RECT 254.305 47.405 255.085 47.470 ;
        POLYGON 254.255 47.405 254.255 47.385 254.240 47.385 ;
        RECT 254.255 47.385 255.085 47.405 ;
        RECT 244.630 47.365 245.465 47.385 ;
        RECT 243.530 47.350 244.095 47.365 ;
        POLYGON 244.095 47.365 244.100 47.350 244.095 47.350 ;
        POLYGON 244.630 47.365 244.635 47.365 244.635 47.360 ;
        RECT 244.635 47.350 245.465 47.365 ;
        RECT 243.530 47.335 244.105 47.350 ;
        POLYGON 244.635 47.350 244.640 47.350 244.640 47.345 ;
        RECT 244.640 47.345 245.465 47.350 ;
        POLYGON 243.530 47.335 243.535 47.335 243.535 47.325 ;
        RECT 243.535 47.325 244.105 47.335 ;
        RECT 242.105 47.240 242.880 47.325 ;
        POLYGON 242.880 47.325 242.910 47.240 242.880 47.240 ;
        POLYGON 243.535 47.325 243.555 47.325 243.555 47.285 ;
        RECT 243.555 47.285 244.105 47.325 ;
        POLYGON 243.555 47.285 243.575 47.285 243.575 47.240 ;
        RECT 243.575 47.260 244.105 47.285 ;
        POLYGON 244.105 47.345 244.150 47.260 244.105 47.260 ;
        POLYGON 244.640 47.345 244.680 47.345 244.680 47.260 ;
        RECT 244.680 47.330 245.465 47.345 ;
        POLYGON 245.465 47.385 245.500 47.330 245.465 47.330 ;
        POLYGON 254.240 47.385 254.240 47.350 254.215 47.350 ;
        RECT 254.240 47.365 255.085 47.385 ;
        POLYGON 255.085 47.470 255.135 47.470 255.085 47.365 ;
        POLYGON 255.620 47.470 255.620 47.455 255.615 47.455 ;
        RECT 255.620 47.455 256.070 47.470 ;
        POLYGON 255.615 47.450 255.615 47.380 255.590 47.380 ;
        RECT 255.615 47.380 256.070 47.455 ;
        POLYGON 255.590 47.380 255.590 47.370 255.585 47.370 ;
        RECT 255.590 47.370 256.070 47.380 ;
        RECT 254.240 47.350 254.965 47.365 ;
        POLYGON 254.215 47.350 254.215 47.330 254.200 47.330 ;
        RECT 254.215 47.330 254.965 47.350 ;
        RECT 244.680 47.295 245.500 47.330 ;
        POLYGON 245.500 47.330 245.520 47.295 245.500 47.295 ;
        POLYGON 254.200 47.330 254.200 47.295 254.175 47.295 ;
        RECT 254.200 47.295 254.965 47.330 ;
        RECT 244.680 47.260 245.520 47.295 ;
        RECT 243.575 47.250 244.150 47.260 ;
        POLYGON 244.150 47.260 244.155 47.250 244.150 47.250 ;
        POLYGON 244.680 47.260 244.685 47.260 244.685 47.250 ;
        RECT 244.685 47.250 245.520 47.260 ;
        RECT 243.575 47.240 244.155 47.250 ;
        RECT 242.105 47.215 242.910 47.240 ;
        POLYGON 242.105 47.215 242.130 47.215 242.130 47.150 ;
        RECT 242.130 47.165 242.910 47.215 ;
        POLYGON 242.910 47.240 242.945 47.165 242.910 47.165 ;
        POLYGON 243.575 47.240 243.605 47.240 243.605 47.175 ;
        RECT 243.605 47.165 244.155 47.240 ;
        POLYGON 244.155 47.250 244.200 47.165 244.155 47.165 ;
        POLYGON 244.685 47.250 244.695 47.250 244.695 47.230 ;
        RECT 244.695 47.240 245.520 47.250 ;
        POLYGON 245.520 47.295 245.550 47.240 245.520 47.240 ;
        POLYGON 254.175 47.295 254.175 47.245 254.140 47.245 ;
        RECT 254.175 47.245 254.965 47.295 ;
        RECT 244.695 47.230 245.550 47.240 ;
        POLYGON 244.695 47.230 244.720 47.230 244.720 47.190 ;
        RECT 244.720 47.225 245.550 47.230 ;
        POLYGON 245.550 47.240 245.565 47.225 245.550 47.225 ;
        POLYGON 254.140 47.240 254.140 47.230 254.130 47.230 ;
        RECT 254.140 47.230 254.965 47.245 ;
        RECT 244.720 47.190 245.565 47.225 ;
        POLYGON 244.720 47.190 244.730 47.190 244.730 47.170 ;
        RECT 244.730 47.165 245.565 47.190 ;
        RECT 242.130 47.160 242.945 47.165 ;
        POLYGON 242.945 47.165 242.950 47.160 242.945 47.160 ;
        POLYGON 243.605 47.165 243.610 47.165 243.610 47.160 ;
        RECT 243.610 47.160 244.200 47.165 ;
        RECT 242.130 47.150 242.950 47.160 ;
        RECT 239.995 47.120 241.150 47.150 ;
        POLYGON 239.995 47.120 240.025 47.120 240.025 47.035 ;
        RECT 240.025 47.035 241.150 47.120 ;
        POLYGON 241.150 47.150 241.190 47.035 241.150 47.035 ;
        POLYGON 242.130 47.150 242.175 47.150 242.175 47.040 ;
        RECT 242.175 47.145 242.950 47.150 ;
        POLYGON 242.950 47.160 242.955 47.145 242.950 47.145 ;
        RECT 242.175 47.115 242.955 47.145 ;
        POLYGON 243.610 47.160 243.620 47.160 243.620 47.140 ;
        RECT 243.620 47.145 244.200 47.160 ;
        POLYGON 244.200 47.165 244.215 47.145 244.200 47.145 ;
        POLYGON 244.730 47.165 244.735 47.165 244.735 47.160 ;
        RECT 244.735 47.160 245.565 47.165 ;
        POLYGON 244.735 47.160 244.740 47.160 244.740 47.150 ;
        RECT 244.740 47.145 245.565 47.160 ;
        RECT 243.620 47.140 244.215 47.145 ;
        POLYGON 242.955 47.140 242.970 47.115 242.955 47.115 ;
        POLYGON 243.620 47.140 243.630 47.140 243.630 47.120 ;
        RECT 243.630 47.135 244.215 47.140 ;
        POLYGON 244.215 47.145 244.220 47.135 244.215 47.135 ;
        POLYGON 244.740 47.145 244.745 47.145 244.745 47.140 ;
        RECT 244.745 47.140 245.565 47.145 ;
        POLYGON 245.565 47.225 245.620 47.140 245.565 47.140 ;
        POLYGON 254.130 47.225 254.130 47.200 254.110 47.200 ;
        RECT 254.130 47.200 254.965 47.230 ;
        POLYGON 254.110 47.200 254.110 47.150 254.075 47.150 ;
        RECT 254.110 47.150 254.965 47.200 ;
        POLYGON 254.075 47.150 254.075 47.140 254.070 47.140 ;
        RECT 254.075 47.140 254.965 47.150 ;
        RECT 244.745 47.135 245.620 47.140 ;
        RECT 243.630 47.115 244.220 47.135 ;
        RECT 242.175 47.105 242.970 47.115 ;
        POLYGON 242.970 47.115 242.975 47.105 242.970 47.105 ;
        POLYGON 243.630 47.115 243.635 47.115 243.635 47.110 ;
        RECT 243.635 47.105 244.220 47.115 ;
        RECT 242.175 47.065 242.975 47.105 ;
        POLYGON 242.975 47.105 242.990 47.065 242.975 47.065 ;
        POLYGON 243.635 47.105 243.655 47.105 243.655 47.075 ;
        RECT 243.655 47.065 244.220 47.105 ;
        RECT 242.175 47.050 242.990 47.065 ;
        POLYGON 242.990 47.065 242.995 47.050 242.990 47.050 ;
        POLYGON 243.655 47.065 243.665 47.065 243.665 47.050 ;
        RECT 243.665 47.050 244.220 47.065 ;
        RECT 240.025 47.030 241.190 47.035 ;
        RECT 242.175 47.030 242.995 47.050 ;
        POLYGON 207.630 47.030 207.645 47.030 207.645 46.970 ;
        RECT 207.645 46.970 222.610 47.030 ;
        RECT 182.935 46.415 197.810 46.970 ;
        POLYGON 197.810 46.970 197.880 46.415 197.810 46.415 ;
        POLYGON 207.645 46.970 207.650 46.970 207.650 46.950 ;
        RECT 207.650 46.945 222.610 46.970 ;
        POLYGON 222.610 47.030 222.630 46.945 222.610 46.945 ;
        POLYGON 229.670 47.030 229.690 47.030 229.690 46.955 ;
        RECT 207.650 46.935 222.630 46.945 ;
        RECT 229.690 46.945 233.710 47.030 ;
        POLYGON 233.710 47.030 233.735 46.945 233.710 46.945 ;
        RECT 229.690 46.935 233.735 46.945 ;
        POLYGON 236.485 47.030 236.510 47.030 236.510 46.940 ;
        RECT 236.510 46.985 238.480 47.030 ;
        POLYGON 238.480 47.030 238.495 46.985 238.480 46.985 ;
        POLYGON 240.025 47.030 240.040 47.030 240.040 46.990 ;
        RECT 240.040 46.985 241.190 47.030 ;
        RECT 236.510 46.935 238.495 46.985 ;
        POLYGON 238.495 46.985 238.510 46.935 238.495 46.935 ;
        POLYGON 240.040 46.985 240.060 46.985 240.060 46.935 ;
        RECT 240.060 46.940 241.190 46.985 ;
        POLYGON 241.190 47.030 241.225 46.940 241.190 46.940 ;
        POLYGON 242.175 47.030 242.185 47.030 242.185 47.015 ;
        RECT 240.060 46.935 241.225 46.940 ;
        RECT 242.185 47.005 242.995 47.030 ;
        POLYGON 242.185 47.005 242.220 47.005 242.220 46.935 ;
        RECT 242.220 46.980 242.995 47.005 ;
        POLYGON 242.995 47.050 243.030 46.980 242.995 46.980 ;
        POLYGON 243.665 47.050 243.700 47.050 243.700 46.980 ;
        RECT 243.700 47.030 244.220 47.050 ;
        POLYGON 244.220 47.135 244.280 47.030 244.220 47.030 ;
        POLYGON 244.745 47.135 244.805 47.135 244.805 47.030 ;
        RECT 244.805 47.065 245.620 47.135 ;
        POLYGON 245.620 47.140 245.670 47.065 245.620 47.065 ;
        POLYGON 254.070 47.140 254.070 47.135 254.065 47.135 ;
        RECT 254.070 47.135 254.965 47.140 ;
        POLYGON 254.965 47.365 255.085 47.365 254.965 47.135 ;
        POLYGON 255.585 47.365 255.585 47.315 255.560 47.315 ;
        RECT 255.585 47.360 256.070 47.370 ;
        POLYGON 256.070 47.610 256.175 47.610 256.070 47.360 ;
        POLYGON 256.725 47.610 256.725 47.580 256.715 47.580 ;
        RECT 256.725 47.580 257.390 47.610 ;
        POLYGON 256.715 47.580 256.715 47.560 256.710 47.560 ;
        RECT 256.715 47.570 257.390 47.580 ;
        POLYGON 257.390 47.650 257.410 47.650 257.390 47.570 ;
        POLYGON 258.215 47.650 258.215 47.600 258.200 47.600 ;
        RECT 258.215 47.600 259.150 47.655 ;
        POLYGON 258.200 47.600 258.200 47.570 258.190 47.570 ;
        RECT 258.200 47.575 259.150 47.600 ;
        POLYGON 259.150 47.685 259.175 47.685 259.150 47.575 ;
        POLYGON 260.370 47.685 260.370 47.590 260.355 47.590 ;
        RECT 260.370 47.590 261.910 47.690 ;
        RECT 258.200 47.570 259.105 47.575 ;
        RECT 256.715 47.560 257.305 47.570 ;
        POLYGON 256.710 47.560 256.710 47.420 256.665 47.420 ;
        RECT 256.710 47.420 257.305 47.560 ;
        POLYGON 256.665 47.420 256.665 47.360 256.645 47.360 ;
        RECT 256.665 47.360 257.305 47.420 ;
        RECT 255.585 47.340 256.065 47.360 ;
        POLYGON 256.065 47.360 256.070 47.360 256.065 47.340 ;
        POLYGON 256.645 47.360 256.645 47.345 256.640 47.345 ;
        RECT 256.645 47.345 257.305 47.360 ;
        RECT 255.585 47.315 256.035 47.340 ;
        POLYGON 255.560 47.315 255.560 47.295 255.555 47.295 ;
        RECT 255.560 47.295 256.035 47.315 ;
        POLYGON 255.555 47.295 255.555 47.220 255.520 47.220 ;
        RECT 255.555 47.275 256.035 47.295 ;
        POLYGON 256.035 47.340 256.065 47.340 256.035 47.275 ;
        POLYGON 256.640 47.340 256.640 47.315 256.630 47.315 ;
        RECT 256.640 47.315 257.305 47.345 ;
        POLYGON 256.630 47.315 256.630 47.275 256.610 47.275 ;
        RECT 256.630 47.290 257.305 47.315 ;
        POLYGON 257.305 47.570 257.390 47.570 257.305 47.290 ;
        POLYGON 258.190 47.565 258.190 47.445 258.155 47.445 ;
        RECT 258.190 47.445 259.105 47.570 ;
        POLYGON 258.155 47.445 258.155 47.390 258.140 47.390 ;
        RECT 258.155 47.390 259.105 47.445 ;
        POLYGON 259.105 47.575 259.150 47.575 259.105 47.395 ;
        POLYGON 260.355 47.575 260.355 47.395 260.325 47.395 ;
        RECT 260.355 47.525 261.910 47.590 ;
        POLYGON 261.910 47.830 261.930 47.830 261.910 47.525 ;
        POLYGON 263.985 47.820 263.985 47.755 263.980 47.755 ;
        RECT 263.985 47.755 266.695 47.830 ;
        POLYGON 263.980 47.755 263.980 47.530 263.950 47.530 ;
        RECT 263.980 47.645 266.695 47.755 ;
        POLYGON 266.695 48.245 266.725 48.245 266.695 47.645 ;
        POLYGON 270.695 48.245 270.695 47.730 270.690 47.730 ;
        RECT 270.695 47.915 277.885 48.520 ;
        POLYGON 277.885 48.520 277.910 47.915 277.885 47.915 ;
        RECT 270.695 47.730 277.910 47.915 ;
        RECT 263.980 47.530 266.645 47.645 ;
        RECT 260.355 47.395 261.880 47.525 ;
        POLYGON 258.140 47.390 258.140 47.310 258.115 47.310 ;
        RECT 258.140 47.380 259.105 47.390 ;
        RECT 258.140 47.310 259.020 47.380 ;
        POLYGON 258.115 47.310 258.115 47.295 258.110 47.295 ;
        RECT 258.115 47.295 259.020 47.310 ;
        RECT 256.630 47.275 257.215 47.290 ;
        RECT 255.555 47.220 255.940 47.275 ;
        POLYGON 255.520 47.220 255.520 47.205 255.515 47.205 ;
        RECT 255.520 47.205 255.940 47.220 ;
        POLYGON 255.515 47.205 255.515 47.135 255.480 47.135 ;
        RECT 255.515 47.135 255.940 47.205 ;
        POLYGON 254.065 47.135 254.065 47.065 254.010 47.065 ;
        RECT 254.065 47.065 254.920 47.135 ;
        RECT 244.805 47.030 245.670 47.065 ;
        POLYGON 245.670 47.065 245.695 47.030 245.670 47.030 ;
        POLYGON 254.010 47.065 254.010 47.055 254.000 47.055 ;
        RECT 254.010 47.055 254.920 47.065 ;
        POLYGON 254.000 47.055 254.000 47.030 253.980 47.030 ;
        RECT 254.000 47.045 254.920 47.055 ;
        POLYGON 254.920 47.135 254.965 47.135 254.920 47.045 ;
        POLYGON 255.480 47.135 255.480 47.110 255.470 47.110 ;
        RECT 255.480 47.110 255.940 47.135 ;
        POLYGON 255.470 47.110 255.470 47.045 255.435 47.045 ;
        RECT 255.470 47.075 255.940 47.110 ;
        POLYGON 255.940 47.275 256.035 47.275 255.940 47.075 ;
        POLYGON 256.610 47.270 256.610 47.225 256.590 47.225 ;
        RECT 256.610 47.225 257.215 47.275 ;
        POLYGON 256.590 47.225 256.590 47.205 256.585 47.205 ;
        RECT 256.590 47.205 257.215 47.225 ;
        POLYGON 256.585 47.205 256.585 47.165 256.570 47.165 ;
        RECT 256.585 47.165 257.215 47.205 ;
        POLYGON 256.570 47.165 256.570 47.155 256.565 47.155 ;
        RECT 256.570 47.155 257.215 47.165 ;
        POLYGON 256.565 47.155 256.565 47.075 256.530 47.075 ;
        RECT 256.565 47.075 257.215 47.155 ;
        RECT 255.470 47.045 255.920 47.075 ;
        RECT 254.000 47.030 254.910 47.045 ;
        POLYGON 254.910 47.045 254.920 47.045 254.910 47.030 ;
        POLYGON 255.435 47.040 255.435 47.035 255.430 47.035 ;
        RECT 255.435 47.035 255.920 47.045 ;
        POLYGON 255.920 47.075 255.940 47.075 255.920 47.035 ;
        POLYGON 256.530 47.075 256.530 47.035 256.515 47.035 ;
        RECT 256.530 47.040 257.215 47.075 ;
        POLYGON 257.215 47.290 257.305 47.290 257.215 47.040 ;
        POLYGON 258.110 47.290 258.110 47.225 258.085 47.225 ;
        RECT 258.110 47.225 259.020 47.295 ;
        POLYGON 258.085 47.225 258.085 47.040 258.025 47.040 ;
        RECT 258.085 47.075 259.020 47.225 ;
        POLYGON 259.020 47.380 259.105 47.380 259.020 47.075 ;
        POLYGON 260.325 47.395 260.325 47.240 260.300 47.240 ;
        RECT 260.325 47.240 261.880 47.395 ;
        POLYGON 260.300 47.240 260.300 47.195 260.290 47.195 ;
        RECT 260.300 47.235 261.880 47.240 ;
        POLYGON 261.880 47.525 261.910 47.525 261.880 47.235 ;
        POLYGON 263.950 47.525 263.950 47.490 263.945 47.490 ;
        RECT 263.950 47.490 266.645 47.530 ;
        POLYGON 263.945 47.490 263.945 47.235 263.915 47.235 ;
        RECT 263.945 47.235 266.645 47.490 ;
        RECT 260.300 47.195 261.850 47.235 ;
        POLYGON 260.290 47.195 260.290 47.075 260.265 47.075 ;
        RECT 260.290 47.075 261.850 47.195 ;
        RECT 258.085 47.040 259.005 47.075 ;
        RECT 256.530 47.035 257.210 47.040 ;
        RECT 255.430 47.030 255.920 47.035 ;
        RECT 256.515 47.030 257.210 47.035 ;
        POLYGON 257.210 47.040 257.215 47.040 257.210 47.030 ;
        POLYGON 258.025 47.040 258.025 47.030 258.020 47.030 ;
        RECT 258.025 47.030 259.005 47.040 ;
        POLYGON 259.005 47.075 259.020 47.075 259.005 47.030 ;
        POLYGON 260.265 47.070 260.265 47.030 260.255 47.030 ;
        RECT 260.265 47.030 261.850 47.075 ;
        POLYGON 261.850 47.235 261.880 47.235 261.850 47.035 ;
        POLYGON 263.915 47.215 263.915 47.035 263.885 47.035 ;
        RECT 263.915 47.035 266.645 47.235 ;
        POLYGON 266.645 47.645 266.695 47.645 266.645 47.040 ;
        POLYGON 270.690 47.645 270.690 47.075 270.685 47.075 ;
        RECT 270.690 47.075 277.910 47.730 ;
        RECT 243.700 47.015 244.280 47.030 ;
        POLYGON 244.280 47.030 244.290 47.015 244.280 47.015 ;
        POLYGON 244.805 47.030 244.810 47.030 244.810 47.020 ;
        RECT 244.810 47.015 245.695 47.030 ;
        RECT 243.700 47.005 244.290 47.015 ;
        POLYGON 244.290 47.015 244.295 47.005 244.290 47.005 ;
        POLYGON 244.810 47.015 244.815 47.015 244.815 47.010 ;
        RECT 244.815 47.005 245.695 47.015 ;
        POLYGON 245.695 47.030 245.715 47.005 245.695 47.005 ;
        POLYGON 253.980 47.030 253.980 47.005 253.960 47.005 ;
        RECT 253.980 47.005 254.850 47.030 ;
        RECT 242.220 46.940 243.030 46.980 ;
        RECT 243.700 46.975 244.295 47.005 ;
        POLYGON 243.030 46.975 243.045 46.940 243.030 46.940 ;
        POLYGON 243.700 46.975 243.720 46.975 243.720 46.940 ;
        RECT 243.720 46.965 244.295 46.975 ;
        POLYGON 244.295 47.005 244.320 46.965 244.295 46.965 ;
        POLYGON 244.815 47.005 244.840 47.005 244.840 46.965 ;
        RECT 244.840 46.965 245.715 47.005 ;
        RECT 243.720 46.940 244.320 46.965 ;
        POLYGON 244.320 46.965 244.335 46.940 244.320 46.940 ;
        POLYGON 244.840 46.965 244.855 46.965 244.855 46.940 ;
        RECT 244.855 46.960 245.715 46.965 ;
        POLYGON 245.715 47.005 245.750 46.960 245.715 46.960 ;
        POLYGON 253.960 47.005 253.960 46.975 253.935 46.975 ;
        RECT 253.960 46.975 254.850 47.005 ;
        RECT 242.220 46.935 243.045 46.940 ;
        RECT 243.720 46.935 244.335 46.940 ;
        RECT 244.855 46.935 245.750 46.960 ;
        POLYGON 253.935 46.975 253.935 46.955 253.920 46.955 ;
        RECT 253.935 46.955 254.850 46.975 ;
        POLYGON 207.650 46.935 207.785 46.935 207.785 46.415 ;
        RECT 207.785 46.415 222.630 46.935 ;
        POLYGON 222.630 46.935 222.755 46.415 222.630 46.415 ;
        POLYGON 229.690 46.935 229.745 46.935 229.745 46.705 ;
        RECT 229.745 46.705 233.735 46.935 ;
        POLYGON 229.745 46.705 229.765 46.705 229.765 46.605 ;
        RECT 229.765 46.630 233.735 46.705 ;
        POLYGON 233.735 46.935 233.815 46.630 233.735 46.630 ;
        POLYGON 236.510 46.935 236.555 46.935 236.555 46.775 ;
        RECT 236.555 46.775 238.510 46.935 ;
        RECT 229.765 46.605 233.815 46.630 ;
        POLYGON 236.555 46.775 236.605 46.775 236.605 46.625 ;
        RECT 236.605 46.670 238.510 46.775 ;
        POLYGON 238.510 46.935 238.595 46.670 238.510 46.670 ;
        POLYGON 240.060 46.935 240.095 46.935 240.095 46.840 ;
        RECT 240.095 46.915 241.225 46.935 ;
        POLYGON 241.225 46.935 241.235 46.915 241.225 46.915 ;
        POLYGON 242.220 46.935 242.230 46.935 242.230 46.915 ;
        RECT 242.230 46.920 243.045 46.935 ;
        POLYGON 243.045 46.935 243.055 46.920 243.045 46.920 ;
        POLYGON 243.720 46.935 243.730 46.935 243.730 46.920 ;
        RECT 243.730 46.920 244.335 46.935 ;
        RECT 242.230 46.915 243.055 46.920 ;
        RECT 240.095 46.840 241.235 46.915 ;
        POLYGON 240.095 46.840 240.140 46.840 240.140 46.715 ;
        RECT 240.140 46.820 241.235 46.840 ;
        POLYGON 241.235 46.915 241.270 46.820 241.235 46.820 ;
        POLYGON 242.230 46.915 242.235 46.915 242.235 46.910 ;
        RECT 242.235 46.910 243.055 46.915 ;
        POLYGON 242.235 46.910 242.275 46.910 242.275 46.820 ;
        RECT 242.275 46.830 243.055 46.910 ;
        POLYGON 243.055 46.920 243.100 46.830 243.055 46.830 ;
        POLYGON 243.730 46.920 243.735 46.920 243.735 46.910 ;
        RECT 243.735 46.910 244.335 46.920 ;
        POLYGON 243.735 46.910 243.760 46.910 243.760 46.865 ;
        RECT 243.760 46.870 244.335 46.910 ;
        POLYGON 244.335 46.935 244.380 46.870 244.335 46.870 ;
        POLYGON 244.855 46.935 244.865 46.935 244.865 46.925 ;
        RECT 244.865 46.925 245.750 46.935 ;
        POLYGON 244.865 46.925 244.875 46.925 244.875 46.910 ;
        RECT 244.875 46.915 245.750 46.925 ;
        POLYGON 245.750 46.955 245.780 46.915 245.750 46.915 ;
        POLYGON 253.920 46.955 253.920 46.915 253.890 46.915 ;
        RECT 253.920 46.935 254.850 46.955 ;
        POLYGON 254.850 47.030 254.910 47.030 254.850 46.935 ;
        POLYGON 255.430 47.030 255.430 46.955 255.390 46.955 ;
        RECT 255.430 46.975 255.890 47.030 ;
        POLYGON 255.890 47.030 255.920 47.030 255.890 46.975 ;
        POLYGON 256.515 47.030 256.515 47.010 256.505 47.010 ;
        RECT 256.515 47.015 257.205 47.030 ;
        POLYGON 257.205 47.030 257.210 47.030 257.205 47.015 ;
        POLYGON 258.020 47.025 258.020 47.015 258.015 47.015 ;
        RECT 258.020 47.015 258.975 47.030 ;
        RECT 256.515 47.010 257.200 47.015 ;
        POLYGON 256.505 47.010 256.505 46.975 256.490 46.975 ;
        RECT 256.505 47.005 257.200 47.010 ;
        POLYGON 257.200 47.015 257.205 47.015 257.200 47.005 ;
        RECT 256.505 46.975 257.175 47.005 ;
        RECT 255.430 46.955 255.870 46.975 ;
        POLYGON 255.390 46.955 255.390 46.935 255.375 46.935 ;
        RECT 255.390 46.935 255.870 46.955 ;
        POLYGON 255.870 46.975 255.890 46.975 255.870 46.935 ;
        POLYGON 256.490 46.975 256.490 46.960 256.485 46.960 ;
        RECT 256.490 46.960 257.175 46.975 ;
        POLYGON 256.485 46.960 256.485 46.935 256.475 46.935 ;
        RECT 256.485 46.935 257.175 46.960 ;
        POLYGON 257.175 47.005 257.200 47.005 257.175 46.940 ;
        POLYGON 258.015 47.005 258.015 46.965 258.000 46.965 ;
        RECT 258.015 46.965 258.975 47.015 ;
        POLYGON 258.000 46.965 258.000 46.940 257.990 46.940 ;
        RECT 258.000 46.940 258.975 46.965 ;
        RECT 257.990 46.935 258.975 46.940 ;
        POLYGON 258.975 47.030 259.005 47.030 258.975 46.935 ;
        POLYGON 260.255 47.020 260.255 46.945 260.240 46.945 ;
        RECT 260.255 46.965 261.840 47.030 ;
        POLYGON 261.840 47.030 261.850 47.030 261.840 46.965 ;
        RECT 263.885 47.030 266.645 47.035 ;
        POLYGON 263.885 47.020 263.885 46.965 263.875 46.965 ;
        RECT 263.885 46.965 266.630 47.030 ;
        RECT 260.255 46.945 261.835 46.965 ;
        RECT 260.240 46.935 261.835 46.945 ;
        POLYGON 261.835 46.965 261.840 46.965 261.835 46.940 ;
        RECT 253.920 46.915 254.730 46.935 ;
        RECT 244.875 46.910 245.780 46.915 ;
        POLYGON 244.875 46.910 244.895 46.910 244.895 46.875 ;
        RECT 244.895 46.870 245.780 46.910 ;
        RECT 243.760 46.865 244.380 46.870 ;
        POLYGON 243.760 46.865 243.775 46.865 243.775 46.835 ;
        RECT 243.775 46.860 244.380 46.865 ;
        POLYGON 244.380 46.870 244.385 46.860 244.380 46.860 ;
        POLYGON 244.895 46.870 244.905 46.870 244.905 46.860 ;
        RECT 244.905 46.860 245.780 46.870 ;
        RECT 243.775 46.830 244.385 46.860 ;
        RECT 242.275 46.820 243.100 46.830 ;
        RECT 240.140 46.715 241.270 46.820 ;
        POLYGON 240.140 46.715 240.155 46.715 240.155 46.675 ;
        RECT 240.155 46.690 241.270 46.715 ;
        POLYGON 241.270 46.820 241.325 46.690 241.270 46.690 ;
        POLYGON 242.275 46.820 242.335 46.820 242.335 46.690 ;
        RECT 242.335 46.815 243.100 46.820 ;
        POLYGON 243.100 46.830 243.110 46.815 243.100 46.815 ;
        POLYGON 243.775 46.830 243.785 46.830 243.785 46.820 ;
        RECT 243.785 46.815 244.385 46.830 ;
        RECT 242.335 46.715 243.110 46.815 ;
        POLYGON 243.110 46.815 243.160 46.715 243.110 46.715 ;
        POLYGON 243.785 46.815 243.840 46.815 243.840 46.720 ;
        RECT 243.840 46.765 244.385 46.815 ;
        POLYGON 244.385 46.860 244.445 46.765 244.385 46.765 ;
        POLYGON 244.905 46.860 244.960 46.860 244.960 46.770 ;
        RECT 244.960 46.780 245.780 46.860 ;
        POLYGON 245.780 46.915 245.885 46.780 245.780 46.780 ;
        POLYGON 253.890 46.915 253.890 46.880 253.865 46.880 ;
        RECT 253.890 46.880 254.730 46.915 ;
        POLYGON 253.865 46.880 253.865 46.820 253.805 46.820 ;
        RECT 253.865 46.820 254.730 46.880 ;
        POLYGON 253.805 46.820 253.805 46.780 253.775 46.780 ;
        RECT 253.805 46.780 254.730 46.820 ;
        RECT 244.960 46.765 245.885 46.780 ;
        POLYGON 245.885 46.780 245.895 46.765 245.885 46.765 ;
        POLYGON 253.775 46.780 253.775 46.765 253.760 46.765 ;
        RECT 253.775 46.765 254.730 46.780 ;
        RECT 243.840 46.715 244.445 46.765 ;
        POLYGON 244.445 46.765 244.480 46.715 244.445 46.715 ;
        POLYGON 244.960 46.765 244.995 46.765 244.995 46.715 ;
        RECT 244.995 46.715 245.895 46.765 ;
        RECT 242.335 46.700 243.160 46.715 ;
        POLYGON 243.160 46.715 243.170 46.700 243.160 46.700 ;
        POLYGON 243.840 46.715 243.850 46.715 243.850 46.705 ;
        RECT 243.850 46.700 244.480 46.715 ;
        POLYGON 244.480 46.715 244.490 46.700 244.480 46.700 ;
        POLYGON 244.995 46.715 245.005 46.715 245.005 46.700 ;
        RECT 245.005 46.700 245.895 46.715 ;
        RECT 240.155 46.685 241.325 46.690 ;
        POLYGON 241.325 46.690 241.330 46.685 241.325 46.685 ;
        RECT 242.335 46.685 243.170 46.700 ;
        RECT 240.155 46.670 241.330 46.685 ;
        RECT 236.605 46.640 238.595 46.670 ;
        POLYGON 238.595 46.670 238.605 46.640 238.595 46.640 ;
        POLYGON 240.155 46.670 240.170 46.670 240.170 46.640 ;
        RECT 240.170 46.640 241.330 46.670 ;
        RECT 236.605 46.620 238.605 46.640 ;
        POLYGON 229.765 46.605 229.810 46.605 229.810 46.420 ;
        RECT 182.935 45.765 197.880 46.415 ;
        RECT 207.785 46.405 222.755 46.415 ;
        RECT 229.810 46.415 233.815 46.605 ;
        POLYGON 233.815 46.620 233.880 46.415 233.815 46.415 ;
        POLYGON 236.605 46.620 236.675 46.620 236.675 46.415 ;
        RECT 236.675 46.555 238.605 46.620 ;
        POLYGON 238.605 46.640 238.635 46.555 238.605 46.555 ;
        POLYGON 240.170 46.640 240.205 46.640 240.205 46.560 ;
        RECT 240.205 46.555 241.330 46.640 ;
        RECT 236.675 46.550 238.635 46.555 ;
        POLYGON 238.635 46.555 238.640 46.550 238.635 46.550 ;
        POLYGON 240.205 46.555 240.210 46.555 240.210 46.550 ;
        RECT 240.210 46.550 241.330 46.555 ;
        RECT 229.810 46.405 233.880 46.415 ;
        RECT 236.675 46.410 238.640 46.550 ;
        POLYGON 238.640 46.550 238.690 46.410 238.640 46.410 ;
        POLYGON 240.210 46.550 240.225 46.550 240.225 46.510 ;
        RECT 240.225 46.510 241.330 46.550 ;
        POLYGON 240.225 46.510 240.265 46.510 240.265 46.410 ;
        RECT 240.265 46.470 241.330 46.510 ;
        POLYGON 241.330 46.685 241.425 46.470 241.330 46.470 ;
        POLYGON 242.335 46.685 242.370 46.685 242.370 46.615 ;
        RECT 242.370 46.615 243.170 46.685 ;
        POLYGON 243.170 46.700 243.215 46.615 243.170 46.615 ;
        POLYGON 243.850 46.700 243.900 46.700 243.900 46.620 ;
        RECT 243.900 46.635 244.490 46.700 ;
        POLYGON 244.490 46.700 244.535 46.635 244.490 46.635 ;
        POLYGON 245.005 46.700 245.025 46.700 245.025 46.670 ;
        RECT 245.025 46.690 245.895 46.700 ;
        POLYGON 245.895 46.765 245.955 46.690 245.895 46.690 ;
        POLYGON 253.760 46.765 253.760 46.695 253.695 46.695 ;
        RECT 253.760 46.740 254.730 46.765 ;
        POLYGON 254.730 46.935 254.850 46.935 254.730 46.740 ;
        POLYGON 255.375 46.935 255.375 46.885 255.345 46.885 ;
        RECT 255.375 46.885 255.805 46.935 ;
        POLYGON 255.345 46.885 255.345 46.835 255.320 46.835 ;
        RECT 255.345 46.835 255.805 46.885 ;
        POLYGON 255.320 46.835 255.320 46.780 255.285 46.780 ;
        RECT 255.320 46.810 255.805 46.835 ;
        POLYGON 255.805 46.935 255.870 46.935 255.805 46.810 ;
        POLYGON 256.475 46.935 256.475 46.900 256.460 46.900 ;
        RECT 256.475 46.900 257.100 46.935 ;
        POLYGON 256.460 46.900 256.460 46.810 256.415 46.810 ;
        RECT 256.460 46.810 257.100 46.900 ;
        RECT 255.320 46.780 255.765 46.810 ;
        POLYGON 255.285 46.780 255.285 46.740 255.260 46.740 ;
        RECT 255.285 46.750 255.765 46.780 ;
        POLYGON 255.765 46.810 255.805 46.810 255.765 46.750 ;
        POLYGON 256.415 46.810 256.415 46.750 256.385 46.750 ;
        RECT 256.415 46.750 257.100 46.810 ;
        RECT 255.285 46.740 255.695 46.750 ;
        RECT 253.760 46.700 254.705 46.740 ;
        POLYGON 254.705 46.740 254.730 46.740 254.705 46.700 ;
        POLYGON 255.260 46.740 255.260 46.705 255.240 46.705 ;
        RECT 255.260 46.705 255.695 46.740 ;
        RECT 253.760 46.695 254.525 46.700 ;
        RECT 245.025 46.670 245.955 46.690 ;
        POLYGON 245.025 46.670 245.040 46.670 245.040 46.645 ;
        RECT 245.040 46.645 245.955 46.670 ;
        POLYGON 245.040 46.645 245.045 46.645 245.045 46.635 ;
        RECT 245.045 46.635 245.955 46.645 ;
        RECT 243.900 46.615 244.535 46.635 ;
        POLYGON 242.370 46.615 242.385 46.615 242.385 46.590 ;
        RECT 242.385 46.590 243.215 46.615 ;
        POLYGON 242.385 46.590 242.450 46.590 242.450 46.470 ;
        RECT 242.450 46.585 243.215 46.590 ;
        POLYGON 243.215 46.615 243.230 46.585 243.215 46.585 ;
        POLYGON 243.900 46.615 243.920 46.615 243.920 46.585 ;
        RECT 243.920 46.585 244.535 46.615 ;
        RECT 242.450 46.490 243.230 46.585 ;
        POLYGON 243.230 46.585 243.285 46.490 243.230 46.490 ;
        POLYGON 243.920 46.585 243.975 46.585 243.975 46.500 ;
        RECT 243.975 46.575 244.535 46.585 ;
        POLYGON 244.535 46.635 244.575 46.575 244.535 46.575 ;
        POLYGON 245.045 46.635 245.085 46.635 245.085 46.580 ;
        RECT 245.085 46.625 245.955 46.635 ;
        POLYGON 245.955 46.690 246.015 46.625 245.955 46.625 ;
        POLYGON 253.695 46.690 253.695 46.665 253.670 46.665 ;
        RECT 253.695 46.665 254.525 46.695 ;
        POLYGON 253.670 46.665 253.670 46.625 253.635 46.625 ;
        RECT 253.670 46.625 254.525 46.665 ;
        RECT 245.085 46.610 246.015 46.625 ;
        POLYGON 246.015 46.625 246.025 46.610 246.015 46.610 ;
        POLYGON 253.635 46.625 253.635 46.610 253.620 46.610 ;
        RECT 253.635 46.610 254.525 46.625 ;
        RECT 245.085 46.575 246.025 46.610 ;
        RECT 243.975 46.555 244.575 46.575 ;
        POLYGON 244.575 46.575 244.595 46.555 244.575 46.555 ;
        POLYGON 245.085 46.575 245.100 46.575 245.100 46.555 ;
        RECT 245.100 46.555 246.025 46.575 ;
        RECT 243.975 46.535 244.595 46.555 ;
        POLYGON 244.595 46.555 244.605 46.535 244.595 46.535 ;
        POLYGON 245.100 46.555 245.115 46.555 245.115 46.535 ;
        RECT 245.115 46.535 246.025 46.555 ;
        RECT 243.975 46.500 244.605 46.535 ;
        POLYGON 243.975 46.500 243.980 46.500 243.980 46.490 ;
        RECT 243.980 46.490 244.605 46.500 ;
        RECT 236.675 46.405 238.690 46.410 ;
        RECT 240.265 46.405 241.425 46.470 ;
        RECT 242.450 46.465 243.285 46.490 ;
        RECT 171.490 45.580 175.575 45.765 ;
        POLYGON 171.435 45.580 171.435 45.395 171.400 45.395 ;
        RECT 171.435 45.395 175.575 45.580 ;
        RECT 166.390 45.275 168.405 45.395 ;
        RECT 163.315 45.250 164.520 45.270 ;
        POLYGON 163.270 45.250 163.270 45.235 163.260 45.235 ;
        RECT 163.270 45.235 164.520 45.250 ;
        RECT 161.240 45.175 162.170 45.235 ;
        POLYGON 161.190 45.175 161.190 45.120 161.150 45.120 ;
        RECT 161.190 45.170 162.170 45.175 ;
        POLYGON 162.170 45.235 162.210 45.235 162.170 45.170 ;
        POLYGON 163.260 45.230 163.260 45.170 163.225 45.170 ;
        RECT 163.260 45.170 164.520 45.235 ;
        RECT 161.190 45.120 162.065 45.170 ;
        RECT 158.190 45.110 158.640 45.120 ;
        RECT 153.325 45.105 156.290 45.110 ;
        POLYGON 156.290 45.110 156.295 45.110 156.290 45.105 ;
        POLYGON 158.115 45.110 158.115 45.105 158.110 45.105 ;
        RECT 158.115 45.105 158.640 45.110 ;
        RECT 153.325 45.095 156.130 45.105 ;
        POLYGON 153.325 45.095 153.360 45.095 153.360 45.085 ;
        RECT 153.360 45.085 156.130 45.095 ;
        RECT 151.010 45.070 151.640 45.085 ;
        POLYGON 151.640 45.085 151.660 45.070 151.640 45.070 ;
        POLYGON 153.365 45.085 153.410 45.085 153.410 45.070 ;
        RECT 153.410 45.070 156.130 45.085 ;
        RECT 151.010 45.065 151.660 45.070 ;
        POLYGON 150.380 45.065 150.400 45.020 150.380 45.020 ;
        POLYGON 151.010 45.065 151.060 45.065 151.060 45.020 ;
        RECT 151.060 45.020 151.660 45.065 ;
        RECT 117.265 45.010 150.400 45.020 ;
        POLYGON 150.400 45.020 150.405 45.010 150.400 45.010 ;
        POLYGON 151.060 45.020 151.075 45.020 151.075 45.010 ;
        RECT 151.075 45.010 151.660 45.020 ;
        RECT 117.265 44.940 150.405 45.010 ;
        POLYGON 150.405 45.010 150.435 44.940 150.405 44.940 ;
        POLYGON 151.075 45.010 151.170 45.010 151.170 44.940 ;
        RECT 151.170 44.985 151.660 45.010 ;
        POLYGON 151.660 45.070 151.805 44.985 151.660 44.985 ;
        POLYGON 153.410 45.070 153.530 45.070 153.530 45.035 ;
        RECT 153.530 45.060 156.130 45.070 ;
        POLYGON 156.130 45.105 156.290 45.105 156.130 45.060 ;
        POLYGON 158.110 45.105 158.110 45.065 158.050 45.065 ;
        RECT 158.110 45.065 158.640 45.105 ;
        POLYGON 158.050 45.065 158.050 45.060 158.045 45.060 ;
        RECT 158.050 45.060 158.640 45.065 ;
        RECT 153.530 45.055 156.120 45.060 ;
        POLYGON 156.120 45.060 156.130 45.060 156.120 45.055 ;
        POLYGON 158.045 45.060 158.045 45.055 158.035 45.055 ;
        RECT 158.045 45.055 158.640 45.060 ;
        RECT 153.530 45.045 156.085 45.055 ;
        POLYGON 156.085 45.055 156.120 45.055 156.085 45.045 ;
        POLYGON 158.035 45.055 158.035 45.045 158.025 45.045 ;
        RECT 158.035 45.045 158.640 45.055 ;
        RECT 153.530 45.035 155.970 45.045 ;
        POLYGON 153.530 45.035 153.575 45.035 153.575 45.025 ;
        RECT 153.575 45.025 155.970 45.035 ;
        POLYGON 153.580 45.025 153.585 45.025 153.585 45.020 ;
        RECT 153.585 45.020 155.970 45.025 ;
        POLYGON 153.585 45.020 153.740 45.020 153.740 44.985 ;
        RECT 153.740 45.015 155.970 45.020 ;
        POLYGON 155.970 45.045 156.085 45.045 155.970 45.015 ;
        POLYGON 158.025 45.045 158.025 45.015 157.985 45.015 ;
        RECT 158.025 45.020 158.640 45.045 ;
        POLYGON 158.640 45.120 158.765 45.120 158.640 45.020 ;
        POLYGON 159.505 45.120 159.505 45.110 159.495 45.110 ;
        RECT 159.505 45.110 160.185 45.120 ;
        POLYGON 159.495 45.110 159.495 45.085 159.465 45.085 ;
        RECT 159.495 45.085 160.185 45.110 ;
        POLYGON 159.465 45.085 159.465 45.020 159.395 45.020 ;
        RECT 159.465 45.020 160.185 45.085 ;
        RECT 158.025 45.015 158.580 45.020 ;
        RECT 153.740 45.010 155.935 45.015 ;
        POLYGON 155.935 45.015 155.970 45.015 155.935 45.010 ;
        POLYGON 157.985 45.015 157.985 45.010 157.980 45.010 ;
        RECT 157.985 45.010 158.580 45.015 ;
        RECT 153.740 44.985 155.805 45.010 ;
        RECT 151.170 44.975 151.810 44.985 ;
        POLYGON 151.810 44.985 151.820 44.975 151.810 44.975 ;
        POLYGON 153.740 44.985 153.760 44.985 153.760 44.980 ;
        RECT 153.760 44.980 155.805 44.985 ;
        POLYGON 155.805 45.010 155.935 45.010 155.805 44.980 ;
        POLYGON 157.980 45.010 157.980 44.995 157.960 44.995 ;
        RECT 157.980 44.995 158.580 45.010 ;
        POLYGON 157.960 44.995 157.960 44.990 157.945 44.990 ;
        RECT 157.960 44.990 158.580 44.995 ;
        POLYGON 157.945 44.990 157.945 44.980 157.930 44.980 ;
        RECT 157.945 44.980 158.580 44.990 ;
        POLYGON 153.760 44.980 153.790 44.980 153.790 44.975 ;
        RECT 153.790 44.975 155.755 44.980 ;
        RECT 151.170 44.950 151.820 44.975 ;
        POLYGON 151.820 44.975 151.875 44.950 151.820 44.950 ;
        POLYGON 153.795 44.975 153.915 44.975 153.915 44.950 ;
        RECT 153.915 44.965 155.755 44.975 ;
        POLYGON 155.755 44.980 155.805 44.980 155.755 44.965 ;
        POLYGON 157.930 44.980 157.930 44.965 157.910 44.965 ;
        RECT 157.930 44.970 158.580 44.980 ;
        POLYGON 158.580 45.020 158.640 45.020 158.580 44.970 ;
        POLYGON 159.395 45.020 159.395 44.985 159.355 44.985 ;
        RECT 159.395 44.985 160.185 45.020 ;
        POLYGON 159.355 44.985 159.355 44.970 159.340 44.970 ;
        RECT 159.355 44.970 160.185 44.985 ;
        RECT 157.930 44.965 158.505 44.970 ;
        RECT 153.915 44.950 155.660 44.965 ;
        POLYGON 155.660 44.965 155.755 44.965 155.660 44.950 ;
        POLYGON 157.910 44.965 157.910 44.950 157.885 44.950 ;
        RECT 157.910 44.950 158.505 44.965 ;
        RECT 151.170 44.940 151.875 44.950 ;
        RECT 117.265 44.930 150.435 44.940 ;
        POLYGON 150.435 44.940 150.440 44.930 150.435 44.930 ;
        RECT 117.265 44.920 150.440 44.930 ;
        POLYGON 151.170 44.940 151.190 44.940 151.190 44.925 ;
        RECT 151.190 44.925 151.875 44.940 ;
        POLYGON 150.440 44.925 150.445 44.920 150.440 44.920 ;
        RECT 117.265 44.885 150.445 44.920 ;
        POLYGON 151.190 44.925 151.210 44.925 151.210 44.910 ;
        RECT 151.210 44.910 151.875 44.925 ;
        POLYGON 150.445 44.910 150.460 44.885 150.445 44.885 ;
        POLYGON 151.210 44.910 151.245 44.910 151.245 44.885 ;
        RECT 151.245 44.905 151.875 44.910 ;
        POLYGON 151.875 44.950 151.955 44.905 151.875 44.905 ;
        POLYGON 153.915 44.950 153.940 44.950 153.940 44.945 ;
        RECT 153.940 44.945 155.635 44.950 ;
        POLYGON 155.635 44.950 155.660 44.950 155.635 44.945 ;
        POLYGON 157.885 44.950 157.885 44.945 157.875 44.945 ;
        RECT 157.885 44.945 158.505 44.950 ;
        POLYGON 153.940 44.945 154.000 44.945 154.000 44.935 ;
        RECT 154.000 44.935 155.570 44.945 ;
        POLYGON 155.570 44.945 155.630 44.945 155.570 44.935 ;
        POLYGON 157.875 44.945 157.875 44.935 157.860 44.935 ;
        RECT 157.875 44.935 158.505 44.945 ;
        POLYGON 154.005 44.935 154.115 44.935 154.115 44.915 ;
        RECT 154.115 44.920 155.460 44.935 ;
        POLYGON 155.460 44.935 155.570 44.935 155.460 44.920 ;
        POLYGON 157.860 44.935 157.860 44.920 157.835 44.920 ;
        RECT 157.860 44.920 158.505 44.935 ;
        POLYGON 158.505 44.970 158.580 44.970 158.505 44.920 ;
        POLYGON 159.340 44.970 159.340 44.920 159.290 44.920 ;
        RECT 159.340 44.945 160.185 44.970 ;
        POLYGON 160.185 45.120 160.345 45.120 160.185 44.945 ;
        POLYGON 161.150 45.120 161.150 44.990 161.060 44.990 ;
        RECT 161.150 45.020 162.065 45.120 ;
        POLYGON 162.065 45.170 162.170 45.170 162.065 45.020 ;
        POLYGON 163.225 45.165 163.225 45.020 163.145 45.020 ;
        RECT 163.225 45.020 164.520 45.170 ;
        RECT 161.150 44.990 161.905 45.020 ;
        POLYGON 161.060 44.990 161.060 44.965 161.040 44.965 ;
        RECT 161.060 44.965 161.905 44.990 ;
        POLYGON 161.040 44.965 161.040 44.945 161.025 44.945 ;
        RECT 161.040 44.945 161.905 44.965 ;
        RECT 159.340 44.920 160.145 44.945 ;
        RECT 154.115 44.915 155.455 44.920 ;
        POLYGON 155.455 44.920 155.460 44.920 155.455 44.915 ;
        POLYGON 157.835 44.920 157.835 44.915 157.830 44.915 ;
        RECT 157.835 44.915 158.385 44.920 ;
        POLYGON 154.140 44.915 154.220 44.915 154.220 44.905 ;
        RECT 154.220 44.910 155.390 44.915 ;
        POLYGON 155.390 44.915 155.450 44.915 155.390 44.910 ;
        POLYGON 157.830 44.915 157.830 44.910 157.820 44.910 ;
        RECT 157.830 44.910 158.385 44.915 ;
        RECT 154.220 44.905 155.280 44.910 ;
        RECT 151.245 44.890 151.955 44.905 ;
        POLYGON 151.955 44.905 151.985 44.890 151.955 44.890 ;
        POLYGON 154.220 44.905 154.295 44.905 154.295 44.895 ;
        RECT 154.295 44.895 155.280 44.905 ;
        POLYGON 155.280 44.910 155.390 44.910 155.280 44.895 ;
        POLYGON 157.820 44.910 157.820 44.895 157.795 44.895 ;
        RECT 157.820 44.895 158.385 44.910 ;
        POLYGON 154.295 44.895 154.360 44.895 154.360 44.890 ;
        RECT 154.360 44.890 155.205 44.895 ;
        POLYGON 155.205 44.895 155.245 44.895 155.205 44.890 ;
        POLYGON 157.795 44.895 157.795 44.890 157.790 44.890 ;
        RECT 157.795 44.890 158.385 44.895 ;
        RECT 151.245 44.885 151.985 44.890 ;
        RECT 117.265 44.810 150.460 44.885 ;
        POLYGON 150.460 44.885 150.490 44.810 150.460 44.810 ;
        POLYGON 151.245 44.885 151.275 44.885 151.275 44.860 ;
        RECT 151.275 44.860 151.985 44.885 ;
        RECT 117.265 44.795 150.490 44.810 ;
        POLYGON 151.275 44.860 151.345 44.860 151.345 44.805 ;
        RECT 151.345 44.840 151.985 44.860 ;
        POLYGON 151.985 44.890 152.070 44.840 151.985 44.840 ;
        POLYGON 154.360 44.890 154.430 44.890 154.430 44.885 ;
        RECT 154.430 44.885 155.050 44.890 ;
        POLYGON 154.430 44.885 154.475 44.885 154.475 44.880 ;
        RECT 154.475 44.880 155.050 44.885 ;
        POLYGON 155.050 44.890 155.205 44.890 155.050 44.880 ;
        POLYGON 157.790 44.890 157.790 44.885 157.780 44.885 ;
        RECT 157.790 44.885 158.385 44.890 ;
        POLYGON 157.780 44.885 157.780 44.880 157.775 44.880 ;
        RECT 157.780 44.880 158.385 44.885 ;
        POLYGON 154.530 44.880 154.635 44.880 154.635 44.875 ;
        RECT 154.635 44.875 155.035 44.880 ;
        POLYGON 155.035 44.880 155.045 44.880 155.035 44.875 ;
        POLYGON 157.775 44.880 157.775 44.875 157.765 44.875 ;
        RECT 157.775 44.875 158.385 44.880 ;
        POLYGON 154.655 44.875 154.840 44.875 154.840 44.870 ;
        POLYGON 154.840 44.875 154.910 44.875 154.840 44.870 ;
        POLYGON 157.765 44.875 157.765 44.870 157.760 44.870 ;
        RECT 157.765 44.870 158.385 44.875 ;
        POLYGON 157.760 44.870 157.760 44.845 157.720 44.845 ;
        RECT 157.760 44.845 158.385 44.870 ;
        POLYGON 157.715 44.845 157.715 44.840 157.705 44.840 ;
        RECT 157.715 44.840 158.385 44.845 ;
        RECT 151.345 44.825 152.070 44.840 ;
        POLYGON 152.070 44.840 152.105 44.825 152.070 44.825 ;
        POLYGON 157.705 44.840 157.705 44.825 157.680 44.825 ;
        RECT 157.705 44.835 158.385 44.840 ;
        POLYGON 158.385 44.920 158.505 44.920 158.385 44.835 ;
        POLYGON 159.290 44.920 159.290 44.895 159.260 44.895 ;
        RECT 159.290 44.905 160.145 44.920 ;
        POLYGON 160.145 44.945 160.185 44.945 160.145 44.905 ;
        POLYGON 161.025 44.945 161.025 44.905 160.995 44.905 ;
        RECT 161.025 44.905 161.905 44.945 ;
        RECT 159.290 44.895 159.940 44.905 ;
        POLYGON 159.260 44.895 159.260 44.835 159.190 44.835 ;
        RECT 159.260 44.835 159.940 44.895 ;
        RECT 157.705 44.825 158.235 44.835 ;
        RECT 151.345 44.805 152.105 44.825 ;
        POLYGON 150.490 44.805 150.495 44.795 150.490 44.795 ;
        RECT 117.265 44.785 150.495 44.795 ;
        POLYGON 151.345 44.805 151.365 44.805 151.365 44.790 ;
        RECT 151.365 44.795 152.105 44.805 ;
        POLYGON 152.105 44.825 152.160 44.795 152.105 44.795 ;
        POLYGON 157.680 44.825 157.680 44.815 157.665 44.815 ;
        RECT 157.680 44.815 158.235 44.825 ;
        POLYGON 157.665 44.815 157.665 44.795 157.630 44.795 ;
        RECT 157.665 44.795 158.235 44.815 ;
        RECT 151.365 44.790 152.165 44.795 ;
        POLYGON 150.495 44.790 150.500 44.785 150.495 44.785 ;
        RECT 117.265 44.780 150.500 44.785 ;
        POLYGON 151.365 44.790 151.380 44.790 151.380 44.780 ;
        RECT 151.380 44.780 152.165 44.790 ;
        RECT 117.265 44.775 150.505 44.780 ;
        POLYGON 150.505 44.780 150.515 44.775 150.505 44.775 ;
        POLYGON 151.380 44.780 151.385 44.780 151.385 44.775 ;
        RECT 151.385 44.775 152.165 44.780 ;
        RECT 117.265 44.755 150.515 44.775 ;
        POLYGON 150.515 44.775 150.540 44.755 150.515 44.755 ;
        POLYGON 151.385 44.775 151.415 44.775 151.415 44.755 ;
        RECT 151.415 44.755 152.165 44.775 ;
        RECT 117.265 44.740 150.540 44.755 ;
        POLYGON 150.540 44.755 150.555 44.740 150.540 44.740 ;
        POLYGON 151.415 44.755 151.435 44.755 151.435 44.740 ;
        RECT 151.435 44.750 152.165 44.755 ;
        POLYGON 152.165 44.795 152.260 44.750 152.165 44.750 ;
        POLYGON 157.630 44.795 157.630 44.750 157.555 44.750 ;
        RECT 157.630 44.750 158.235 44.795 ;
        RECT 151.435 44.740 152.260 44.750 ;
        RECT 117.265 44.730 150.555 44.740 ;
        POLYGON 117.265 44.730 117.270 44.730 117.270 44.670 ;
        RECT 117.270 44.705 150.555 44.730 ;
        POLYGON 150.555 44.740 150.600 44.705 150.555 44.705 ;
        POLYGON 151.435 44.740 151.465 44.740 151.465 44.720 ;
        RECT 151.465 44.720 152.260 44.740 ;
        POLYGON 151.465 44.720 151.485 44.720 151.485 44.710 ;
        RECT 151.485 44.715 152.260 44.720 ;
        POLYGON 152.260 44.750 152.330 44.715 152.260 44.715 ;
        POLYGON 157.555 44.750 157.555 44.745 157.545 44.745 ;
        RECT 157.555 44.745 158.235 44.750 ;
        POLYGON 157.545 44.745 157.545 44.715 157.495 44.715 ;
        RECT 157.545 44.730 158.235 44.745 ;
        POLYGON 158.235 44.835 158.385 44.835 158.235 44.730 ;
        POLYGON 159.190 44.835 159.190 44.780 159.130 44.780 ;
        RECT 159.190 44.780 159.940 44.835 ;
        POLYGON 159.125 44.780 159.125 44.745 159.085 44.745 ;
        RECT 159.125 44.745 159.940 44.780 ;
        POLYGON 159.085 44.745 159.085 44.730 159.065 44.730 ;
        RECT 159.085 44.730 159.940 44.745 ;
        RECT 157.545 44.715 158.190 44.730 ;
        RECT 151.485 44.710 152.330 44.715 ;
        POLYGON 152.330 44.715 152.345 44.710 152.330 44.710 ;
        POLYGON 157.495 44.715 157.495 44.710 157.485 44.710 ;
        RECT 157.495 44.710 158.190 44.715 ;
        POLYGON 151.485 44.710 151.490 44.710 151.490 44.705 ;
        RECT 151.490 44.705 152.350 44.710 ;
        RECT 117.270 44.695 150.600 44.705 ;
        POLYGON 150.600 44.705 150.615 44.695 150.600 44.695 ;
        POLYGON 151.490 44.705 151.505 44.705 151.505 44.695 ;
        RECT 151.505 44.695 152.350 44.705 ;
        RECT 117.270 44.635 150.615 44.695 ;
        POLYGON 150.615 44.695 150.695 44.635 150.615 44.635 ;
        POLYGON 151.505 44.695 151.585 44.695 151.585 44.645 ;
        RECT 151.585 44.680 152.350 44.695 ;
        POLYGON 152.350 44.710 152.415 44.680 152.350 44.680 ;
        POLYGON 157.485 44.710 157.485 44.680 157.420 44.680 ;
        RECT 157.485 44.695 158.190 44.710 ;
        POLYGON 158.190 44.730 158.235 44.730 158.190 44.695 ;
        POLYGON 159.065 44.730 159.065 44.695 159.020 44.695 ;
        RECT 159.065 44.695 159.940 44.730 ;
        POLYGON 159.940 44.905 160.145 44.905 159.940 44.695 ;
        POLYGON 160.995 44.905 160.995 44.880 160.975 44.880 ;
        RECT 160.995 44.880 161.905 44.905 ;
        POLYGON 160.975 44.880 160.975 44.790 160.905 44.790 ;
        RECT 160.975 44.790 161.905 44.880 ;
        POLYGON 161.905 45.020 162.065 45.020 161.905 44.790 ;
        POLYGON 163.145 45.020 163.145 44.985 163.125 44.985 ;
        RECT 163.145 44.985 164.520 45.020 ;
        POLYGON 163.125 44.985 163.125 44.970 163.120 44.970 ;
        RECT 163.125 44.970 164.520 44.985 ;
        POLYGON 163.120 44.970 163.120 44.935 163.095 44.935 ;
        RECT 163.120 44.935 164.520 44.970 ;
        POLYGON 163.095 44.935 163.095 44.790 163.005 44.790 ;
        RECT 163.095 44.865 164.520 44.935 ;
        POLYGON 164.520 45.270 164.705 45.270 164.520 44.865 ;
        POLYGON 166.325 45.270 166.325 45.215 166.300 45.215 ;
        RECT 166.325 45.215 168.405 45.275 ;
        POLYGON 166.300 45.215 166.300 45.090 166.250 45.090 ;
        RECT 166.300 45.090 168.405 45.215 ;
        POLYGON 166.250 45.090 166.250 44.965 166.190 44.965 ;
        RECT 166.250 44.965 168.405 45.090 ;
        POLYGON 166.190 44.965 166.190 44.900 166.165 44.900 ;
        RECT 166.190 44.905 168.405 44.965 ;
        POLYGON 168.405 45.395 168.555 45.395 168.405 44.905 ;
        POLYGON 171.400 45.395 171.400 45.205 171.365 45.205 ;
        RECT 171.400 45.205 175.575 45.395 ;
        POLYGON 171.365 45.205 171.365 45.135 171.350 45.135 ;
        RECT 171.365 45.135 175.575 45.205 ;
        POLYGON 171.350 45.135 171.350 44.905 171.295 44.905 ;
        RECT 171.350 44.905 175.575 45.135 ;
        RECT 166.190 44.900 168.255 44.905 ;
        POLYGON 166.165 44.900 166.165 44.870 166.150 44.870 ;
        RECT 166.165 44.870 168.255 44.900 ;
        RECT 163.095 44.810 164.495 44.865 ;
        POLYGON 164.495 44.865 164.520 44.865 164.495 44.810 ;
        POLYGON 166.150 44.865 166.150 44.810 166.120 44.810 ;
        RECT 166.150 44.810 168.255 44.870 ;
        RECT 163.095 44.790 164.435 44.810 ;
        POLYGON 160.905 44.790 160.905 44.700 160.830 44.700 ;
        RECT 160.905 44.765 161.890 44.790 ;
        POLYGON 161.890 44.790 161.905 44.790 161.890 44.765 ;
        POLYGON 163.005 44.785 163.005 44.770 162.995 44.770 ;
        RECT 163.005 44.770 164.435 44.790 ;
        POLYGON 162.995 44.770 162.995 44.765 162.990 44.765 ;
        RECT 162.995 44.765 164.435 44.770 ;
        RECT 160.905 44.700 161.675 44.765 ;
        RECT 157.485 44.680 158.130 44.695 ;
        RECT 151.585 44.645 152.415 44.680 ;
        POLYGON 152.415 44.680 152.500 44.645 152.415 44.645 ;
        POLYGON 157.420 44.680 157.420 44.665 157.385 44.665 ;
        RECT 157.420 44.665 158.130 44.680 ;
        POLYGON 157.385 44.665 157.385 44.655 157.370 44.655 ;
        RECT 157.385 44.660 158.130 44.665 ;
        POLYGON 158.130 44.695 158.190 44.695 158.130 44.660 ;
        POLYGON 159.020 44.695 159.020 44.690 159.015 44.690 ;
        RECT 159.020 44.690 159.775 44.695 ;
        POLYGON 159.015 44.690 159.015 44.660 158.975 44.660 ;
        RECT 159.015 44.660 159.775 44.690 ;
        RECT 157.385 44.655 157.960 44.660 ;
        POLYGON 157.365 44.655 157.365 44.645 157.345 44.645 ;
        RECT 157.365 44.645 157.960 44.655 ;
        POLYGON 151.585 44.645 151.600 44.645 151.600 44.635 ;
        RECT 151.600 44.635 152.505 44.645 ;
        RECT 117.270 44.630 150.695 44.635 ;
        POLYGON 150.695 44.635 150.700 44.630 150.695 44.630 ;
        POLYGON 151.600 44.635 151.605 44.635 151.605 44.630 ;
        RECT 151.605 44.630 152.505 44.635 ;
        POLYGON 152.505 44.645 152.535 44.630 152.505 44.630 ;
        POLYGON 157.345 44.645 157.345 44.630 157.315 44.630 ;
        RECT 157.345 44.630 157.960 44.645 ;
        RECT 117.270 44.570 150.700 44.630 ;
        POLYGON 117.270 44.570 117.285 44.570 117.285 43.870 ;
        RECT 117.285 44.555 150.700 44.570 ;
        POLYGON 150.700 44.630 150.805 44.555 150.700 44.555 ;
        POLYGON 151.605 44.630 151.680 44.630 151.680 44.580 ;
        RECT 151.680 44.615 152.535 44.630 ;
        POLYGON 152.535 44.630 152.575 44.615 152.535 44.615 ;
        POLYGON 157.315 44.630 157.315 44.615 157.280 44.615 ;
        RECT 157.315 44.615 157.960 44.630 ;
        RECT 151.680 44.605 152.575 44.615 ;
        POLYGON 152.575 44.615 152.600 44.605 152.575 44.605 ;
        POLYGON 157.280 44.615 157.280 44.605 157.260 44.605 ;
        RECT 157.280 44.605 157.960 44.615 ;
        RECT 151.680 44.580 152.600 44.605 ;
        POLYGON 151.680 44.580 151.720 44.580 151.720 44.555 ;
        RECT 151.720 44.565 152.600 44.580 ;
        POLYGON 152.600 44.605 152.715 44.565 152.600 44.565 ;
        POLYGON 157.260 44.605 157.260 44.595 157.240 44.595 ;
        RECT 157.260 44.595 157.960 44.605 ;
        POLYGON 157.240 44.595 157.240 44.575 157.195 44.575 ;
        RECT 157.240 44.575 157.960 44.595 ;
        POLYGON 157.195 44.575 157.195 44.565 157.175 44.565 ;
        RECT 157.195 44.565 157.960 44.575 ;
        RECT 151.720 44.560 152.715 44.565 ;
        POLYGON 152.715 44.565 152.730 44.560 152.715 44.560 ;
        POLYGON 157.175 44.565 157.175 44.560 157.160 44.560 ;
        RECT 157.175 44.560 157.960 44.565 ;
        RECT 151.720 44.555 152.730 44.560 ;
        POLYGON 152.730 44.560 152.735 44.555 152.730 44.555 ;
        POLYGON 157.160 44.560 157.160 44.555 157.150 44.555 ;
        RECT 157.160 44.555 157.960 44.560 ;
        POLYGON 157.960 44.660 158.130 44.660 157.960 44.555 ;
        POLYGON 158.975 44.660 158.975 44.640 158.950 44.640 ;
        RECT 158.975 44.640 159.775 44.660 ;
        POLYGON 158.950 44.640 158.950 44.585 158.885 44.585 ;
        RECT 158.950 44.585 159.775 44.640 ;
        POLYGON 158.885 44.585 158.885 44.555 158.845 44.555 ;
        RECT 158.885 44.555 159.775 44.585 ;
        RECT 117.285 44.475 150.805 44.555 ;
        POLYGON 150.805 44.555 150.920 44.475 150.805 44.475 ;
        POLYGON 151.720 44.555 151.730 44.555 151.730 44.550 ;
        RECT 151.730 44.550 152.740 44.555 ;
        POLYGON 151.730 44.550 151.850 44.550 151.850 44.475 ;
        RECT 151.850 44.505 152.740 44.550 ;
        POLYGON 152.740 44.555 152.880 44.505 152.740 44.505 ;
        POLYGON 157.150 44.555 157.150 44.540 157.110 44.540 ;
        RECT 157.150 44.540 157.865 44.555 ;
        POLYGON 157.110 44.540 157.110 44.505 157.030 44.505 ;
        RECT 157.110 44.505 157.865 44.540 ;
        RECT 151.850 44.495 152.880 44.505 ;
        POLYGON 152.880 44.505 152.905 44.495 152.880 44.495 ;
        POLYGON 157.030 44.505 157.030 44.495 157.010 44.495 ;
        RECT 157.030 44.495 157.865 44.505 ;
        POLYGON 157.865 44.555 157.960 44.555 157.865 44.495 ;
        POLYGON 158.845 44.555 158.845 44.495 158.765 44.495 ;
        RECT 158.845 44.540 159.775 44.555 ;
        POLYGON 159.775 44.695 159.940 44.695 159.775 44.540 ;
        POLYGON 160.830 44.695 160.830 44.555 160.710 44.555 ;
        RECT 160.830 44.555 161.675 44.700 ;
        POLYGON 160.710 44.555 160.710 44.540 160.695 44.540 ;
        RECT 160.710 44.540 161.675 44.555 ;
        RECT 158.845 44.510 159.740 44.540 ;
        POLYGON 159.740 44.540 159.775 44.540 159.740 44.510 ;
        POLYGON 160.695 44.540 160.695 44.510 160.670 44.510 ;
        RECT 160.695 44.510 161.675 44.540 ;
        RECT 158.845 44.495 159.720 44.510 ;
        RECT 151.850 44.490 152.905 44.495 ;
        POLYGON 152.905 44.495 152.925 44.490 152.905 44.490 ;
        POLYGON 157.010 44.495 157.010 44.490 156.995 44.490 ;
        RECT 157.010 44.490 157.780 44.495 ;
        RECT 151.850 44.475 152.930 44.490 ;
        RECT 117.285 44.420 150.920 44.475 ;
        POLYGON 150.920 44.475 151.010 44.420 150.920 44.420 ;
        POLYGON 151.850 44.475 151.875 44.475 151.875 44.460 ;
        RECT 151.875 44.460 152.930 44.475 ;
        POLYGON 151.875 44.460 151.940 44.460 151.940 44.420 ;
        RECT 151.940 44.445 152.930 44.460 ;
        POLYGON 152.930 44.490 153.070 44.445 152.930 44.445 ;
        POLYGON 156.995 44.490 156.995 44.485 156.975 44.485 ;
        RECT 156.995 44.485 157.780 44.490 ;
        POLYGON 156.975 44.485 156.975 44.470 156.940 44.470 ;
        RECT 156.975 44.470 157.780 44.485 ;
        POLYGON 156.940 44.470 156.940 44.445 156.860 44.445 ;
        RECT 156.940 44.445 157.780 44.470 ;
        POLYGON 157.780 44.495 157.865 44.495 157.780 44.445 ;
        POLYGON 158.765 44.495 158.765 44.445 158.695 44.445 ;
        RECT 158.765 44.490 159.720 44.495 ;
        POLYGON 159.720 44.510 159.740 44.510 159.720 44.490 ;
        POLYGON 160.670 44.510 160.670 44.490 160.655 44.490 ;
        RECT 160.670 44.490 161.675 44.510 ;
        POLYGON 161.675 44.765 161.890 44.765 161.675 44.490 ;
        POLYGON 162.990 44.760 162.990 44.545 162.860 44.545 ;
        RECT 162.990 44.700 164.435 44.765 ;
        POLYGON 164.435 44.810 164.495 44.810 164.435 44.700 ;
        POLYGON 166.120 44.805 166.120 44.755 166.095 44.755 ;
        RECT 166.120 44.755 168.255 44.810 ;
        POLYGON 166.095 44.755 166.095 44.700 166.070 44.700 ;
        RECT 166.095 44.700 168.255 44.755 ;
        RECT 162.990 44.545 164.260 44.700 ;
        POLYGON 162.860 44.545 162.860 44.495 162.825 44.495 ;
        RECT 162.860 44.495 164.260 44.545 ;
        RECT 158.765 44.445 159.495 44.490 ;
        RECT 151.940 44.430 153.070 44.445 ;
        POLYGON 153.070 44.445 153.125 44.430 153.070 44.430 ;
        POLYGON 156.860 44.445 156.860 44.440 156.845 44.440 ;
        RECT 156.860 44.440 157.690 44.445 ;
        POLYGON 156.840 44.440 156.840 44.430 156.810 44.430 ;
        RECT 156.840 44.430 157.690 44.440 ;
        RECT 151.940 44.425 153.125 44.430 ;
        POLYGON 153.125 44.430 153.145 44.425 153.125 44.425 ;
        POLYGON 156.810 44.430 156.810 44.425 156.795 44.425 ;
        RECT 156.810 44.425 157.690 44.430 ;
        RECT 151.940 44.420 153.145 44.425 ;
        RECT 117.285 44.410 151.010 44.420 ;
        POLYGON 151.010 44.420 151.020 44.410 151.010 44.410 ;
        POLYGON 151.940 44.420 151.955 44.420 151.955 44.410 ;
        RECT 151.955 44.415 153.145 44.420 ;
        POLYGON 153.145 44.425 153.170 44.415 153.145 44.415 ;
        POLYGON 156.795 44.425 156.795 44.415 156.770 44.415 ;
        RECT 156.795 44.415 157.690 44.425 ;
        RECT 151.955 44.410 153.170 44.415 ;
        RECT 117.285 44.380 151.020 44.410 ;
        POLYGON 151.020 44.410 151.075 44.380 151.020 44.380 ;
        POLYGON 151.955 44.410 151.975 44.410 151.975 44.400 ;
        RECT 151.975 44.400 153.170 44.410 ;
        POLYGON 153.170 44.415 153.240 44.400 153.170 44.400 ;
        POLYGON 156.770 44.415 156.770 44.400 156.725 44.400 ;
        RECT 156.770 44.400 157.690 44.415 ;
        POLYGON 151.975 44.400 152.010 44.400 152.010 44.380 ;
        RECT 152.010 44.380 153.240 44.400 ;
        RECT 117.285 44.320 151.075 44.380 ;
        POLYGON 151.075 44.380 151.170 44.320 151.075 44.320 ;
        POLYGON 152.010 44.380 152.115 44.380 152.115 44.320 ;
        RECT 152.115 44.375 153.240 44.380 ;
        POLYGON 153.240 44.400 153.325 44.375 153.240 44.375 ;
        POLYGON 156.725 44.400 156.725 44.395 156.715 44.395 ;
        RECT 156.725 44.395 157.690 44.400 ;
        POLYGON 157.690 44.445 157.780 44.445 157.690 44.395 ;
        POLYGON 158.695 44.445 158.695 44.405 158.640 44.405 ;
        RECT 158.695 44.405 159.495 44.445 ;
        POLYGON 158.640 44.405 158.640 44.400 158.635 44.400 ;
        RECT 158.640 44.400 159.495 44.405 ;
        POLYGON 158.635 44.400 158.635 44.395 158.625 44.395 ;
        RECT 158.635 44.395 159.495 44.400 ;
        POLYGON 156.715 44.395 156.715 44.380 156.665 44.380 ;
        RECT 156.715 44.380 157.590 44.395 ;
        POLYGON 156.665 44.380 156.665 44.375 156.645 44.375 ;
        RECT 156.665 44.375 157.590 44.380 ;
        RECT 152.115 44.365 153.325 44.375 ;
        POLYGON 153.325 44.375 153.360 44.365 153.325 44.365 ;
        POLYGON 156.645 44.375 156.645 44.365 156.610 44.365 ;
        RECT 156.645 44.365 157.590 44.375 ;
        RECT 152.115 44.355 153.365 44.365 ;
        POLYGON 153.365 44.365 153.410 44.355 153.365 44.355 ;
        POLYGON 156.610 44.365 156.610 44.355 156.570 44.355 ;
        RECT 156.610 44.355 157.590 44.365 ;
        RECT 152.115 44.340 153.410 44.355 ;
        POLYGON 153.410 44.355 153.460 44.340 153.410 44.340 ;
        POLYGON 156.570 44.355 156.570 44.340 156.510 44.340 ;
        RECT 156.570 44.340 157.590 44.355 ;
        POLYGON 157.590 44.395 157.690 44.395 157.590 44.340 ;
        POLYGON 158.625 44.395 158.625 44.365 158.580 44.365 ;
        RECT 158.625 44.365 159.495 44.395 ;
        POLYGON 158.580 44.365 158.580 44.340 158.545 44.340 ;
        RECT 158.580 44.340 159.495 44.365 ;
        RECT 152.115 44.325 153.460 44.340 ;
        POLYGON 153.460 44.340 153.530 44.325 153.460 44.325 ;
        POLYGON 156.510 44.340 156.510 44.330 156.485 44.330 ;
        RECT 156.510 44.330 157.425 44.340 ;
        POLYGON 156.480 44.330 156.480 44.325 156.460 44.325 ;
        RECT 156.480 44.325 157.425 44.330 ;
        RECT 152.115 44.320 153.530 44.325 ;
        POLYGON 153.530 44.325 153.575 44.320 153.530 44.320 ;
        POLYGON 156.460 44.325 156.460 44.320 156.440 44.320 ;
        RECT 156.460 44.320 157.425 44.325 ;
        RECT 117.285 44.270 151.170 44.320 ;
        POLYGON 151.170 44.320 151.245 44.270 151.170 44.270 ;
        POLYGON 152.115 44.320 152.210 44.320 152.210 44.270 ;
        RECT 152.210 44.315 153.580 44.320 ;
        POLYGON 156.440 44.320 156.440 44.315 156.415 44.315 ;
        RECT 156.440 44.315 157.425 44.320 ;
        RECT 152.210 44.285 153.585 44.315 ;
        POLYGON 153.585 44.315 153.735 44.285 153.585 44.285 ;
        POLYGON 156.415 44.315 156.415 44.290 156.300 44.290 ;
        RECT 156.415 44.290 157.425 44.315 ;
        POLYGON 156.295 44.290 156.295 44.285 156.290 44.285 ;
        RECT 156.295 44.285 157.425 44.290 ;
        RECT 152.210 44.280 153.740 44.285 ;
        POLYGON 153.740 44.285 153.760 44.280 153.740 44.280 ;
        POLYGON 156.285 44.285 156.285 44.280 156.260 44.280 ;
        RECT 156.285 44.280 157.425 44.285 ;
        RECT 152.210 44.275 153.765 44.280 ;
        POLYGON 153.765 44.280 153.790 44.275 153.765 44.275 ;
        POLYGON 156.260 44.280 156.260 44.275 156.235 44.275 ;
        RECT 156.260 44.275 157.425 44.280 ;
        RECT 152.210 44.270 153.795 44.275 ;
        RECT 117.285 44.145 151.245 44.270 ;
        POLYGON 151.245 44.270 151.465 44.145 151.245 44.145 ;
        POLYGON 152.210 44.270 152.220 44.270 152.220 44.265 ;
        RECT 152.220 44.265 153.795 44.270 ;
        POLYGON 152.220 44.265 152.290 44.265 152.290 44.225 ;
        RECT 152.290 44.255 153.795 44.265 ;
        POLYGON 153.795 44.275 153.935 44.255 153.795 44.255 ;
        POLYGON 156.235 44.275 156.235 44.270 156.210 44.270 ;
        RECT 156.235 44.270 157.425 44.275 ;
        POLYGON 156.210 44.270 156.210 44.255 156.130 44.255 ;
        RECT 156.210 44.255 157.425 44.270 ;
        RECT 152.290 44.240 153.940 44.255 ;
        POLYGON 153.940 44.255 154.005 44.240 153.940 44.240 ;
        POLYGON 156.120 44.255 156.120 44.250 156.085 44.250 ;
        RECT 156.120 44.250 157.425 44.255 ;
        POLYGON 157.425 44.340 157.590 44.340 157.425 44.250 ;
        POLYGON 158.545 44.340 158.545 44.315 158.505 44.315 ;
        RECT 158.545 44.315 159.495 44.340 ;
        POLYGON 158.505 44.315 158.505 44.250 158.410 44.250 ;
        RECT 158.505 44.295 159.495 44.315 ;
        POLYGON 159.495 44.490 159.720 44.490 159.495 44.295 ;
        POLYGON 160.655 44.490 160.655 44.445 160.615 44.445 ;
        RECT 160.655 44.445 161.620 44.490 ;
        POLYGON 160.615 44.445 160.615 44.360 160.540 44.360 ;
        RECT 160.615 44.420 161.620 44.445 ;
        POLYGON 161.620 44.490 161.675 44.490 161.620 44.420 ;
        POLYGON 162.825 44.490 162.825 44.445 162.790 44.445 ;
        RECT 162.825 44.445 164.260 44.495 ;
        POLYGON 162.790 44.445 162.790 44.425 162.775 44.425 ;
        RECT 162.790 44.425 164.260 44.445 ;
        RECT 160.615 44.360 161.555 44.420 ;
        POLYGON 160.540 44.360 160.540 44.350 160.535 44.350 ;
        RECT 160.540 44.350 161.555 44.360 ;
        POLYGON 160.535 44.350 160.535 44.295 160.485 44.295 ;
        RECT 160.535 44.345 161.555 44.350 ;
        POLYGON 161.555 44.420 161.620 44.420 161.555 44.345 ;
        POLYGON 162.775 44.420 162.775 44.350 162.725 44.350 ;
        RECT 162.775 44.365 164.260 44.425 ;
        POLYGON 164.260 44.700 164.435 44.700 164.260 44.365 ;
        POLYGON 166.070 44.700 166.070 44.575 166.015 44.575 ;
        RECT 166.070 44.575 168.255 44.700 ;
        POLYGON 166.015 44.575 166.015 44.425 165.945 44.425 ;
        RECT 166.015 44.465 168.255 44.575 ;
        POLYGON 168.255 44.905 168.405 44.905 168.255 44.465 ;
        POLYGON 171.295 44.905 171.295 44.755 171.260 44.755 ;
        RECT 171.295 44.755 175.575 44.905 ;
        POLYGON 171.260 44.755 171.260 44.485 171.195 44.485 ;
        RECT 171.260 44.485 175.575 44.755 ;
        POLYGON 171.195 44.485 171.195 44.465 171.190 44.465 ;
        RECT 171.195 44.465 175.575 44.485 ;
        RECT 166.015 44.425 168.240 44.465 ;
        POLYGON 165.945 44.425 165.945 44.365 165.915 44.365 ;
        RECT 165.945 44.420 168.240 44.425 ;
        POLYGON 168.240 44.465 168.255 44.465 168.240 44.420 ;
        POLYGON 171.190 44.465 171.190 44.420 171.180 44.420 ;
        RECT 171.190 44.420 175.575 44.465 ;
        RECT 165.945 44.365 168.050 44.420 ;
        RECT 162.775 44.350 164.065 44.365 ;
        RECT 160.535 44.295 161.305 44.345 ;
        RECT 158.505 44.250 159.375 44.295 ;
        POLYGON 156.080 44.250 156.080 44.240 156.025 44.240 ;
        RECT 156.080 44.240 157.365 44.250 ;
        RECT 152.290 44.225 154.005 44.240 ;
        POLYGON 154.005 44.240 154.110 44.225 154.005 44.225 ;
        POLYGON 156.025 44.240 156.025 44.230 155.970 44.230 ;
        RECT 156.025 44.230 157.365 44.240 ;
        POLYGON 155.970 44.230 155.970 44.225 155.935 44.225 ;
        RECT 155.970 44.225 157.365 44.230 ;
        POLYGON 152.290 44.225 152.450 44.225 152.450 44.145 ;
        RECT 152.450 44.215 154.140 44.225 ;
        POLYGON 154.140 44.225 154.220 44.215 154.140 44.215 ;
        POLYGON 155.935 44.225 155.935 44.220 155.870 44.220 ;
        RECT 155.935 44.220 157.365 44.225 ;
        POLYGON 155.870 44.220 155.870 44.215 155.840 44.215 ;
        RECT 155.870 44.215 157.365 44.220 ;
        POLYGON 157.365 44.250 157.425 44.250 157.365 44.215 ;
        POLYGON 158.410 44.250 158.410 44.245 158.400 44.245 ;
        RECT 158.410 44.245 159.375 44.250 ;
        POLYGON 158.400 44.245 158.400 44.235 158.385 44.235 ;
        RECT 158.400 44.235 159.375 44.245 ;
        POLYGON 158.385 44.235 158.385 44.215 158.350 44.215 ;
        RECT 158.385 44.215 159.375 44.235 ;
        RECT 152.450 44.205 154.220 44.215 ;
        POLYGON 154.220 44.215 154.295 44.205 154.220 44.205 ;
        POLYGON 155.840 44.215 155.840 44.210 155.805 44.210 ;
        RECT 155.840 44.210 157.315 44.215 ;
        POLYGON 155.800 44.210 155.800 44.205 155.755 44.205 ;
        RECT 155.800 44.205 157.315 44.210 ;
        RECT 152.450 44.195 154.295 44.205 ;
        POLYGON 154.295 44.205 154.390 44.195 154.295 44.195 ;
        POLYGON 155.755 44.205 155.755 44.195 155.660 44.195 ;
        RECT 155.755 44.195 157.315 44.205 ;
        RECT 152.450 44.190 154.430 44.195 ;
        POLYGON 154.430 44.195 154.470 44.190 154.430 44.190 ;
        POLYGON 155.650 44.195 155.650 44.190 155.635 44.190 ;
        RECT 155.650 44.190 157.315 44.195 ;
        POLYGON 157.315 44.215 157.365 44.215 157.315 44.190 ;
        POLYGON 158.350 44.215 158.350 44.190 158.310 44.190 ;
        RECT 158.350 44.200 159.375 44.215 ;
        POLYGON 159.375 44.295 159.495 44.295 159.375 44.200 ;
        POLYGON 160.485 44.295 160.485 44.205 160.395 44.205 ;
        RECT 160.485 44.205 161.305 44.295 ;
        RECT 158.350 44.190 159.290 44.200 ;
        RECT 152.450 44.185 154.475 44.190 ;
        POLYGON 154.475 44.190 154.530 44.185 154.475 44.185 ;
        POLYGON 155.570 44.190 155.570 44.185 155.515 44.185 ;
        RECT 155.570 44.185 157.160 44.190 ;
        RECT 152.450 44.180 154.530 44.185 ;
        POLYGON 154.530 44.185 154.640 44.180 154.530 44.180 ;
        POLYGON 155.515 44.185 155.515 44.180 155.460 44.180 ;
        RECT 155.515 44.180 157.160 44.185 ;
        RECT 152.450 44.175 154.655 44.180 ;
        POLYGON 154.655 44.180 154.715 44.175 154.655 44.175 ;
        POLYGON 155.445 44.180 155.445 44.175 155.390 44.175 ;
        RECT 155.445 44.175 157.160 44.180 ;
        RECT 152.450 44.170 154.715 44.175 ;
        POLYGON 154.715 44.175 154.905 44.170 154.715 44.170 ;
        POLYGON 155.280 44.175 155.280 44.170 155.250 44.170 ;
        RECT 155.280 44.170 157.160 44.175 ;
        RECT 152.450 44.145 157.160 44.170 ;
        RECT 117.285 44.085 151.465 44.145 ;
        POLYGON 151.465 44.145 151.585 44.085 151.465 44.085 ;
        POLYGON 152.450 44.145 152.470 44.145 152.470 44.135 ;
        RECT 152.470 44.135 157.160 44.145 ;
        POLYGON 152.470 44.135 152.505 44.135 152.505 44.120 ;
        RECT 152.505 44.120 157.160 44.135 ;
        POLYGON 152.505 44.120 152.575 44.120 152.575 44.085 ;
        RECT 152.575 44.115 157.160 44.120 ;
        POLYGON 157.160 44.190 157.315 44.190 157.160 44.115 ;
        POLYGON 158.310 44.190 158.310 44.145 158.235 44.145 ;
        RECT 158.310 44.145 159.290 44.190 ;
        POLYGON 158.235 44.145 158.235 44.115 158.190 44.115 ;
        RECT 158.235 44.135 159.290 44.145 ;
        POLYGON 159.290 44.200 159.375 44.200 159.290 44.135 ;
        POLYGON 160.395 44.200 160.395 44.135 160.330 44.135 ;
        RECT 160.395 44.135 161.305 44.205 ;
        RECT 158.235 44.115 159.260 44.135 ;
        RECT 152.575 44.110 157.150 44.115 ;
        POLYGON 157.150 44.115 157.160 44.115 157.150 44.110 ;
        POLYGON 158.190 44.115 158.190 44.110 158.180 44.110 ;
        RECT 158.190 44.110 159.260 44.115 ;
        POLYGON 159.260 44.135 159.290 44.135 159.260 44.110 ;
        POLYGON 160.330 44.135 160.330 44.110 160.305 44.110 ;
        RECT 160.330 44.110 161.305 44.135 ;
        RECT 152.575 44.085 157.030 44.110 ;
        RECT 117.285 44.015 151.585 44.085 ;
        POLYGON 151.585 44.085 151.710 44.015 151.585 44.015 ;
        POLYGON 152.575 44.085 152.690 44.085 152.690 44.030 ;
        RECT 152.690 44.055 157.030 44.085 ;
        POLYGON 157.030 44.110 157.150 44.110 157.030 44.055 ;
        POLYGON 158.180 44.110 158.180 44.100 158.165 44.100 ;
        RECT 158.180 44.100 159.015 44.110 ;
        POLYGON 158.165 44.100 158.165 44.080 158.130 44.080 ;
        RECT 158.165 44.080 159.015 44.100 ;
        POLYGON 158.130 44.080 158.130 44.055 158.085 44.055 ;
        RECT 158.130 44.055 159.015 44.080 ;
        RECT 152.690 44.030 156.940 44.055 ;
        POLYGON 152.690 44.030 152.715 44.030 152.715 44.020 ;
        RECT 152.715 44.020 156.940 44.030 ;
        POLYGON 152.720 44.020 152.730 44.020 152.730 44.015 ;
        RECT 152.730 44.015 156.940 44.020 ;
        POLYGON 156.940 44.055 157.030 44.055 156.940 44.015 ;
        POLYGON 158.085 44.055 158.085 44.015 158.015 44.015 ;
        RECT 158.085 44.015 159.015 44.055 ;
        RECT 117.285 44.010 151.710 44.015 ;
        POLYGON 151.710 44.015 151.730 44.010 151.710 44.010 ;
        POLYGON 152.730 44.015 152.740 44.015 152.740 44.010 ;
        RECT 152.740 44.010 156.890 44.015 ;
        RECT 117.285 43.940 151.730 44.010 ;
        POLYGON 151.730 44.010 151.875 43.940 151.730 43.940 ;
        POLYGON 152.740 44.010 152.905 44.010 152.905 43.940 ;
        RECT 152.905 43.995 156.890 44.010 ;
        POLYGON 156.890 44.015 156.940 44.015 156.890 43.995 ;
        POLYGON 158.015 44.015 158.015 43.995 157.980 43.995 ;
        RECT 158.015 43.995 159.015 44.015 ;
        RECT 152.905 43.940 156.745 43.995 ;
        RECT 117.285 43.920 151.875 43.940 ;
        POLYGON 151.875 43.940 151.915 43.920 151.875 43.920 ;
        POLYGON 152.905 43.940 152.930 43.940 152.930 43.930 ;
        RECT 152.930 43.935 156.745 43.940 ;
        POLYGON 156.745 43.995 156.890 43.995 156.745 43.935 ;
        POLYGON 157.980 43.995 157.980 43.965 157.920 43.965 ;
        RECT 157.980 43.965 159.015 43.995 ;
        POLYGON 157.920 43.965 157.920 43.935 157.865 43.935 ;
        RECT 157.920 43.935 159.015 43.965 ;
        POLYGON 159.015 44.110 159.260 44.110 159.015 43.935 ;
        POLYGON 160.305 44.110 160.305 44.065 160.260 44.065 ;
        RECT 160.305 44.065 161.305 44.110 ;
        POLYGON 160.260 44.065 160.260 43.995 160.185 43.995 ;
        RECT 160.260 44.060 161.305 44.065 ;
        POLYGON 161.305 44.345 161.555 44.345 161.305 44.060 ;
        POLYGON 162.725 44.345 162.725 44.205 162.630 44.205 ;
        RECT 162.725 44.205 164.065 44.350 ;
        POLYGON 162.630 44.205 162.630 44.065 162.525 44.065 ;
        RECT 162.630 44.065 164.065 44.205 ;
        POLYGON 162.525 44.065 162.525 44.060 162.520 44.060 ;
        RECT 162.525 44.060 164.065 44.065 ;
        RECT 160.260 44.015 161.265 44.060 ;
        POLYGON 161.265 44.060 161.305 44.060 161.265 44.015 ;
        POLYGON 162.520 44.060 162.520 44.015 162.490 44.015 ;
        RECT 162.520 44.030 164.065 44.060 ;
        POLYGON 164.065 44.365 164.260 44.365 164.065 44.030 ;
        POLYGON 165.915 44.365 165.915 44.240 165.850 44.240 ;
        RECT 165.915 44.240 168.050 44.365 ;
        POLYGON 165.850 44.240 165.850 44.220 165.845 44.220 ;
        RECT 165.850 44.220 168.050 44.240 ;
        POLYGON 165.845 44.220 165.845 44.115 165.790 44.115 ;
        RECT 165.845 44.115 168.050 44.220 ;
        POLYGON 165.790 44.115 165.790 44.030 165.750 44.030 ;
        RECT 165.790 44.030 168.050 44.115 ;
        RECT 162.520 44.015 164.010 44.030 ;
        RECT 160.260 43.995 161.210 44.015 ;
        POLYGON 160.185 43.995 160.185 43.970 160.165 43.970 ;
        RECT 160.185 43.970 161.210 43.995 ;
        POLYGON 160.165 43.970 160.165 43.955 160.145 43.955 ;
        RECT 160.165 43.960 161.210 43.970 ;
        POLYGON 161.210 44.015 161.265 44.015 161.210 43.960 ;
        POLYGON 162.490 44.015 162.490 43.960 162.450 43.960 ;
        RECT 162.490 43.960 164.010 44.015 ;
        RECT 160.165 43.955 160.975 43.960 ;
        POLYGON 160.145 43.955 160.145 43.935 160.125 43.935 ;
        RECT 160.145 43.935 160.975 43.955 ;
        RECT 152.930 43.930 156.725 43.935 ;
        POLYGON 152.930 43.930 152.955 43.930 152.955 43.920 ;
        RECT 152.955 43.925 156.725 43.930 ;
        POLYGON 156.725 43.935 156.745 43.935 156.725 43.925 ;
        POLYGON 157.865 43.935 157.865 43.925 157.845 43.925 ;
        RECT 157.865 43.925 158.970 43.935 ;
        RECT 152.955 43.920 156.625 43.925 ;
        RECT 117.285 43.910 151.915 43.920 ;
        POLYGON 151.915 43.920 151.940 43.910 151.915 43.910 ;
        POLYGON 152.955 43.920 152.970 43.920 152.970 43.915 ;
        RECT 152.970 43.915 156.625 43.920 ;
        POLYGON 152.970 43.915 152.980 43.915 152.980 43.910 ;
        RECT 152.980 43.910 156.625 43.915 ;
        RECT 117.285 43.895 151.940 43.910 ;
        POLYGON 151.940 43.910 151.975 43.895 151.940 43.895 ;
        POLYGON 152.980 43.910 153.020 43.910 153.020 43.895 ;
        RECT 153.020 43.895 156.625 43.910 ;
        RECT 117.285 43.885 151.975 43.895 ;
        POLYGON 151.975 43.895 151.990 43.885 151.975 43.885 ;
        POLYGON 153.020 43.895 153.045 43.895 153.045 43.885 ;
        RECT 153.045 43.890 156.625 43.895 ;
        POLYGON 156.625 43.925 156.725 43.925 156.625 43.890 ;
        POLYGON 157.845 43.925 157.845 43.895 157.780 43.895 ;
        RECT 157.845 43.900 158.970 43.925 ;
        POLYGON 158.970 43.935 159.015 43.935 158.970 43.900 ;
        POLYGON 160.125 43.935 160.125 43.900 160.085 43.900 ;
        RECT 160.125 43.900 160.975 43.935 ;
        RECT 157.845 43.895 158.825 43.900 ;
        POLYGON 157.780 43.895 157.780 43.890 157.770 43.890 ;
        RECT 157.780 43.890 158.825 43.895 ;
        RECT 153.045 43.885 156.510 43.890 ;
        RECT 117.285 43.785 151.990 43.885 ;
        POLYGON 151.990 43.885 152.220 43.785 151.990 43.785 ;
        POLYGON 153.045 43.885 153.085 43.885 153.085 43.870 ;
        RECT 153.085 43.870 156.510 43.885 ;
        POLYGON 153.090 43.870 153.145 43.870 153.145 43.845 ;
        RECT 153.145 43.845 156.510 43.870 ;
        POLYGON 156.510 43.890 156.625 43.890 156.510 43.845 ;
        POLYGON 157.770 43.890 157.770 43.850 157.690 43.850 ;
        RECT 157.770 43.850 158.825 43.890 ;
        POLYGON 157.690 43.850 157.690 43.845 157.675 43.845 ;
        RECT 157.690 43.845 158.825 43.850 ;
        POLYGON 153.145 43.845 153.225 43.845 153.225 43.820 ;
        RECT 153.225 43.820 156.360 43.845 ;
        POLYGON 153.225 43.820 153.330 43.820 153.330 43.785 ;
        RECT 153.330 43.795 156.360 43.820 ;
        POLYGON 156.360 43.845 156.510 43.845 156.360 43.795 ;
        POLYGON 157.675 43.845 157.675 43.805 157.590 43.805 ;
        RECT 157.675 43.810 158.825 43.845 ;
        POLYGON 158.825 43.900 158.965 43.900 158.825 43.810 ;
        POLYGON 160.085 43.900 160.085 43.810 159.990 43.810 ;
        RECT 160.085 43.810 160.975 43.900 ;
        RECT 157.675 43.805 158.765 43.810 ;
        POLYGON 157.590 43.805 157.590 43.795 157.570 43.795 ;
        RECT 157.590 43.795 158.765 43.805 ;
        RECT 153.330 43.785 156.295 43.795 ;
        RECT 117.285 43.765 152.220 43.785 ;
        POLYGON 152.220 43.785 152.265 43.765 152.220 43.765 ;
        POLYGON 153.330 43.785 153.365 43.785 153.365 43.775 ;
        RECT 153.365 43.775 156.295 43.785 ;
        POLYGON 153.365 43.775 153.395 43.775 153.395 43.765 ;
        RECT 153.395 43.770 156.295 43.775 ;
        POLYGON 156.295 43.795 156.360 43.795 156.295 43.770 ;
        POLYGON 157.570 43.795 157.570 43.770 157.515 43.770 ;
        RECT 157.570 43.770 158.765 43.795 ;
        RECT 153.395 43.765 156.155 43.770 ;
        RECT 117.285 43.755 152.265 43.765 ;
        POLYGON 152.265 43.765 152.290 43.755 152.265 43.755 ;
        POLYGON 153.395 43.765 153.430 43.765 153.430 43.755 ;
        RECT 153.430 43.755 156.155 43.765 ;
        RECT 117.285 43.750 152.290 43.755 ;
        POLYGON 152.290 43.755 152.310 43.750 152.290 43.750 ;
        POLYGON 153.430 43.755 153.445 43.755 153.445 43.750 ;
        RECT 153.445 43.750 156.155 43.755 ;
        RECT 117.285 43.690 152.310 43.750 ;
        POLYGON 152.310 43.750 152.470 43.690 152.310 43.690 ;
        POLYGON 153.445 43.750 153.480 43.750 153.480 43.740 ;
        RECT 153.480 43.740 156.155 43.750 ;
        POLYGON 153.480 43.740 153.495 43.740 153.495 43.735 ;
        RECT 153.495 43.735 156.155 43.740 ;
        POLYGON 153.495 43.735 153.580 43.735 153.580 43.710 ;
        RECT 153.580 43.730 156.155 43.735 ;
        POLYGON 156.155 43.770 156.295 43.770 156.155 43.730 ;
        POLYGON 157.515 43.770 157.515 43.730 157.425 43.730 ;
        RECT 157.515 43.765 158.765 43.770 ;
        POLYGON 158.765 43.810 158.825 43.810 158.765 43.765 ;
        POLYGON 159.990 43.810 159.990 43.795 159.975 43.795 ;
        RECT 159.990 43.795 160.975 43.810 ;
        POLYGON 159.975 43.795 159.975 43.765 159.940 43.765 ;
        RECT 159.975 43.765 160.975 43.795 ;
        RECT 157.515 43.730 158.550 43.765 ;
        RECT 153.580 43.710 156.095 43.730 ;
        POLYGON 156.095 43.730 156.155 43.730 156.095 43.710 ;
        POLYGON 157.425 43.730 157.425 43.710 157.375 43.710 ;
        RECT 157.425 43.710 158.550 43.730 ;
        POLYGON 153.580 43.710 153.645 43.710 153.645 43.690 ;
        RECT 153.645 43.690 155.870 43.710 ;
        RECT 117.285 43.680 152.470 43.690 ;
        RECT 117.285 43.655 151.000 43.680 ;
        POLYGON 151.000 43.680 151.010 43.680 151.010 43.675 ;
        RECT 151.010 43.675 152.470 43.680 ;
        POLYGON 152.470 43.690 152.500 43.675 152.470 43.675 ;
        POLYGON 153.645 43.690 153.700 43.690 153.700 43.675 ;
        RECT 153.700 43.675 155.870 43.690 ;
        POLYGON 151.000 43.675 151.010 43.655 151.000 43.655 ;
        RECT 117.285 43.615 151.010 43.655 ;
        POLYGON 151.010 43.675 151.050 43.675 151.050 43.650 ;
        RECT 151.050 43.660 152.505 43.675 ;
        POLYGON 152.505 43.675 152.540 43.660 152.505 43.660 ;
        POLYGON 153.705 43.675 153.735 43.675 153.735 43.670 ;
        RECT 153.735 43.670 155.870 43.675 ;
        POLYGON 153.735 43.670 153.775 43.670 153.775 43.660 ;
        RECT 153.775 43.660 155.870 43.670 ;
        RECT 151.050 43.650 152.540 43.660 ;
        POLYGON 117.285 43.615 117.295 43.615 117.295 43.340 ;
        RECT 117.295 43.570 151.010 43.615 ;
        POLYGON 151.010 43.650 151.050 43.570 151.010 43.570 ;
        POLYGON 151.050 43.650 151.175 43.650 151.175 43.570 ;
        RECT 151.175 43.610 152.540 43.650 ;
        POLYGON 152.540 43.660 152.690 43.610 152.540 43.610 ;
        POLYGON 153.775 43.660 153.915 43.660 153.915 43.625 ;
        RECT 153.915 43.655 155.870 43.660 ;
        POLYGON 155.870 43.710 156.085 43.710 155.870 43.655 ;
        POLYGON 157.375 43.710 157.375 43.705 157.365 43.705 ;
        RECT 157.375 43.705 158.550 43.710 ;
        POLYGON 157.365 43.705 157.365 43.685 157.315 43.685 ;
        RECT 157.365 43.685 158.550 43.705 ;
        POLYGON 157.310 43.685 157.310 43.655 157.235 43.655 ;
        RECT 157.310 43.655 158.550 43.685 ;
        RECT 153.915 43.650 155.855 43.655 ;
        POLYGON 155.855 43.655 155.870 43.655 155.855 43.650 ;
        POLYGON 157.235 43.655 157.235 43.650 157.220 43.650 ;
        RECT 157.235 43.650 158.550 43.655 ;
        RECT 153.915 43.645 155.830 43.650 ;
        POLYGON 155.830 43.650 155.850 43.650 155.830 43.645 ;
        POLYGON 157.220 43.650 157.220 43.645 157.210 43.645 ;
        RECT 157.220 43.645 158.550 43.650 ;
        RECT 153.915 43.625 155.660 43.645 ;
        POLYGON 153.915 43.625 153.995 43.625 153.995 43.610 ;
        RECT 153.995 43.610 155.660 43.625 ;
        POLYGON 155.660 43.645 155.830 43.645 155.660 43.610 ;
        POLYGON 157.210 43.645 157.210 43.630 157.170 43.630 ;
        RECT 157.210 43.635 158.550 43.645 ;
        POLYGON 158.550 43.765 158.765 43.765 158.550 43.635 ;
        POLYGON 159.940 43.765 159.940 43.635 159.785 43.635 ;
        RECT 159.940 43.710 160.975 43.765 ;
        POLYGON 160.975 43.960 161.210 43.960 160.975 43.710 ;
        POLYGON 162.450 43.960 162.450 43.945 162.440 43.945 ;
        RECT 162.450 43.945 164.010 43.960 ;
        POLYGON 162.440 43.945 162.440 43.910 162.410 43.910 ;
        RECT 162.440 43.930 164.010 43.945 ;
        POLYGON 164.010 44.030 164.065 44.030 164.010 43.930 ;
        POLYGON 165.750 44.030 165.750 43.930 165.700 43.930 ;
        RECT 165.750 43.940 168.050 44.030 ;
        POLYGON 168.050 44.420 168.240 44.420 168.050 43.940 ;
        POLYGON 171.180 44.420 171.180 43.940 171.045 43.940 ;
        RECT 171.180 44.045 175.575 44.420 ;
        POLYGON 175.575 45.765 175.685 45.765 175.575 44.045 ;
        POLYGON 182.900 45.625 182.900 44.210 182.810 44.210 ;
        RECT 182.900 44.610 197.880 45.765 ;
        POLYGON 197.880 46.405 198.000 44.610 197.880 44.610 ;
        POLYGON 207.785 46.405 207.930 46.405 207.930 45.845 ;
        RECT 207.930 45.845 222.755 46.405 ;
        POLYGON 207.930 45.845 207.980 45.845 207.980 45.700 ;
        RECT 207.980 45.700 222.755 45.845 ;
        POLYGON 207.980 45.700 208.330 45.700 208.330 44.610 ;
        RECT 208.330 45.640 222.755 45.700 ;
        POLYGON 222.755 46.405 222.965 45.640 222.755 45.640 ;
        POLYGON 229.810 46.405 229.910 46.405 229.910 46.020 ;
        RECT 229.910 46.020 233.880 46.405 ;
        POLYGON 229.910 46.020 229.930 46.020 229.930 45.945 ;
        RECT 229.930 46.005 233.880 46.020 ;
        POLYGON 233.880 46.405 234.010 46.005 233.880 46.005 ;
        POLYGON 236.675 46.405 236.725 46.405 236.725 46.265 ;
        RECT 236.725 46.265 238.690 46.405 ;
        POLYGON 236.725 46.265 236.800 46.265 236.800 46.035 ;
        RECT 236.800 46.180 238.690 46.265 ;
        POLYGON 238.690 46.405 238.775 46.180 238.690 46.180 ;
        POLYGON 240.265 46.405 240.325 46.405 240.325 46.265 ;
        RECT 240.325 46.385 241.425 46.405 ;
        POLYGON 241.425 46.465 241.465 46.385 241.425 46.385 ;
        POLYGON 242.450 46.465 242.485 46.465 242.485 46.405 ;
        RECT 242.485 46.460 243.285 46.465 ;
        POLYGON 243.285 46.490 243.300 46.460 243.285 46.460 ;
        POLYGON 243.980 46.490 244.000 46.490 244.000 46.460 ;
        RECT 242.485 46.405 243.300 46.460 ;
        RECT 244.000 46.455 244.605 46.490 ;
        POLYGON 243.300 46.455 243.330 46.405 243.300 46.405 ;
        POLYGON 244.000 46.455 244.015 46.455 244.015 46.435 ;
        RECT 244.015 46.435 244.605 46.455 ;
        POLYGON 244.015 46.435 244.030 46.435 244.030 46.410 ;
        RECT 244.030 46.415 244.605 46.435 ;
        POLYGON 244.605 46.535 244.695 46.415 244.605 46.415 ;
        POLYGON 245.115 46.535 245.165 46.535 245.165 46.465 ;
        RECT 245.165 46.495 246.025 46.535 ;
        POLYGON 246.025 46.610 246.130 46.495 246.025 46.495 ;
        POLYGON 253.620 46.610 253.620 46.495 253.505 46.495 ;
        RECT 253.620 46.495 254.525 46.610 ;
        RECT 245.165 46.465 246.130 46.495 ;
        POLYGON 245.165 46.465 245.190 46.465 245.190 46.435 ;
        RECT 245.190 46.450 246.130 46.465 ;
        POLYGON 246.130 46.495 246.175 46.450 246.130 46.450 ;
        RECT 245.190 46.435 246.175 46.450 ;
        POLYGON 253.505 46.495 253.505 46.445 253.455 46.445 ;
        RECT 253.505 46.445 254.525 46.495 ;
        POLYGON 254.525 46.700 254.705 46.700 254.525 46.445 ;
        POLYGON 255.240 46.700 255.240 46.695 255.235 46.695 ;
        RECT 255.240 46.695 255.695 46.705 ;
        POLYGON 255.235 46.695 255.235 46.600 255.175 46.600 ;
        RECT 255.235 46.625 255.695 46.695 ;
        POLYGON 255.695 46.750 255.765 46.750 255.695 46.625 ;
        POLYGON 256.385 46.745 256.385 46.680 256.355 46.680 ;
        RECT 256.385 46.740 257.100 46.750 ;
        POLYGON 257.100 46.935 257.175 46.935 257.100 46.740 ;
        POLYGON 257.990 46.935 257.990 46.890 257.975 46.890 ;
        RECT 257.990 46.890 258.925 46.935 ;
        POLYGON 257.975 46.890 257.975 46.845 257.955 46.845 ;
        RECT 257.975 46.845 258.925 46.890 ;
        POLYGON 257.955 46.845 257.955 46.740 257.915 46.740 ;
        RECT 257.955 46.775 258.925 46.845 ;
        POLYGON 258.925 46.935 258.975 46.935 258.925 46.775 ;
        POLYGON 260.240 46.935 260.240 46.870 260.225 46.870 ;
        RECT 260.240 46.870 261.790 46.935 ;
        POLYGON 260.225 46.870 260.225 46.780 260.205 46.780 ;
        RECT 260.225 46.780 261.790 46.870 ;
        RECT 257.955 46.740 258.830 46.775 ;
        RECT 256.385 46.680 256.995 46.740 ;
        POLYGON 256.355 46.680 256.355 46.630 256.330 46.630 ;
        RECT 256.355 46.630 256.995 46.680 ;
        RECT 255.235 46.600 255.655 46.625 ;
        POLYGON 255.175 46.600 255.175 46.585 255.160 46.585 ;
        RECT 255.175 46.585 255.655 46.600 ;
        POLYGON 255.160 46.585 255.160 46.545 255.135 46.545 ;
        RECT 255.160 46.555 255.655 46.585 ;
        POLYGON 255.655 46.625 255.695 46.625 255.655 46.555 ;
        POLYGON 256.330 46.625 256.330 46.555 256.295 46.555 ;
        RECT 256.330 46.555 256.995 46.630 ;
        RECT 255.160 46.545 255.560 46.555 ;
        POLYGON 255.135 46.545 255.135 46.475 255.085 46.475 ;
        RECT 255.135 46.475 255.560 46.545 ;
        POLYGON 255.085 46.475 255.085 46.445 255.065 46.445 ;
        RECT 255.085 46.445 255.560 46.475 ;
        POLYGON 245.190 46.435 245.205 46.435 245.205 46.415 ;
        RECT 245.205 46.415 246.175 46.435 ;
        RECT 244.030 46.405 244.695 46.415 ;
        POLYGON 244.695 46.415 244.700 46.405 244.695 46.405 ;
        POLYGON 245.205 46.415 245.210 46.415 245.210 46.405 ;
        RECT 245.210 46.405 246.175 46.415 ;
        POLYGON 242.485 46.405 242.495 46.405 242.495 46.385 ;
        RECT 242.495 46.385 243.330 46.405 ;
        RECT 240.325 46.290 241.465 46.385 ;
        POLYGON 241.465 46.385 241.510 46.290 241.465 46.290 ;
        POLYGON 242.495 46.385 242.525 46.385 242.525 46.335 ;
        RECT 242.525 46.360 243.330 46.385 ;
        POLYGON 243.330 46.405 243.360 46.360 243.330 46.360 ;
        POLYGON 244.030 46.405 244.060 46.405 244.060 46.360 ;
        RECT 244.060 46.385 244.700 46.405 ;
        POLYGON 244.700 46.405 244.720 46.385 244.700 46.385 ;
        POLYGON 245.210 46.405 245.225 46.405 245.225 46.390 ;
        RECT 245.225 46.385 246.175 46.405 ;
        RECT 244.060 46.365 244.720 46.385 ;
        POLYGON 244.720 46.385 244.735 46.365 244.720 46.365 ;
        POLYGON 245.225 46.385 245.240 46.385 245.240 46.370 ;
        RECT 245.240 46.365 246.175 46.385 ;
        RECT 244.060 46.360 244.735 46.365 ;
        RECT 242.525 46.330 243.360 46.360 ;
        POLYGON 243.360 46.360 243.375 46.330 243.360 46.330 ;
        POLYGON 244.060 46.360 244.080 46.360 244.080 46.330 ;
        RECT 244.080 46.330 244.735 46.360 ;
        POLYGON 242.525 46.330 242.545 46.330 242.545 46.290 ;
        RECT 242.545 46.300 243.375 46.330 ;
        POLYGON 243.375 46.330 243.395 46.300 243.375 46.300 ;
        POLYGON 244.080 46.330 244.100 46.330 244.100 46.300 ;
        RECT 244.100 46.300 244.735 46.330 ;
        RECT 240.325 46.285 241.510 46.290 ;
        POLYGON 241.510 46.290 241.515 46.285 241.510 46.285 ;
        RECT 242.545 46.285 243.395 46.300 ;
        RECT 240.325 46.265 241.515 46.285 ;
        POLYGON 241.515 46.285 241.525 46.265 241.515 46.265 ;
        POLYGON 242.545 46.285 242.560 46.285 242.560 46.265 ;
        POLYGON 240.325 46.265 240.330 46.265 240.330 46.255 ;
        RECT 240.330 46.255 241.525 46.265 ;
        RECT 242.560 46.260 243.395 46.285 ;
        POLYGON 241.525 46.260 241.530 46.255 241.525 46.255 ;
        POLYGON 242.560 46.260 242.565 46.260 242.565 46.255 ;
        RECT 242.565 46.255 243.395 46.260 ;
        POLYGON 240.330 46.255 240.360 46.255 240.360 46.185 ;
        RECT 240.360 46.215 241.530 46.255 ;
        POLYGON 241.530 46.255 241.550 46.215 241.530 46.215 ;
        POLYGON 242.565 46.255 242.585 46.255 242.585 46.220 ;
        RECT 242.585 46.215 243.395 46.255 ;
        RECT 240.360 46.200 241.550 46.215 ;
        POLYGON 241.550 46.215 241.560 46.200 241.550 46.200 ;
        POLYGON 242.585 46.215 242.595 46.215 242.595 46.200 ;
        RECT 242.595 46.200 243.395 46.215 ;
        POLYGON 243.395 46.300 243.455 46.200 243.395 46.200 ;
        POLYGON 244.100 46.300 244.130 46.300 244.130 46.265 ;
        RECT 244.130 46.265 244.735 46.300 ;
        POLYGON 244.130 46.265 244.170 46.265 244.170 46.205 ;
        RECT 244.170 46.210 244.735 46.265 ;
        POLYGON 244.735 46.365 244.855 46.210 244.735 46.210 ;
        POLYGON 245.240 46.365 245.335 46.365 245.335 46.245 ;
        RECT 245.335 46.295 246.175 46.365 ;
        POLYGON 246.175 46.445 246.325 46.295 246.175 46.295 ;
        POLYGON 253.455 46.445 253.455 46.405 253.410 46.405 ;
        RECT 253.455 46.440 254.525 46.445 ;
        RECT 253.455 46.405 254.495 46.440 ;
        POLYGON 254.495 46.440 254.525 46.440 254.495 46.405 ;
        POLYGON 255.065 46.445 255.065 46.405 255.035 46.405 ;
        RECT 255.065 46.405 255.560 46.445 ;
        POLYGON 255.560 46.555 255.655 46.555 255.560 46.405 ;
        POLYGON 256.295 46.555 256.295 46.505 256.270 46.505 ;
        RECT 256.295 46.510 256.995 46.555 ;
        POLYGON 256.995 46.740 257.100 46.740 256.995 46.510 ;
        POLYGON 257.915 46.740 257.915 46.625 257.870 46.625 ;
        RECT 257.915 46.625 258.830 46.740 ;
        POLYGON 257.870 46.625 257.870 46.510 257.820 46.510 ;
        RECT 257.870 46.510 258.830 46.625 ;
        POLYGON 258.830 46.775 258.925 46.775 258.830 46.510 ;
        POLYGON 260.205 46.775 260.205 46.715 260.190 46.715 ;
        RECT 260.205 46.715 261.790 46.780 ;
        POLYGON 260.190 46.715 260.190 46.520 260.140 46.520 ;
        RECT 260.190 46.700 261.790 46.715 ;
        POLYGON 261.790 46.935 261.835 46.935 261.790 46.700 ;
        POLYGON 263.875 46.940 263.875 46.935 263.870 46.935 ;
        RECT 263.875 46.935 266.630 46.965 ;
        POLYGON 266.630 47.030 266.645 47.030 266.630 46.935 ;
        POLYGON 263.870 46.925 263.870 46.710 263.835 46.710 ;
        RECT 263.870 46.920 266.630 46.935 ;
        RECT 263.870 46.710 266.570 46.920 ;
        RECT 260.190 46.565 261.760 46.700 ;
        POLYGON 261.760 46.700 261.790 46.700 261.760 46.565 ;
        POLYGON 263.835 46.700 263.835 46.680 263.830 46.680 ;
        RECT 263.835 46.680 266.570 46.710 ;
        POLYGON 263.830 46.680 263.830 46.615 263.820 46.615 ;
        RECT 263.830 46.615 266.570 46.680 ;
        POLYGON 263.820 46.615 263.820 46.565 263.810 46.565 ;
        RECT 263.820 46.565 266.570 46.615 ;
        RECT 260.190 46.520 261.735 46.565 ;
        RECT 256.295 46.505 256.985 46.510 ;
        POLYGON 256.270 46.505 256.270 46.500 256.265 46.500 ;
        RECT 256.270 46.500 256.985 46.505 ;
        POLYGON 256.265 46.500 256.265 46.460 256.245 46.460 ;
        RECT 256.265 46.475 256.985 46.500 ;
        POLYGON 256.985 46.510 256.995 46.510 256.985 46.475 ;
        POLYGON 257.820 46.510 257.820 46.485 257.810 46.485 ;
        RECT 257.820 46.485 258.820 46.510 ;
        POLYGON 257.810 46.485 257.810 46.475 257.805 46.475 ;
        RECT 257.810 46.475 258.820 46.485 ;
        POLYGON 258.820 46.510 258.830 46.510 258.820 46.475 ;
        POLYGON 260.140 46.510 260.140 46.480 260.130 46.480 ;
        RECT 260.140 46.480 261.735 46.520 ;
        RECT 256.265 46.470 256.980 46.475 ;
        POLYGON 256.980 46.475 256.985 46.475 256.980 46.470 ;
        RECT 256.265 46.460 256.950 46.470 ;
        POLYGON 256.245 46.460 256.245 46.405 256.215 46.405 ;
        RECT 256.245 46.405 256.950 46.460 ;
        POLYGON 256.950 46.470 256.980 46.470 256.950 46.410 ;
        POLYGON 257.805 46.470 257.805 46.450 257.795 46.450 ;
        RECT 257.805 46.450 258.795 46.475 ;
        POLYGON 257.795 46.450 257.795 46.415 257.780 46.415 ;
        RECT 257.795 46.415 258.795 46.450 ;
        POLYGON 253.410 46.405 253.410 46.380 253.385 46.380 ;
        RECT 253.410 46.380 254.445 46.405 ;
        POLYGON 253.385 46.380 253.385 46.295 253.295 46.295 ;
        RECT 253.385 46.340 254.445 46.380 ;
        POLYGON 254.445 46.405 254.495 46.405 254.445 46.340 ;
        POLYGON 255.035 46.405 255.035 46.340 254.985 46.340 ;
        RECT 255.035 46.340 255.495 46.405 ;
        RECT 253.385 46.295 254.310 46.340 ;
        RECT 245.335 46.270 246.325 46.295 ;
        POLYGON 246.325 46.295 246.355 46.270 246.325 46.270 ;
        POLYGON 253.295 46.295 253.295 46.270 253.270 46.270 ;
        RECT 253.295 46.270 254.310 46.295 ;
        RECT 245.335 46.245 246.355 46.270 ;
        POLYGON 245.335 46.245 245.365 46.245 245.365 46.215 ;
        RECT 245.365 46.220 246.355 46.245 ;
        POLYGON 246.355 46.270 246.405 46.220 246.355 46.220 ;
        POLYGON 253.270 46.270 253.270 46.250 253.245 46.250 ;
        RECT 253.270 46.250 254.310 46.270 ;
        POLYGON 253.245 46.250 253.245 46.220 253.215 46.220 ;
        RECT 253.245 46.220 254.310 46.250 ;
        RECT 245.365 46.210 246.405 46.220 ;
        RECT 244.170 46.200 244.855 46.210 ;
        RECT 240.360 46.180 241.560 46.200 ;
        RECT 236.800 46.140 238.775 46.180 ;
        POLYGON 238.775 46.180 238.795 46.140 238.775 46.140 ;
        POLYGON 240.360 46.180 240.380 46.180 240.380 46.145 ;
        RECT 240.380 46.145 241.560 46.180 ;
        POLYGON 241.560 46.200 241.590 46.145 241.560 46.145 ;
        POLYGON 242.595 46.200 242.605 46.200 242.605 46.185 ;
        RECT 242.605 46.190 243.455 46.200 ;
        POLYGON 243.455 46.200 243.460 46.190 243.455 46.190 ;
        POLYGON 244.170 46.200 244.180 46.200 244.180 46.190 ;
        RECT 244.180 46.190 244.855 46.200 ;
        POLYGON 244.855 46.210 244.875 46.190 244.855 46.190 ;
        POLYGON 245.365 46.210 245.385 46.210 245.385 46.190 ;
        RECT 245.385 46.190 246.405 46.210 ;
        RECT 242.605 46.185 243.460 46.190 ;
        POLYGON 242.605 46.185 242.625 46.185 242.625 46.150 ;
        RECT 242.625 46.145 243.460 46.185 ;
        RECT 240.380 46.140 241.590 46.145 ;
        RECT 236.800 46.035 238.795 46.140 ;
        POLYGON 236.800 46.035 236.810 46.035 236.810 46.005 ;
        RECT 236.810 46.005 238.795 46.035 ;
        RECT 229.930 45.945 234.010 46.005 ;
        POLYGON 229.930 45.945 230.015 45.945 230.015 45.645 ;
        RECT 230.015 45.770 234.010 45.945 ;
        POLYGON 234.010 46.005 234.080 45.770 234.010 45.770 ;
        POLYGON 236.810 46.005 236.900 46.005 236.900 45.775 ;
        RECT 236.900 45.770 238.795 46.005 ;
        RECT 230.015 45.725 234.080 45.770 ;
        POLYGON 234.080 45.770 234.095 45.725 234.080 45.725 ;
        POLYGON 236.900 45.770 236.920 45.770 236.920 45.725 ;
        RECT 236.920 45.740 238.795 45.770 ;
        POLYGON 238.795 46.140 238.965 45.740 238.795 45.740 ;
        POLYGON 240.380 46.140 240.460 46.140 240.460 45.970 ;
        RECT 240.460 46.070 241.590 46.140 ;
        POLYGON 241.590 46.145 241.630 46.070 241.590 46.070 ;
        POLYGON 242.625 46.145 242.675 46.145 242.675 46.070 ;
        RECT 242.675 46.085 243.460 46.145 ;
        POLYGON 243.460 46.190 243.530 46.085 243.460 46.085 ;
        POLYGON 244.180 46.190 244.240 46.190 244.240 46.105 ;
        RECT 244.240 46.105 244.875 46.190 ;
        POLYGON 244.240 46.105 244.250 46.105 244.250 46.090 ;
        RECT 244.250 46.085 244.875 46.105 ;
        RECT 242.675 46.070 243.530 46.085 ;
        RECT 240.460 46.045 241.630 46.070 ;
        POLYGON 241.630 46.070 241.645 46.045 241.630 46.045 ;
        POLYGON 242.675 46.070 242.685 46.070 242.685 46.055 ;
        RECT 242.685 46.055 243.530 46.070 ;
        POLYGON 242.685 46.055 242.690 46.055 242.690 46.045 ;
        RECT 242.690 46.050 243.530 46.055 ;
        POLYGON 243.530 46.085 243.555 46.050 243.530 46.050 ;
        POLYGON 244.250 46.085 244.265 46.085 244.265 46.070 ;
        RECT 244.265 46.070 244.875 46.085 ;
        POLYGON 244.265 46.070 244.280 46.070 244.280 46.050 ;
        RECT 244.280 46.050 244.875 46.070 ;
        RECT 242.690 46.045 243.555 46.050 ;
        RECT 240.460 45.970 241.645 46.045 ;
        POLYGON 240.460 45.970 240.530 45.970 240.530 45.825 ;
        RECT 240.530 45.925 241.645 45.970 ;
        POLYGON 241.645 46.045 241.710 45.925 241.645 45.925 ;
        POLYGON 242.690 46.045 242.765 46.045 242.765 45.925 ;
        RECT 242.765 45.950 243.555 46.045 ;
        POLYGON 243.555 46.050 243.620 45.950 243.555 45.950 ;
        POLYGON 244.280 46.050 244.350 46.050 244.350 45.960 ;
        RECT 244.350 46.035 244.875 46.050 ;
        POLYGON 244.875 46.190 245.005 46.035 244.875 46.035 ;
        POLYGON 245.385 46.190 245.415 46.190 245.415 46.155 ;
        RECT 245.415 46.155 246.405 46.190 ;
        POLYGON 245.415 46.155 245.520 46.155 245.520 46.035 ;
        RECT 245.520 46.150 246.405 46.155 ;
        POLYGON 246.405 46.220 246.485 46.150 246.405 46.150 ;
        POLYGON 253.215 46.220 253.215 46.150 253.130 46.150 ;
        RECT 253.215 46.170 254.310 46.220 ;
        POLYGON 254.310 46.340 254.445 46.340 254.310 46.170 ;
        POLYGON 254.985 46.340 254.985 46.315 254.965 46.315 ;
        RECT 254.985 46.315 255.495 46.340 ;
        POLYGON 254.965 46.315 254.965 46.255 254.920 46.255 ;
        RECT 254.965 46.300 255.495 46.315 ;
        POLYGON 255.495 46.405 255.560 46.405 255.495 46.305 ;
        POLYGON 256.215 46.400 256.215 46.325 256.175 46.325 ;
        RECT 256.215 46.325 256.855 46.405 ;
        POLYGON 256.175 46.325 256.175 46.310 256.165 46.310 ;
        RECT 256.175 46.310 256.855 46.325 ;
        POLYGON 256.165 46.305 256.165 46.300 256.160 46.300 ;
        RECT 256.165 46.300 256.855 46.310 ;
        RECT 254.965 46.280 255.480 46.300 ;
        POLYGON 255.480 46.300 255.495 46.300 255.480 46.280 ;
        POLYGON 256.160 46.300 256.160 46.285 256.150 46.285 ;
        RECT 256.160 46.285 256.855 46.300 ;
        RECT 254.965 46.255 255.320 46.280 ;
        POLYGON 254.920 46.255 254.920 46.250 254.915 46.250 ;
        RECT 254.920 46.250 255.320 46.255 ;
        POLYGON 254.915 46.250 254.915 46.170 254.850 46.170 ;
        RECT 254.915 46.170 255.320 46.250 ;
        RECT 253.215 46.160 254.305 46.170 ;
        POLYGON 254.305 46.170 254.310 46.170 254.305 46.160 ;
        POLYGON 254.850 46.170 254.850 46.160 254.840 46.160 ;
        RECT 254.850 46.160 255.320 46.170 ;
        RECT 253.215 46.150 254.185 46.160 ;
        RECT 245.520 46.105 246.485 46.150 ;
        POLYGON 246.485 46.150 246.535 46.105 246.485 46.105 ;
        POLYGON 253.130 46.150 253.130 46.120 253.095 46.120 ;
        RECT 253.130 46.120 254.185 46.150 ;
        POLYGON 253.095 46.120 253.095 46.105 253.080 46.105 ;
        RECT 253.095 46.105 254.185 46.120 ;
        RECT 245.520 46.035 246.535 46.105 ;
        RECT 244.350 46.015 245.005 46.035 ;
        POLYGON 245.005 46.035 245.025 46.015 245.005 46.015 ;
        RECT 244.350 45.995 245.025 46.015 ;
        POLYGON 245.520 46.035 245.540 46.035 245.540 46.010 ;
        RECT 245.540 46.015 246.535 46.035 ;
        POLYGON 246.535 46.105 246.645 46.015 246.535 46.015 ;
        POLYGON 253.080 46.105 253.080 46.090 253.060 46.090 ;
        RECT 253.080 46.090 254.185 46.105 ;
        POLYGON 253.060 46.090 253.060 46.030 252.985 46.030 ;
        RECT 253.060 46.030 254.185 46.090 ;
        POLYGON 254.185 46.160 254.305 46.160 254.185 46.030 ;
        POLYGON 254.840 46.160 254.840 46.080 254.775 46.080 ;
        RECT 254.840 46.080 255.320 46.160 ;
        POLYGON 254.775 46.080 254.775 46.030 254.730 46.030 ;
        RECT 254.775 46.055 255.320 46.080 ;
        POLYGON 255.320 46.280 255.480 46.280 255.320 46.055 ;
        POLYGON 256.150 46.280 256.150 46.145 256.070 46.145 ;
        RECT 256.150 46.210 256.855 46.285 ;
        POLYGON 256.855 46.405 256.950 46.405 256.855 46.210 ;
        POLYGON 257.780 46.410 257.780 46.405 257.775 46.405 ;
        RECT 257.780 46.405 258.795 46.415 ;
        POLYGON 258.795 46.475 258.820 46.475 258.795 46.410 ;
        POLYGON 260.130 46.475 260.130 46.460 260.125 46.460 ;
        RECT 260.130 46.460 261.735 46.480 ;
        POLYGON 260.125 46.460 260.125 46.410 260.110 46.410 ;
        RECT 260.125 46.445 261.735 46.460 ;
        POLYGON 261.735 46.565 261.760 46.565 261.735 46.445 ;
        POLYGON 263.810 46.565 263.810 46.445 263.785 46.445 ;
        RECT 263.810 46.445 266.570 46.565 ;
        POLYGON 266.570 46.920 266.630 46.920 266.570 46.445 ;
        POLYGON 270.685 46.935 270.685 46.445 270.680 46.445 ;
        RECT 270.685 46.780 277.910 47.075 ;
        POLYGON 287.930 47.030 287.930 46.970 287.925 46.970 ;
        RECT 287.930 46.970 303.120 51.515 ;
        POLYGON 277.910 46.935 277.915 46.780 277.910 46.780 ;
        RECT 270.685 46.445 277.905 46.780 ;
        RECT 260.125 46.410 261.725 46.445 ;
        POLYGON 261.725 46.445 261.735 46.445 261.725 46.410 ;
        POLYGON 263.785 46.445 263.785 46.420 263.780 46.420 ;
        RECT 263.785 46.420 266.565 46.445 ;
        RECT 260.110 46.405 261.725 46.410 ;
        POLYGON 257.775 46.400 257.775 46.295 257.730 46.295 ;
        RECT 257.775 46.395 258.790 46.405 ;
        POLYGON 258.790 46.405 258.795 46.405 258.790 46.395 ;
        POLYGON 260.110 46.405 260.110 46.395 260.105 46.395 ;
        RECT 260.110 46.395 261.665 46.405 ;
        RECT 257.775 46.295 258.705 46.395 ;
        POLYGON 257.730 46.295 257.730 46.210 257.690 46.210 ;
        RECT 257.730 46.210 258.705 46.295 ;
        RECT 256.150 46.145 256.765 46.210 ;
        POLYGON 256.070 46.145 256.070 46.130 256.065 46.130 ;
        RECT 256.070 46.130 256.765 46.145 ;
        POLYGON 256.065 46.130 256.065 46.055 256.020 46.055 ;
        RECT 256.065 46.055 256.765 46.130 ;
        RECT 254.775 46.030 255.290 46.055 ;
        POLYGON 252.985 46.030 252.985 46.015 252.965 46.015 ;
        RECT 252.985 46.015 254.095 46.030 ;
        RECT 245.540 46.010 246.645 46.015 ;
        POLYGON 245.025 46.010 245.040 45.995 245.025 45.995 ;
        POLYGON 245.540 46.010 245.555 46.010 245.555 45.995 ;
        RECT 245.555 46.005 246.645 46.010 ;
        POLYGON 246.645 46.015 246.650 46.005 246.645 46.005 ;
        POLYGON 252.965 46.015 252.965 46.005 252.955 46.005 ;
        RECT 252.965 46.005 254.095 46.015 ;
        RECT 245.555 45.995 246.650 46.005 ;
        RECT 244.350 45.960 245.040 45.995 ;
        POLYGON 244.350 45.960 244.355 45.960 244.355 45.950 ;
        RECT 244.355 45.950 245.040 45.960 ;
        RECT 242.765 45.935 243.620 45.950 ;
        POLYGON 243.620 45.950 243.630 45.935 243.620 45.935 ;
        POLYGON 244.355 45.950 244.365 45.950 244.365 45.940 ;
        RECT 244.365 45.935 245.040 45.950 ;
        RECT 242.765 45.925 243.630 45.935 ;
        RECT 240.530 45.915 241.710 45.925 ;
        POLYGON 241.710 45.925 241.715 45.915 241.710 45.915 ;
        POLYGON 242.765 45.925 242.770 45.925 242.770 45.915 ;
        RECT 242.770 45.915 243.630 45.925 ;
        RECT 240.530 45.895 241.715 45.915 ;
        POLYGON 241.715 45.915 241.730 45.895 241.715 45.895 ;
        POLYGON 242.770 45.915 242.780 45.915 242.780 45.900 ;
        RECT 242.780 45.905 243.630 45.915 ;
        POLYGON 243.630 45.935 243.655 45.905 243.630 45.905 ;
        POLYGON 244.365 45.935 244.385 45.935 244.385 45.915 ;
        RECT 244.385 45.915 245.040 45.935 ;
        POLYGON 244.385 45.915 244.390 45.915 244.390 45.905 ;
        RECT 244.390 45.905 245.040 45.915 ;
        RECT 242.780 45.895 243.655 45.905 ;
        RECT 240.530 45.825 241.730 45.895 ;
        POLYGON 240.530 45.825 240.570 45.825 240.570 45.745 ;
        RECT 240.570 45.795 241.730 45.825 ;
        POLYGON 241.730 45.895 241.790 45.795 241.730 45.795 ;
        POLYGON 242.780 45.895 242.845 45.895 242.845 45.795 ;
        RECT 242.845 45.795 243.655 45.895 ;
        RECT 240.570 45.740 241.790 45.795 ;
        RECT 236.920 45.725 238.965 45.740 ;
        RECT 208.330 45.400 222.965 45.640 ;
        RECT 230.015 45.630 234.095 45.725 ;
        POLYGON 222.965 45.630 223.035 45.400 222.965 45.400 ;
        POLYGON 230.015 45.630 230.085 45.630 230.085 45.400 ;
        RECT 230.085 45.400 234.095 45.630 ;
        RECT 208.330 44.740 223.035 45.400 ;
        POLYGON 223.035 45.400 223.235 44.740 223.035 44.740 ;
        POLYGON 230.085 45.400 230.115 45.400 230.115 45.290 ;
        RECT 230.115 45.290 234.095 45.400 ;
        POLYGON 230.115 45.290 230.285 45.290 230.285 44.760 ;
        RECT 230.285 44.965 234.095 45.290 ;
        POLYGON 234.095 45.725 234.380 44.965 234.095 44.965 ;
        POLYGON 236.920 45.725 237.005 45.725 237.005 45.510 ;
        RECT 237.005 45.695 238.965 45.725 ;
        POLYGON 238.965 45.740 238.980 45.695 238.965 45.695 ;
        POLYGON 240.570 45.740 240.595 45.740 240.595 45.695 ;
        RECT 240.595 45.695 241.790 45.740 ;
        RECT 237.005 45.510 238.980 45.695 ;
        POLYGON 237.005 45.510 237.025 45.510 237.025 45.465 ;
        RECT 237.025 45.465 238.980 45.510 ;
        POLYGON 237.025 45.465 237.085 45.465 237.085 45.315 ;
        RECT 237.085 45.395 238.980 45.465 ;
        POLYGON 238.980 45.695 239.125 45.395 238.980 45.395 ;
        POLYGON 240.595 45.695 240.600 45.695 240.600 45.685 ;
        RECT 240.600 45.690 241.790 45.695 ;
        POLYGON 241.790 45.795 241.855 45.690 241.790 45.690 ;
        POLYGON 242.845 45.795 242.850 45.795 242.850 45.790 ;
        RECT 242.850 45.790 243.655 45.795 ;
        POLYGON 242.850 45.790 242.880 45.790 242.880 45.745 ;
        RECT 242.880 45.785 243.655 45.790 ;
        POLYGON 243.655 45.905 243.735 45.785 243.655 45.785 ;
        POLYGON 244.390 45.905 244.410 45.905 244.410 45.880 ;
        RECT 244.410 45.880 245.040 45.905 ;
        POLYGON 244.410 45.880 244.485 45.880 244.485 45.785 ;
        RECT 244.485 45.865 245.040 45.880 ;
        POLYGON 245.040 45.995 245.165 45.865 245.040 45.865 ;
        POLYGON 245.555 45.995 245.615 45.995 245.615 45.935 ;
        RECT 245.615 45.985 246.650 45.995 ;
        POLYGON 246.650 46.005 246.675 45.985 246.650 45.985 ;
        POLYGON 252.955 46.005 252.955 45.995 252.940 45.995 ;
        RECT 252.955 45.995 254.095 46.005 ;
        POLYGON 252.940 45.995 252.940 45.985 252.930 45.985 ;
        RECT 252.940 45.985 254.095 45.995 ;
        RECT 245.615 45.935 246.675 45.985 ;
        POLYGON 245.615 45.935 245.680 45.935 245.680 45.865 ;
        RECT 245.680 45.875 246.675 45.935 ;
        POLYGON 246.675 45.985 246.820 45.875 246.675 45.875 ;
        POLYGON 252.930 45.985 252.930 45.955 252.895 45.955 ;
        RECT 252.930 45.955 254.095 45.985 ;
        POLYGON 252.895 45.955 252.895 45.905 252.820 45.905 ;
        RECT 252.895 45.930 254.095 45.955 ;
        POLYGON 254.095 46.030 254.185 46.030 254.095 45.930 ;
        POLYGON 254.730 46.030 254.730 46.000 254.705 46.000 ;
        RECT 254.730 46.010 255.290 46.030 ;
        POLYGON 255.290 46.055 255.320 46.055 255.290 46.010 ;
        POLYGON 256.020 46.055 256.020 46.010 255.990 46.010 ;
        RECT 256.020 46.045 256.765 46.055 ;
        POLYGON 256.765 46.210 256.855 46.210 256.765 46.045 ;
        POLYGON 257.690 46.205 257.690 46.185 257.680 46.185 ;
        RECT 257.690 46.185 258.705 46.210 ;
        POLYGON 257.680 46.185 257.680 46.170 257.670 46.170 ;
        RECT 257.680 46.175 258.705 46.185 ;
        POLYGON 258.705 46.395 258.790 46.395 258.705 46.175 ;
        POLYGON 260.105 46.390 260.105 46.370 260.100 46.370 ;
        RECT 260.105 46.370 261.665 46.395 ;
        POLYGON 260.100 46.370 260.100 46.295 260.080 46.295 ;
        RECT 260.100 46.295 261.665 46.370 ;
        POLYGON 260.080 46.295 260.080 46.215 260.055 46.215 ;
        RECT 260.080 46.215 261.665 46.295 ;
        POLYGON 260.055 46.215 260.055 46.185 260.045 46.185 ;
        RECT 260.055 46.190 261.665 46.215 ;
        POLYGON 261.665 46.405 261.725 46.405 261.665 46.190 ;
        POLYGON 263.780 46.410 263.780 46.405 263.775 46.405 ;
        RECT 263.780 46.405 266.565 46.420 ;
        POLYGON 266.565 46.445 266.570 46.445 266.565 46.415 ;
        POLYGON 263.775 46.395 263.775 46.195 263.735 46.195 ;
        RECT 263.775 46.195 266.475 46.405 ;
        RECT 260.055 46.185 261.580 46.190 ;
        RECT 257.680 46.170 258.580 46.175 ;
        POLYGON 257.670 46.170 257.670 46.135 257.655 46.135 ;
        RECT 257.670 46.135 258.580 46.170 ;
        POLYGON 257.655 46.135 257.655 46.070 257.625 46.070 ;
        RECT 257.655 46.070 258.580 46.135 ;
        POLYGON 257.625 46.070 257.625 46.045 257.615 46.045 ;
        RECT 257.625 46.045 258.580 46.070 ;
        RECT 256.020 46.020 256.755 46.045 ;
        POLYGON 256.755 46.045 256.765 46.045 256.755 46.020 ;
        POLYGON 257.615 46.045 257.615 46.025 257.605 46.025 ;
        RECT 257.615 46.025 258.580 46.045 ;
        RECT 256.020 46.010 256.715 46.020 ;
        RECT 254.730 46.000 255.175 46.010 ;
        POLYGON 254.705 46.000 254.705 45.930 254.640 45.930 ;
        RECT 254.705 45.930 255.175 46.000 ;
        RECT 252.895 45.905 254.065 45.930 ;
        POLYGON 252.820 45.905 252.820 45.875 252.785 45.875 ;
        RECT 252.820 45.895 254.065 45.905 ;
        POLYGON 254.065 45.930 254.095 45.930 254.065 45.895 ;
        POLYGON 254.640 45.930 254.640 45.895 254.605 45.895 ;
        RECT 254.640 45.895 255.175 45.930 ;
        RECT 252.820 45.875 253.935 45.895 ;
        RECT 245.680 45.865 246.820 45.875 ;
        POLYGON 246.820 45.875 246.830 45.865 246.820 45.865 ;
        POLYGON 252.785 45.875 252.785 45.865 252.770 45.865 ;
        RECT 252.785 45.865 253.935 45.875 ;
        RECT 244.485 45.840 245.165 45.865 ;
        POLYGON 245.165 45.865 245.190 45.840 245.165 45.840 ;
        POLYGON 245.680 45.865 245.705 45.865 245.705 45.840 ;
        RECT 245.705 45.840 246.830 45.865 ;
        RECT 244.485 45.800 245.190 45.840 ;
        POLYGON 245.190 45.840 245.225 45.800 245.190 45.800 ;
        POLYGON 245.705 45.840 245.715 45.840 245.715 45.830 ;
        RECT 245.715 45.830 246.830 45.840 ;
        POLYGON 245.715 45.830 245.750 45.830 245.750 45.800 ;
        RECT 245.750 45.825 246.830 45.830 ;
        POLYGON 246.830 45.865 246.890 45.825 246.830 45.825 ;
        POLYGON 252.770 45.865 252.770 45.830 252.725 45.830 ;
        RECT 252.770 45.830 253.935 45.865 ;
        POLYGON 252.725 45.830 252.725 45.825 252.720 45.825 ;
        RECT 252.725 45.825 253.935 45.830 ;
        RECT 245.750 45.800 246.890 45.825 ;
        RECT 244.485 45.785 245.225 45.800 ;
        RECT 242.880 45.755 243.735 45.785 ;
        POLYGON 243.735 45.785 243.760 45.755 243.735 45.755 ;
        POLYGON 244.485 45.785 244.510 45.785 244.510 45.755 ;
        RECT 244.510 45.755 245.225 45.785 ;
        RECT 242.880 45.745 243.760 45.755 ;
        POLYGON 242.880 45.745 242.915 45.745 242.915 45.690 ;
        RECT 242.915 45.705 243.760 45.745 ;
        POLYGON 243.760 45.755 243.795 45.705 243.760 45.705 ;
        POLYGON 244.510 45.755 244.535 45.755 244.535 45.725 ;
        RECT 244.535 45.725 245.225 45.755 ;
        POLYGON 244.535 45.725 244.555 45.725 244.555 45.705 ;
        RECT 244.555 45.705 245.225 45.725 ;
        RECT 242.915 45.690 243.795 45.705 ;
        RECT 240.600 45.685 241.855 45.690 ;
        POLYGON 240.600 45.685 240.755 45.685 240.755 45.395 ;
        RECT 240.755 45.645 241.855 45.685 ;
        POLYGON 241.855 45.690 241.885 45.645 241.855 45.645 ;
        POLYGON 242.915 45.690 242.945 45.690 242.945 45.645 ;
        RECT 242.945 45.645 243.795 45.690 ;
        RECT 240.755 45.565 241.885 45.645 ;
        POLYGON 241.885 45.645 241.930 45.565 241.885 45.565 ;
        POLYGON 242.945 45.645 243.000 45.645 243.000 45.565 ;
        RECT 243.000 45.635 243.795 45.645 ;
        POLYGON 243.795 45.705 243.850 45.635 243.795 45.635 ;
        POLYGON 244.555 45.705 244.565 45.705 244.565 45.695 ;
        RECT 244.565 45.695 245.225 45.705 ;
        POLYGON 244.565 45.695 244.615 45.695 244.615 45.635 ;
        RECT 244.615 45.685 245.225 45.695 ;
        POLYGON 245.225 45.800 245.335 45.685 245.225 45.685 ;
        POLYGON 245.750 45.800 245.865 45.800 245.865 45.685 ;
        RECT 245.865 45.770 246.890 45.800 ;
        POLYGON 246.890 45.825 246.965 45.770 246.890 45.770 ;
        POLYGON 252.720 45.825 252.720 45.810 252.695 45.810 ;
        RECT 252.720 45.810 253.935 45.825 ;
        POLYGON 252.695 45.810 252.695 45.800 252.675 45.800 ;
        RECT 252.695 45.800 253.935 45.810 ;
        POLYGON 252.675 45.800 252.675 45.770 252.630 45.770 ;
        RECT 252.675 45.770 253.935 45.800 ;
        RECT 245.865 45.685 246.965 45.770 ;
        RECT 244.615 45.660 245.335 45.685 ;
        POLYGON 245.335 45.685 245.355 45.660 245.335 45.660 ;
        POLYGON 245.865 45.685 245.890 45.685 245.890 45.660 ;
        RECT 245.890 45.670 246.965 45.685 ;
        POLYGON 246.965 45.770 247.115 45.670 246.965 45.670 ;
        POLYGON 252.630 45.770 252.630 45.765 252.625 45.765 ;
        RECT 252.630 45.765 253.935 45.770 ;
        POLYGON 253.935 45.895 254.065 45.895 253.935 45.765 ;
        POLYGON 254.605 45.895 254.605 45.805 254.525 45.805 ;
        RECT 254.605 45.860 255.175 45.895 ;
        POLYGON 255.175 46.010 255.290 46.010 255.175 45.860 ;
        POLYGON 255.990 46.010 255.990 45.930 255.940 45.930 ;
        RECT 255.990 45.950 256.715 46.010 ;
        POLYGON 256.715 46.020 256.755 46.020 256.715 45.950 ;
        POLYGON 257.605 46.020 257.605 45.985 257.585 45.985 ;
        RECT 257.605 45.985 258.580 46.025 ;
        POLYGON 257.585 45.985 257.585 45.965 257.575 45.965 ;
        RECT 257.585 45.965 258.580 45.985 ;
        POLYGON 257.575 45.965 257.575 45.950 257.565 45.950 ;
        RECT 257.575 45.950 258.580 45.965 ;
        RECT 255.990 45.930 256.570 45.950 ;
        POLYGON 255.940 45.930 255.940 45.915 255.930 45.915 ;
        RECT 255.940 45.915 256.570 45.930 ;
        POLYGON 255.930 45.915 255.930 45.865 255.895 45.865 ;
        RECT 255.930 45.865 256.570 45.915 ;
        RECT 254.605 45.810 255.135 45.860 ;
        POLYGON 255.135 45.860 255.175 45.860 255.135 45.810 ;
        POLYGON 255.895 45.860 255.895 45.855 255.890 45.855 ;
        RECT 255.895 45.855 256.570 45.865 ;
        POLYGON 255.890 45.855 255.890 45.810 255.860 45.810 ;
        RECT 255.890 45.810 256.570 45.855 ;
        RECT 254.605 45.805 255.070 45.810 ;
        POLYGON 254.525 45.805 254.525 45.765 254.485 45.765 ;
        RECT 254.525 45.765 255.070 45.805 ;
        POLYGON 252.625 45.765 252.625 45.715 252.550 45.715 ;
        RECT 252.625 45.750 253.925 45.765 ;
        POLYGON 253.925 45.765 253.935 45.765 253.925 45.750 ;
        POLYGON 254.485 45.765 254.485 45.750 254.470 45.750 ;
        RECT 254.485 45.750 255.070 45.765 ;
        RECT 252.625 45.715 253.870 45.750 ;
        POLYGON 252.550 45.715 252.550 45.700 252.525 45.700 ;
        RECT 252.550 45.700 253.870 45.715 ;
        POLYGON 253.870 45.750 253.920 45.750 253.870 45.700 ;
        POLYGON 254.470 45.750 254.470 45.720 254.445 45.720 ;
        RECT 254.470 45.735 255.070 45.750 ;
        POLYGON 255.070 45.810 255.135 45.810 255.070 45.735 ;
        POLYGON 255.860 45.810 255.860 45.735 255.810 45.735 ;
        RECT 255.860 45.735 256.570 45.810 ;
        RECT 254.470 45.720 254.940 45.735 ;
        POLYGON 254.445 45.720 254.445 45.700 254.425 45.700 ;
        RECT 254.445 45.700 254.940 45.720 ;
        POLYGON 252.525 45.700 252.525 45.670 252.480 45.670 ;
        RECT 252.525 45.670 253.805 45.700 ;
        RECT 245.890 45.660 247.115 45.670 ;
        RECT 244.615 45.655 245.355 45.660 ;
        POLYGON 245.355 45.660 245.365 45.655 245.355 45.655 ;
        POLYGON 245.890 45.660 245.895 45.660 245.895 45.655 ;
        RECT 245.895 45.655 247.115 45.660 ;
        RECT 244.615 45.635 245.365 45.655 ;
        RECT 243.000 45.605 243.850 45.635 ;
        POLYGON 243.850 45.635 243.875 45.605 243.850 45.605 ;
        POLYGON 244.615 45.635 244.640 45.635 244.640 45.605 ;
        RECT 244.640 45.605 245.365 45.635 ;
        POLYGON 245.365 45.655 245.415 45.605 245.365 45.605 ;
        POLYGON 245.895 45.655 245.955 45.655 245.955 45.610 ;
        RECT 245.955 45.650 247.115 45.655 ;
        POLYGON 247.115 45.670 247.150 45.650 247.115 45.650 ;
        POLYGON 252.480 45.670 252.480 45.655 252.460 45.655 ;
        RECT 252.480 45.655 253.805 45.670 ;
        POLYGON 252.460 45.655 252.460 45.650 252.450 45.650 ;
        RECT 252.460 45.650 253.805 45.655 ;
        RECT 245.955 45.635 247.150 45.650 ;
        POLYGON 247.150 45.650 247.175 45.635 247.150 45.635 ;
        POLYGON 252.450 45.650 252.450 45.635 252.430 45.635 ;
        RECT 252.450 45.640 253.805 45.650 ;
        POLYGON 253.805 45.700 253.870 45.700 253.805 45.640 ;
        POLYGON 254.425 45.700 254.425 45.640 254.360 45.640 ;
        RECT 254.425 45.640 254.940 45.700 ;
        RECT 252.450 45.635 253.670 45.640 ;
        RECT 245.955 45.610 247.175 45.635 ;
        POLYGON 245.955 45.610 245.960 45.610 245.960 45.605 ;
        RECT 245.960 45.605 247.175 45.610 ;
        RECT 243.000 45.565 243.875 45.605 ;
        RECT 240.755 45.480 241.930 45.565 ;
        POLYGON 241.930 45.565 241.990 45.480 241.930 45.480 ;
        POLYGON 243.000 45.565 243.040 45.565 243.040 45.510 ;
        RECT 243.040 45.510 243.875 45.565 ;
        POLYGON 243.040 45.510 243.060 45.510 243.060 45.480 ;
        RECT 243.060 45.480 243.875 45.510 ;
        POLYGON 243.875 45.605 243.975 45.480 243.875 45.480 ;
        POLYGON 244.640 45.605 244.695 45.605 244.695 45.545 ;
        RECT 244.695 45.545 245.415 45.605 ;
        POLYGON 244.695 45.545 244.725 45.545 244.725 45.515 ;
        RECT 244.725 45.515 245.415 45.545 ;
        POLYGON 244.725 45.515 244.755 45.515 244.755 45.480 ;
        RECT 244.755 45.510 245.415 45.515 ;
        POLYGON 245.415 45.605 245.520 45.510 245.415 45.510 ;
        POLYGON 245.960 45.605 246.035 45.605 246.035 45.540 ;
        RECT 246.035 45.575 247.175 45.605 ;
        POLYGON 247.175 45.635 247.270 45.575 247.175 45.575 ;
        POLYGON 252.430 45.635 252.430 45.615 252.395 45.615 ;
        RECT 252.430 45.615 253.670 45.635 ;
        POLYGON 252.395 45.615 252.395 45.605 252.380 45.605 ;
        RECT 252.395 45.605 253.670 45.615 ;
        POLYGON 252.375 45.605 252.375 45.575 252.325 45.575 ;
        RECT 252.375 45.575 253.670 45.605 ;
        RECT 246.035 45.540 247.270 45.575 ;
        POLYGON 246.035 45.540 246.070 45.540 246.070 45.510 ;
        RECT 246.070 45.535 247.270 45.540 ;
        POLYGON 247.270 45.575 247.345 45.535 247.270 45.535 ;
        POLYGON 252.325 45.575 252.325 45.555 252.295 45.555 ;
        RECT 252.325 45.555 253.670 45.575 ;
        POLYGON 252.290 45.555 252.290 45.535 252.255 45.535 ;
        RECT 252.290 45.535 253.670 45.555 ;
        RECT 246.070 45.525 247.345 45.535 ;
        POLYGON 247.345 45.535 247.360 45.525 247.345 45.525 ;
        POLYGON 252.255 45.535 252.255 45.525 252.240 45.525 ;
        RECT 252.255 45.525 253.670 45.535 ;
        RECT 246.070 45.510 247.360 45.525 ;
        RECT 244.755 45.480 245.520 45.510 ;
        POLYGON 245.520 45.510 245.550 45.480 245.520 45.480 ;
        POLYGON 246.070 45.510 246.105 45.510 246.105 45.480 ;
        RECT 246.105 45.495 247.360 45.510 ;
        POLYGON 247.360 45.525 247.415 45.495 247.360 45.495 ;
        POLYGON 252.240 45.525 252.240 45.515 252.220 45.515 ;
        RECT 252.240 45.520 253.670 45.525 ;
        POLYGON 253.670 45.640 253.805 45.640 253.670 45.520 ;
        POLYGON 254.360 45.640 254.360 45.585 254.305 45.585 ;
        RECT 254.360 45.585 254.940 45.640 ;
        POLYGON 254.305 45.585 254.305 45.520 254.235 45.520 ;
        RECT 254.305 45.580 254.940 45.585 ;
        POLYGON 254.940 45.735 255.070 45.735 254.940 45.580 ;
        POLYGON 255.810 45.735 255.810 45.730 255.805 45.730 ;
        RECT 255.810 45.730 256.570 45.735 ;
        POLYGON 255.805 45.725 255.805 45.675 255.765 45.675 ;
        RECT 255.805 45.695 256.570 45.730 ;
        POLYGON 256.570 45.950 256.715 45.950 256.570 45.695 ;
        POLYGON 257.565 45.945 257.565 45.880 257.530 45.880 ;
        RECT 257.565 45.880 258.580 45.950 ;
        POLYGON 258.580 46.175 258.705 46.175 258.580 45.880 ;
        POLYGON 260.045 46.175 260.045 45.975 259.980 45.975 ;
        RECT 260.045 45.975 261.580 46.185 ;
        POLYGON 259.980 45.975 259.980 45.905 259.955 45.905 ;
        RECT 259.980 45.935 261.580 45.975 ;
        POLYGON 261.580 46.190 261.665 46.190 261.580 45.935 ;
        POLYGON 263.735 46.190 263.735 46.145 263.725 46.145 ;
        RECT 263.735 46.145 266.475 46.195 ;
        POLYGON 263.725 46.145 263.725 45.935 263.675 45.935 ;
        RECT 263.725 45.935 266.475 46.145 ;
        RECT 259.980 45.905 261.485 45.935 ;
        POLYGON 259.955 45.905 259.955 45.880 259.945 45.880 ;
        RECT 259.955 45.880 261.485 45.905 ;
        POLYGON 257.530 45.880 257.530 45.760 257.465 45.760 ;
        RECT 257.530 45.810 258.545 45.880 ;
        POLYGON 258.545 45.880 258.580 45.880 258.545 45.810 ;
        POLYGON 259.945 45.875 259.945 45.810 259.920 45.810 ;
        RECT 259.945 45.810 261.485 45.880 ;
        RECT 257.530 45.760 258.445 45.810 ;
        POLYGON 257.465 45.760 257.465 45.700 257.435 45.700 ;
        RECT 257.465 45.700 258.445 45.760 ;
        RECT 255.805 45.675 256.525 45.695 ;
        POLYGON 255.765 45.675 255.765 45.580 255.700 45.580 ;
        RECT 255.765 45.630 256.525 45.675 ;
        POLYGON 256.525 45.695 256.570 45.695 256.525 45.630 ;
        POLYGON 257.435 45.695 257.435 45.680 257.425 45.680 ;
        RECT 257.435 45.680 258.445 45.700 ;
        POLYGON 257.425 45.680 257.425 45.655 257.410 45.655 ;
        RECT 257.425 45.655 258.445 45.680 ;
        POLYGON 257.410 45.655 257.410 45.635 257.400 45.635 ;
        RECT 257.410 45.635 258.445 45.655 ;
        RECT 255.765 45.610 256.515 45.630 ;
        POLYGON 256.515 45.630 256.525 45.630 256.515 45.610 ;
        POLYGON 257.400 45.630 257.400 45.615 257.390 45.615 ;
        RECT 257.400 45.615 258.445 45.635 ;
        POLYGON 257.390 45.615 257.390 45.610 257.385 45.610 ;
        RECT 257.390 45.610 258.445 45.615 ;
        RECT 255.765 45.580 256.410 45.610 ;
        RECT 254.305 45.570 254.935 45.580 ;
        POLYGON 254.935 45.580 254.940 45.580 254.935 45.570 ;
        POLYGON 255.700 45.580 255.700 45.570 255.690 45.570 ;
        RECT 255.700 45.570 256.410 45.580 ;
        RECT 254.305 45.520 254.850 45.570 ;
        RECT 252.240 45.515 253.660 45.520 ;
        POLYGON 252.220 45.515 252.220 45.505 252.205 45.505 ;
        RECT 252.220 45.510 253.660 45.515 ;
        POLYGON 253.660 45.520 253.670 45.520 253.660 45.510 ;
        POLYGON 254.235 45.520 254.235 45.510 254.225 45.510 ;
        RECT 254.235 45.510 254.850 45.520 ;
        RECT 252.220 45.505 253.640 45.510 ;
        POLYGON 252.205 45.505 252.205 45.495 252.185 45.495 ;
        RECT 252.205 45.495 253.640 45.505 ;
        POLYGON 253.640 45.510 253.660 45.510 253.640 45.495 ;
        POLYGON 254.225 45.510 254.225 45.495 254.205 45.495 ;
        RECT 254.225 45.495 254.850 45.510 ;
        RECT 246.105 45.485 247.415 45.495 ;
        POLYGON 247.415 45.495 247.430 45.485 247.415 45.485 ;
        POLYGON 252.185 45.495 252.185 45.485 252.165 45.485 ;
        RECT 252.185 45.485 253.535 45.495 ;
        RECT 246.105 45.480 247.430 45.485 ;
        RECT 240.755 45.450 241.990 45.480 ;
        POLYGON 241.990 45.480 242.010 45.450 241.990 45.450 ;
        POLYGON 243.060 45.480 243.080 45.480 243.080 45.450 ;
        RECT 243.080 45.460 243.975 45.480 ;
        POLYGON 243.975 45.480 243.985 45.460 243.975 45.460 ;
        POLYGON 244.755 45.480 244.775 45.480 244.775 45.460 ;
        RECT 244.775 45.460 245.550 45.480 ;
        RECT 243.080 45.450 243.985 45.460 ;
        POLYGON 243.985 45.460 244.000 45.450 243.985 45.450 ;
        POLYGON 244.775 45.460 244.785 45.460 244.785 45.450 ;
        RECT 244.785 45.450 245.550 45.460 ;
        RECT 237.085 45.385 239.125 45.395 ;
        POLYGON 239.125 45.395 239.130 45.385 239.125 45.385 ;
        RECT 240.755 45.385 242.010 45.450 ;
        RECT 237.085 45.350 239.130 45.385 ;
        POLYGON 239.130 45.385 239.145 45.350 239.130 45.350 ;
        POLYGON 240.755 45.385 240.775 45.385 240.775 45.355 ;
        RECT 240.775 45.350 242.010 45.385 ;
        RECT 237.085 45.315 239.145 45.350 ;
        POLYGON 237.085 45.315 237.245 45.315 237.245 44.965 ;
        RECT 237.245 45.225 239.145 45.315 ;
        POLYGON 239.145 45.350 239.205 45.225 239.145 45.225 ;
        POLYGON 240.775 45.350 240.830 45.350 240.830 45.260 ;
        RECT 240.830 45.310 242.010 45.350 ;
        POLYGON 242.010 45.450 242.105 45.310 242.010 45.310 ;
        POLYGON 243.080 45.450 243.110 45.450 243.110 45.410 ;
        RECT 243.110 45.430 244.000 45.450 ;
        POLYGON 244.000 45.450 244.015 45.430 244.000 45.430 ;
        POLYGON 244.785 45.450 244.800 45.450 244.800 45.430 ;
        RECT 244.800 45.430 245.550 45.450 ;
        RECT 243.110 45.410 244.015 45.430 ;
        POLYGON 243.110 45.410 243.190 45.410 243.190 45.310 ;
        RECT 243.190 45.325 244.015 45.410 ;
        POLYGON 244.015 45.430 244.100 45.325 244.015 45.325 ;
        POLYGON 244.800 45.430 244.905 45.430 244.905 45.325 ;
        RECT 244.905 45.420 245.550 45.430 ;
        POLYGON 245.550 45.480 245.615 45.420 245.550 45.420 ;
        POLYGON 246.105 45.480 246.130 45.480 246.130 45.460 ;
        RECT 246.130 45.460 247.430 45.480 ;
        POLYGON 246.130 45.460 246.175 45.460 246.175 45.425 ;
        RECT 246.175 45.425 247.430 45.460 ;
        POLYGON 246.175 45.425 246.180 45.425 246.180 45.420 ;
        RECT 246.180 45.420 247.430 45.425 ;
        POLYGON 247.430 45.485 247.550 45.420 247.430 45.420 ;
        POLYGON 252.165 45.485 252.165 45.465 252.125 45.465 ;
        RECT 252.165 45.465 253.535 45.485 ;
        POLYGON 252.125 45.465 252.125 45.450 252.100 45.450 ;
        RECT 252.125 45.450 253.535 45.465 ;
        POLYGON 252.100 45.450 252.100 45.420 252.040 45.420 ;
        RECT 252.100 45.420 253.535 45.450 ;
        RECT 244.905 45.330 245.615 45.420 ;
        POLYGON 245.615 45.420 245.710 45.330 245.615 45.330 ;
        POLYGON 246.180 45.420 246.260 45.420 246.260 45.365 ;
        RECT 246.260 45.400 247.550 45.420 ;
        POLYGON 247.550 45.420 247.590 45.400 247.550 45.400 ;
        POLYGON 252.040 45.420 252.040 45.400 252.000 45.400 ;
        RECT 252.040 45.405 253.535 45.420 ;
        POLYGON 253.535 45.495 253.640 45.495 253.535 45.405 ;
        POLYGON 254.205 45.495 254.205 45.475 254.185 45.475 ;
        RECT 254.205 45.480 254.850 45.495 ;
        POLYGON 254.850 45.570 254.935 45.570 254.850 45.480 ;
        POLYGON 255.690 45.570 255.690 45.545 255.675 45.545 ;
        RECT 255.690 45.545 256.410 45.570 ;
        POLYGON 255.675 45.545 255.675 45.520 255.655 45.520 ;
        RECT 255.675 45.520 256.410 45.545 ;
        POLYGON 255.655 45.520 255.655 45.480 255.625 45.480 ;
        RECT 255.655 45.480 256.410 45.520 ;
        RECT 254.205 45.475 254.730 45.480 ;
        POLYGON 254.185 45.475 254.185 45.430 254.135 45.430 ;
        RECT 254.185 45.430 254.730 45.475 ;
        POLYGON 254.135 45.430 254.135 45.405 254.105 45.405 ;
        RECT 254.135 45.405 254.730 45.430 ;
        RECT 252.040 45.400 253.410 45.405 ;
        RECT 246.260 45.390 247.590 45.400 ;
        POLYGON 247.590 45.400 247.615 45.390 247.590 45.390 ;
        POLYGON 252.000 45.400 252.000 45.390 251.980 45.390 ;
        RECT 252.000 45.390 253.410 45.400 ;
        RECT 246.260 45.365 247.615 45.390 ;
        POLYGON 246.260 45.365 246.300 45.365 246.300 45.330 ;
        RECT 246.300 45.355 247.615 45.365 ;
        POLYGON 247.615 45.390 247.690 45.355 247.615 45.355 ;
        POLYGON 251.980 45.390 251.980 45.375 251.950 45.375 ;
        RECT 251.980 45.375 253.410 45.390 ;
        POLYGON 251.950 45.375 251.950 45.360 251.915 45.360 ;
        RECT 251.950 45.360 253.410 45.375 ;
        POLYGON 251.915 45.360 251.915 45.355 251.905 45.355 ;
        RECT 251.915 45.355 253.410 45.360 ;
        RECT 246.300 45.330 247.690 45.355 ;
        RECT 244.905 45.325 245.715 45.330 ;
        RECT 243.190 45.310 244.100 45.325 ;
        RECT 240.830 45.260 242.105 45.310 ;
        POLYGON 240.830 45.260 240.850 45.260 240.850 45.225 ;
        RECT 240.850 45.225 242.105 45.260 ;
        RECT 237.245 44.970 239.205 45.225 ;
        POLYGON 239.205 45.225 239.340 44.970 239.205 44.970 ;
        POLYGON 240.850 45.225 240.915 45.225 240.915 45.120 ;
        RECT 240.915 45.220 242.105 45.225 ;
        POLYGON 242.105 45.310 242.165 45.220 242.105 45.220 ;
        POLYGON 243.190 45.310 243.235 45.310 243.235 45.255 ;
        RECT 243.235 45.295 244.100 45.310 ;
        POLYGON 244.100 45.325 244.130 45.295 244.100 45.295 ;
        POLYGON 244.905 45.325 244.935 45.325 244.935 45.295 ;
        RECT 244.935 45.295 245.715 45.325 ;
        RECT 243.235 45.255 244.130 45.295 ;
        POLYGON 243.235 45.255 243.245 45.255 243.245 45.235 ;
        RECT 243.245 45.235 244.130 45.255 ;
        POLYGON 243.245 45.235 243.255 45.235 243.255 45.220 ;
        RECT 243.255 45.225 244.130 45.235 ;
        POLYGON 244.130 45.295 244.185 45.225 244.130 45.225 ;
        POLYGON 244.935 45.295 245.005 45.295 245.005 45.225 ;
        RECT 245.005 45.240 245.715 45.295 ;
        POLYGON 245.715 45.330 245.820 45.240 245.715 45.240 ;
        POLYGON 246.300 45.330 246.355 45.330 246.355 45.290 ;
        RECT 246.355 45.325 247.690 45.330 ;
        POLYGON 247.690 45.355 247.750 45.325 247.690 45.325 ;
        POLYGON 251.905 45.355 251.905 45.325 251.850 45.325 ;
        RECT 251.905 45.325 253.410 45.355 ;
        RECT 246.355 45.290 247.750 45.325 ;
        POLYGON 246.355 45.290 246.405 45.290 246.405 45.255 ;
        RECT 246.405 45.265 247.750 45.290 ;
        POLYGON 247.750 45.325 247.890 45.265 247.750 45.265 ;
        POLYGON 251.850 45.325 251.850 45.310 251.805 45.310 ;
        RECT 251.850 45.310 253.410 45.325 ;
        POLYGON 251.805 45.310 251.805 45.295 251.775 45.295 ;
        RECT 251.805 45.305 253.410 45.310 ;
        POLYGON 253.410 45.405 253.535 45.405 253.410 45.305 ;
        POLYGON 254.105 45.405 254.105 45.365 254.065 45.365 ;
        RECT 254.105 45.365 254.730 45.405 ;
        POLYGON 254.065 45.365 254.065 45.305 253.990 45.305 ;
        RECT 254.065 45.350 254.730 45.365 ;
        POLYGON 254.730 45.480 254.850 45.480 254.730 45.350 ;
        POLYGON 255.625 45.480 255.625 45.365 255.535 45.365 ;
        RECT 255.625 45.445 256.410 45.480 ;
        POLYGON 256.410 45.610 256.515 45.610 256.410 45.445 ;
        POLYGON 257.385 45.605 257.385 45.465 257.305 45.465 ;
        RECT 257.385 45.590 258.445 45.610 ;
        POLYGON 258.445 45.810 258.545 45.810 258.445 45.590 ;
        POLYGON 259.920 45.805 259.920 45.745 259.900 45.745 ;
        RECT 259.920 45.745 261.485 45.810 ;
        POLYGON 259.900 45.745 259.900 45.685 259.875 45.685 ;
        RECT 259.900 45.685 261.485 45.745 ;
        POLYGON 259.875 45.685 259.875 45.595 259.835 45.595 ;
        RECT 259.875 45.665 261.485 45.685 ;
        POLYGON 261.485 45.935 261.580 45.935 261.485 45.665 ;
        POLYGON 263.675 45.935 263.675 45.890 263.665 45.890 ;
        RECT 263.675 45.890 266.475 45.935 ;
        POLYGON 263.665 45.890 263.665 45.675 263.615 45.675 ;
        RECT 263.665 45.850 266.475 45.890 ;
        POLYGON 266.475 46.405 266.565 46.405 266.475 45.850 ;
        POLYGON 270.680 46.405 270.680 45.850 270.675 45.850 ;
        RECT 270.680 46.395 277.905 46.445 ;
        POLYGON 277.905 46.780 277.915 46.780 277.905 46.405 ;
        POLYGON 287.925 46.935 287.925 46.445 287.900 46.445 ;
        RECT 287.925 46.445 303.120 46.970 ;
        RECT 270.680 45.850 277.885 46.395 ;
        RECT 263.665 45.820 266.470 45.850 ;
        POLYGON 266.470 45.850 266.475 45.850 266.470 45.820 ;
        RECT 263.665 45.675 266.365 45.820 ;
        RECT 259.875 45.595 261.250 45.665 ;
        RECT 257.385 45.520 258.410 45.590 ;
        POLYGON 258.410 45.590 258.445 45.590 258.410 45.520 ;
        POLYGON 259.835 45.590 259.835 45.560 259.820 45.560 ;
        RECT 259.835 45.560 261.250 45.595 ;
        POLYGON 259.820 45.560 259.820 45.520 259.805 45.520 ;
        RECT 259.820 45.520 261.250 45.560 ;
        RECT 257.385 45.465 258.295 45.520 ;
        POLYGON 257.305 45.465 257.305 45.450 257.295 45.450 ;
        RECT 257.305 45.450 258.295 45.465 ;
        RECT 255.625 45.365 256.275 45.445 ;
        POLYGON 255.535 45.365 255.535 45.355 255.525 45.355 ;
        RECT 255.535 45.355 256.275 45.365 ;
        RECT 254.065 45.305 254.615 45.350 ;
        RECT 251.805 45.295 253.390 45.305 ;
        POLYGON 251.775 45.295 251.775 45.290 251.760 45.290 ;
        RECT 251.775 45.290 253.390 45.295 ;
        POLYGON 253.390 45.305 253.405 45.305 253.390 45.290 ;
        POLYGON 253.990 45.305 253.990 45.290 253.975 45.290 ;
        RECT 253.990 45.290 254.615 45.305 ;
        POLYGON 251.760 45.290 251.760 45.265 251.705 45.265 ;
        RECT 251.760 45.265 253.250 45.290 ;
        RECT 246.405 45.255 247.895 45.265 ;
        POLYGON 246.405 45.255 246.425 45.255 246.425 45.240 ;
        RECT 246.425 45.250 247.895 45.255 ;
        POLYGON 247.895 45.265 247.915 45.250 247.895 45.250 ;
        POLYGON 251.705 45.265 251.705 45.250 251.670 45.250 ;
        RECT 251.705 45.250 253.250 45.265 ;
        RECT 246.425 45.245 247.915 45.250 ;
        POLYGON 247.915 45.250 247.935 45.245 247.915 45.245 ;
        POLYGON 251.670 45.250 251.670 45.245 251.660 45.245 ;
        RECT 251.670 45.245 253.250 45.250 ;
        RECT 246.425 45.240 247.935 45.245 ;
        RECT 245.005 45.225 245.820 45.240 ;
        RECT 243.255 45.220 244.185 45.225 ;
        RECT 240.915 45.195 242.165 45.220 ;
        POLYGON 242.165 45.220 242.185 45.195 242.165 45.195 ;
        RECT 240.915 45.130 242.185 45.195 ;
        POLYGON 243.255 45.220 243.280 45.220 243.280 45.190 ;
        RECT 243.280 45.190 244.185 45.220 ;
        POLYGON 242.185 45.190 242.235 45.130 242.185 45.130 ;
        POLYGON 243.280 45.190 243.325 45.190 243.325 45.130 ;
        RECT 243.325 45.170 244.185 45.190 ;
        POLYGON 244.185 45.225 244.240 45.170 244.185 45.170 ;
        POLYGON 245.005 45.225 245.040 45.225 245.040 45.195 ;
        RECT 245.040 45.195 245.820 45.225 ;
        POLYGON 245.040 45.195 245.065 45.195 245.065 45.170 ;
        RECT 245.065 45.170 245.820 45.195 ;
        RECT 243.325 45.140 244.240 45.170 ;
        POLYGON 244.240 45.170 244.265 45.140 244.240 45.140 ;
        POLYGON 245.065 45.170 245.095 45.170 245.095 45.140 ;
        RECT 245.095 45.160 245.820 45.170 ;
        POLYGON 245.820 45.240 245.915 45.160 245.820 45.160 ;
        POLYGON 246.425 45.240 246.490 45.240 246.490 45.200 ;
        RECT 246.490 45.230 247.935 45.240 ;
        POLYGON 247.935 45.245 247.975 45.230 247.935 45.230 ;
        POLYGON 251.660 45.245 251.660 45.230 251.620 45.230 ;
        RECT 251.660 45.230 253.250 45.245 ;
        RECT 246.490 45.200 247.975 45.230 ;
        POLYGON 246.490 45.200 246.545 45.200 246.545 45.160 ;
        RECT 246.545 45.185 247.975 45.200 ;
        POLYGON 247.975 45.230 248.085 45.185 247.975 45.185 ;
        POLYGON 251.620 45.230 251.620 45.225 251.605 45.225 ;
        RECT 251.620 45.225 253.250 45.230 ;
        POLYGON 251.605 45.225 251.605 45.220 251.595 45.220 ;
        RECT 251.605 45.220 253.250 45.225 ;
        POLYGON 251.595 45.220 251.595 45.190 251.515 45.190 ;
        RECT 251.595 45.190 253.250 45.220 ;
        POLYGON 253.250 45.290 253.390 45.290 253.250 45.190 ;
        POLYGON 253.975 45.290 253.975 45.275 253.955 45.275 ;
        RECT 253.975 45.275 254.615 45.290 ;
        POLYGON 253.955 45.275 253.955 45.255 253.935 45.255 ;
        RECT 253.955 45.255 254.615 45.275 ;
        POLYGON 253.935 45.255 253.935 45.245 253.920 45.245 ;
        RECT 253.935 45.245 254.615 45.255 ;
        POLYGON 253.920 45.245 253.920 45.205 253.870 45.205 ;
        RECT 253.920 45.235 254.615 45.245 ;
        POLYGON 254.615 45.350 254.730 45.350 254.615 45.235 ;
        POLYGON 255.525 45.350 255.525 45.315 255.495 45.315 ;
        RECT 255.525 45.315 256.275 45.355 ;
        POLYGON 255.495 45.310 255.495 45.295 255.480 45.295 ;
        RECT 255.495 45.295 256.275 45.315 ;
        POLYGON 255.480 45.295 255.480 45.235 255.430 45.235 ;
        RECT 255.480 45.245 256.275 45.295 ;
        POLYGON 256.275 45.445 256.410 45.445 256.275 45.245 ;
        POLYGON 257.295 45.445 257.295 45.330 257.225 45.330 ;
        RECT 257.295 45.330 258.295 45.450 ;
        POLYGON 257.225 45.330 257.225 45.320 257.215 45.320 ;
        RECT 257.225 45.320 258.295 45.330 ;
        POLYGON 257.215 45.320 257.215 45.300 257.205 45.300 ;
        RECT 257.215 45.300 258.295 45.320 ;
        POLYGON 258.295 45.520 258.410 45.520 258.295 45.300 ;
        POLYGON 259.805 45.520 259.805 45.470 259.785 45.470 ;
        RECT 259.805 45.470 261.250 45.520 ;
        POLYGON 259.785 45.470 259.785 45.300 259.715 45.300 ;
        RECT 259.785 45.300 261.250 45.470 ;
        POLYGON 257.205 45.300 257.205 45.295 257.200 45.295 ;
        RECT 257.205 45.295 258.245 45.300 ;
        POLYGON 257.200 45.295 257.200 45.245 257.170 45.245 ;
        RECT 257.200 45.245 258.245 45.295 ;
        RECT 255.480 45.235 256.265 45.245 ;
        POLYGON 256.265 45.245 256.275 45.245 256.265 45.235 ;
        POLYGON 257.170 45.245 257.170 45.235 257.165 45.235 ;
        RECT 257.170 45.235 258.245 45.245 ;
        RECT 253.920 45.205 254.525 45.235 ;
        POLYGON 253.870 45.205 253.870 45.190 253.850 45.190 ;
        RECT 253.870 45.190 254.525 45.205 ;
        POLYGON 251.515 45.190 251.515 45.185 251.505 45.185 ;
        RECT 251.515 45.185 253.245 45.190 ;
        POLYGON 253.245 45.190 253.250 45.190 253.245 45.185 ;
        POLYGON 253.850 45.190 253.850 45.185 253.845 45.185 ;
        RECT 253.850 45.185 254.525 45.190 ;
        RECT 246.545 45.170 248.085 45.185 ;
        POLYGON 248.085 45.185 248.135 45.170 248.085 45.170 ;
        POLYGON 251.505 45.185 251.505 45.180 251.490 45.180 ;
        RECT 251.505 45.180 253.170 45.185 ;
        POLYGON 251.490 45.180 251.490 45.170 251.465 45.170 ;
        RECT 251.490 45.170 253.170 45.180 ;
        RECT 246.545 45.160 248.135 45.170 ;
        RECT 245.095 45.140 245.915 45.160 ;
        RECT 243.325 45.130 244.265 45.140 ;
        RECT 240.915 45.120 242.235 45.130 ;
        POLYGON 240.915 45.120 241.000 45.120 241.000 44.970 ;
        RECT 241.000 44.970 242.235 45.120 ;
        RECT 237.245 44.965 239.340 44.970 ;
        RECT 230.285 44.935 234.380 44.965 ;
        POLYGON 234.380 44.965 234.390 44.935 234.380 44.935 ;
        POLYGON 237.245 44.965 237.255 44.965 237.255 44.940 ;
        RECT 237.255 44.935 239.340 44.965 ;
        RECT 230.285 44.830 234.390 44.935 ;
        POLYGON 234.390 44.935 234.430 44.830 234.390 44.830 ;
        POLYGON 237.255 44.935 237.305 44.935 237.305 44.835 ;
        RECT 237.305 44.830 239.340 44.935 ;
        RECT 230.285 44.760 234.430 44.830 ;
        POLYGON 230.285 44.760 230.290 44.760 230.290 44.740 ;
        RECT 230.290 44.740 234.430 44.760 ;
        RECT 182.900 44.210 198.000 44.610 ;
        POLYGON 182.810 44.210 182.810 44.075 182.795 44.075 ;
        RECT 182.810 44.095 198.000 44.210 ;
        POLYGON 198.000 44.610 198.035 44.095 198.000 44.095 ;
        RECT 208.330 44.605 223.235 44.740 ;
        POLYGON 223.235 44.740 223.280 44.605 223.235 44.605 ;
        POLYGON 230.290 44.740 230.320 44.740 230.320 44.645 ;
        RECT 230.320 44.645 234.430 44.740 ;
        RECT 208.330 44.600 223.280 44.605 ;
        POLYGON 230.320 44.645 230.335 44.645 230.335 44.600 ;
        RECT 230.335 44.605 234.430 44.645 ;
        POLYGON 234.430 44.830 234.525 44.605 234.430 44.605 ;
        POLYGON 237.305 44.830 237.335 44.830 237.335 44.770 ;
        RECT 237.335 44.770 239.340 44.830 ;
        POLYGON 237.335 44.770 237.410 44.770 237.410 44.605 ;
        RECT 237.410 44.760 239.340 44.770 ;
        POLYGON 239.340 44.970 239.450 44.760 239.340 44.760 ;
        POLYGON 241.000 44.970 241.005 44.970 241.005 44.965 ;
        RECT 241.005 44.965 242.235 44.970 ;
        POLYGON 241.005 44.965 241.090 44.965 241.090 44.835 ;
        RECT 241.090 44.940 242.235 44.965 ;
        POLYGON 242.235 45.130 242.370 44.940 242.235 44.940 ;
        POLYGON 243.325 45.130 243.395 45.130 243.395 45.045 ;
        RECT 243.395 45.050 244.265 45.130 ;
        POLYGON 244.265 45.140 244.350 45.050 244.265 45.050 ;
        POLYGON 245.095 45.140 245.200 45.140 245.200 45.050 ;
        RECT 245.200 45.125 245.915 45.140 ;
        POLYGON 245.915 45.160 245.955 45.125 245.915 45.125 ;
        POLYGON 246.545 45.160 246.590 45.160 246.590 45.130 ;
        RECT 246.590 45.155 248.135 45.160 ;
        POLYGON 248.135 45.170 248.180 45.155 248.135 45.155 ;
        POLYGON 251.465 45.170 251.465 45.165 251.450 45.165 ;
        RECT 251.465 45.165 253.170 45.170 ;
        POLYGON 251.450 45.165 251.450 45.155 251.425 45.155 ;
        RECT 251.450 45.155 253.170 45.165 ;
        RECT 246.590 45.130 248.180 45.155 ;
        POLYGON 248.180 45.155 248.250 45.130 248.180 45.130 ;
        POLYGON 251.425 45.155 251.425 45.150 251.410 45.150 ;
        RECT 251.425 45.150 253.170 45.155 ;
        POLYGON 251.410 45.150 251.410 45.140 251.375 45.140 ;
        RECT 251.410 45.140 253.170 45.150 ;
        POLYGON 246.590 45.130 246.595 45.130 246.595 45.125 ;
        RECT 246.595 45.125 248.250 45.130 ;
        POLYGON 251.375 45.140 251.375 45.125 251.335 45.125 ;
        RECT 251.375 45.135 253.170 45.140 ;
        POLYGON 253.170 45.185 253.245 45.185 253.170 45.135 ;
        POLYGON 253.845 45.185 253.845 45.155 253.805 45.155 ;
        RECT 253.845 45.155 254.525 45.185 ;
        POLYGON 253.805 45.155 253.805 45.135 253.780 45.135 ;
        RECT 253.805 45.140 254.525 45.155 ;
        POLYGON 254.525 45.235 254.615 45.235 254.525 45.140 ;
        POLYGON 255.430 45.235 255.430 45.185 255.390 45.185 ;
        RECT 255.430 45.205 256.245 45.235 ;
        POLYGON 256.245 45.235 256.265 45.235 256.245 45.205 ;
        POLYGON 257.165 45.235 257.165 45.205 257.145 45.205 ;
        RECT 257.165 45.210 258.245 45.235 ;
        POLYGON 258.245 45.300 258.295 45.300 258.245 45.210 ;
        POLYGON 259.715 45.300 259.715 45.275 259.705 45.275 ;
        RECT 259.715 45.275 261.250 45.300 ;
        POLYGON 259.705 45.275 259.705 45.245 259.695 45.245 ;
        RECT 259.705 45.245 261.250 45.275 ;
        POLYGON 259.695 45.245 259.695 45.210 259.680 45.210 ;
        RECT 259.695 45.210 261.250 45.245 ;
        RECT 257.165 45.205 258.140 45.210 ;
        RECT 255.430 45.185 256.070 45.205 ;
        POLYGON 255.390 45.185 255.390 45.140 255.350 45.140 ;
        RECT 255.390 45.140 256.070 45.185 ;
        RECT 253.805 45.135 254.475 45.140 ;
        RECT 251.375 45.125 253.115 45.135 ;
        RECT 245.200 45.060 245.955 45.125 ;
        POLYGON 245.955 45.125 246.035 45.060 245.955 45.060 ;
        POLYGON 246.595 45.125 246.640 45.125 246.640 45.100 ;
        RECT 246.640 45.100 248.265 45.125 ;
        POLYGON 248.265 45.125 248.335 45.100 248.265 45.100 ;
        POLYGON 251.335 45.125 251.335 45.115 251.310 45.115 ;
        RECT 251.335 45.115 253.115 45.125 ;
        POLYGON 251.295 45.115 251.295 45.100 251.250 45.100 ;
        RECT 251.295 45.100 253.115 45.115 ;
        POLYGON 246.645 45.100 246.705 45.100 246.705 45.060 ;
        RECT 246.705 45.075 248.340 45.100 ;
        POLYGON 248.340 45.100 248.425 45.075 248.340 45.075 ;
        POLYGON 251.250 45.100 251.250 45.095 251.235 45.095 ;
        RECT 251.250 45.095 253.115 45.100 ;
        POLYGON 253.115 45.135 253.170 45.135 253.115 45.095 ;
        POLYGON 253.780 45.135 253.780 45.095 253.730 45.095 ;
        RECT 253.780 45.095 254.475 45.135 ;
        POLYGON 251.235 45.095 251.235 45.090 251.225 45.090 ;
        RECT 251.235 45.090 253.095 45.095 ;
        POLYGON 251.225 45.090 251.225 45.075 251.175 45.075 ;
        RECT 251.225 45.080 253.095 45.090 ;
        POLYGON 253.095 45.095 253.115 45.095 253.095 45.080 ;
        POLYGON 253.730 45.095 253.730 45.080 253.715 45.080 ;
        RECT 253.730 45.090 254.475 45.095 ;
        POLYGON 254.475 45.140 254.525 45.140 254.475 45.090 ;
        POLYGON 255.350 45.140 255.350 45.105 255.320 45.105 ;
        RECT 255.350 45.105 256.070 45.140 ;
        POLYGON 255.320 45.105 255.320 45.090 255.310 45.090 ;
        RECT 255.320 45.090 256.070 45.105 ;
        RECT 253.730 45.080 254.380 45.090 ;
        RECT 251.225 45.075 252.975 45.080 ;
        RECT 246.705 45.060 248.425 45.075 ;
        POLYGON 248.425 45.075 248.470 45.060 248.425 45.060 ;
        POLYGON 251.175 45.075 251.175 45.065 251.140 45.065 ;
        RECT 251.175 45.065 252.975 45.075 ;
        POLYGON 251.140 45.065 251.140 45.060 251.130 45.060 ;
        RECT 251.140 45.060 252.975 45.065 ;
        RECT 245.200 45.050 246.035 45.060 ;
        RECT 243.395 45.045 244.350 45.050 ;
        POLYGON 243.395 45.045 243.435 45.045 243.435 45.000 ;
        RECT 243.435 45.015 244.350 45.045 ;
        POLYGON 244.350 45.050 244.385 45.015 244.350 45.015 ;
        POLYGON 245.200 45.050 245.225 45.050 245.225 45.030 ;
        RECT 245.225 45.030 246.035 45.050 ;
        POLYGON 245.225 45.030 245.240 45.030 245.240 45.015 ;
        RECT 245.240 45.015 246.035 45.030 ;
        POLYGON 246.035 45.060 246.085 45.015 246.035 45.015 ;
        POLYGON 246.705 45.060 246.725 45.060 246.725 45.050 ;
        RECT 246.725 45.050 248.475 45.060 ;
        POLYGON 246.725 45.050 246.780 45.050 246.780 45.015 ;
        RECT 246.780 45.040 248.475 45.050 ;
        POLYGON 248.475 45.060 248.545 45.040 248.475 45.040 ;
        POLYGON 251.130 45.060 251.130 45.055 251.095 45.055 ;
        RECT 251.130 45.055 252.975 45.060 ;
        POLYGON 251.095 45.055 251.095 45.040 251.035 45.040 ;
        RECT 251.095 45.040 252.975 45.055 ;
        RECT 246.780 45.035 248.545 45.040 ;
        POLYGON 248.545 45.040 248.565 45.035 248.545 45.035 ;
        POLYGON 251.035 45.040 251.035 45.035 251.015 45.035 ;
        RECT 251.035 45.035 252.975 45.040 ;
        RECT 246.780 45.030 248.565 45.035 ;
        POLYGON 248.565 45.035 248.595 45.030 248.565 45.030 ;
        RECT 246.780 45.015 248.595 45.030 ;
        POLYGON 251.015 45.035 251.015 45.025 250.980 45.025 ;
        RECT 251.015 45.025 252.975 45.035 ;
        RECT 243.435 45.000 244.385 45.015 ;
        POLYGON 243.435 45.000 243.485 45.000 243.485 44.940 ;
        RECT 243.485 44.995 244.385 45.000 ;
        POLYGON 244.385 45.015 244.400 44.995 244.385 44.995 ;
        POLYGON 245.240 45.015 245.260 45.015 245.260 44.995 ;
        RECT 245.260 44.995 246.085 45.015 ;
        RECT 243.485 44.940 244.400 44.995 ;
        RECT 241.090 44.925 242.370 44.940 ;
        POLYGON 242.370 44.940 242.385 44.925 242.370 44.925 ;
        POLYGON 243.485 44.940 243.500 44.940 243.500 44.925 ;
        RECT 243.500 44.925 244.400 44.940 ;
        RECT 241.090 44.875 242.385 44.925 ;
        POLYGON 242.385 44.925 242.420 44.875 242.385 44.875 ;
        POLYGON 243.500 44.925 243.545 44.925 243.545 44.875 ;
        RECT 243.545 44.875 244.400 44.925 ;
        RECT 241.090 44.835 242.420 44.875 ;
        POLYGON 241.090 44.835 241.135 44.835 241.135 44.765 ;
        RECT 241.135 44.760 242.420 44.835 ;
        RECT 237.410 44.605 239.450 44.760 ;
        POLYGON 239.450 44.760 239.545 44.605 239.450 44.605 ;
        RECT 230.335 44.600 234.525 44.605 ;
        RECT 237.410 44.600 239.545 44.605 ;
        POLYGON 241.135 44.760 241.240 44.760 241.240 44.600 ;
        RECT 241.240 44.745 242.420 44.760 ;
        POLYGON 242.420 44.875 242.525 44.745 242.420 44.745 ;
        POLYGON 243.545 44.875 243.630 44.875 243.630 44.780 ;
        RECT 243.630 44.860 244.400 44.875 ;
        POLYGON 244.400 44.995 244.535 44.860 244.400 44.860 ;
        POLYGON 245.260 44.995 245.415 44.995 245.415 44.865 ;
        RECT 245.415 44.985 246.085 44.995 ;
        POLYGON 246.085 45.015 246.130 44.985 246.085 44.985 ;
        POLYGON 246.780 45.015 246.830 45.015 246.830 44.985 ;
        RECT 246.830 44.990 248.595 45.015 ;
        POLYGON 248.595 45.025 248.750 44.990 248.595 44.990 ;
        POLYGON 250.980 45.025 250.980 45.020 250.960 45.020 ;
        RECT 250.980 45.020 252.975 45.025 ;
        POLYGON 250.960 45.020 250.960 45.015 250.945 45.015 ;
        RECT 250.960 45.015 252.975 45.020 ;
        POLYGON 250.945 45.015 250.945 44.990 250.845 44.990 ;
        RECT 250.945 45.005 252.975 45.015 ;
        POLYGON 252.975 45.080 253.095 45.080 252.975 45.005 ;
        POLYGON 253.715 45.080 253.715 45.045 253.670 45.045 ;
        RECT 253.715 45.045 254.380 45.080 ;
        POLYGON 253.670 45.045 253.670 45.035 253.660 45.035 ;
        RECT 253.670 45.035 254.380 45.045 ;
        POLYGON 253.655 45.035 253.655 45.025 253.640 45.025 ;
        RECT 253.655 45.025 254.380 45.035 ;
        POLYGON 253.640 45.025 253.640 45.005 253.615 45.005 ;
        RECT 253.640 45.005 254.380 45.025 ;
        POLYGON 254.380 45.090 254.475 45.090 254.380 45.005 ;
        POLYGON 255.310 45.090 255.310 45.065 255.290 45.065 ;
        RECT 255.310 45.065 256.070 45.090 ;
        POLYGON 255.290 45.065 255.290 45.005 255.230 45.005 ;
        RECT 255.290 45.005 256.070 45.065 ;
        RECT 250.945 44.990 252.940 45.005 ;
        RECT 246.830 44.985 248.750 44.990 ;
        POLYGON 248.750 44.990 248.770 44.985 248.750 44.985 ;
        POLYGON 250.830 44.990 250.830 44.985 250.810 44.985 ;
        RECT 250.830 44.985 252.940 44.990 ;
        POLYGON 252.940 45.005 252.975 45.005 252.940 44.985 ;
        POLYGON 253.615 45.005 253.615 44.985 253.590 44.985 ;
        RECT 253.615 44.985 254.310 45.005 ;
        RECT 245.415 44.950 246.130 44.985 ;
        POLYGON 246.130 44.985 246.175 44.950 246.130 44.950 ;
        POLYGON 246.830 44.985 246.890 44.985 246.890 44.950 ;
        RECT 246.890 44.965 248.775 44.985 ;
        POLYGON 248.775 44.985 248.870 44.965 248.775 44.965 ;
        POLYGON 250.810 44.985 250.810 44.975 250.765 44.975 ;
        RECT 250.810 44.980 252.930 44.985 ;
        POLYGON 252.930 44.985 252.940 44.985 252.930 44.980 ;
        POLYGON 253.590 44.985 253.590 44.980 253.585 44.980 ;
        RECT 253.590 44.980 254.310 44.985 ;
        RECT 250.810 44.975 252.830 44.980 ;
        POLYGON 250.765 44.975 250.765 44.965 250.705 44.965 ;
        RECT 250.765 44.965 252.830 44.975 ;
        RECT 246.890 44.955 248.875 44.965 ;
        POLYGON 248.875 44.965 248.945 44.955 248.875 44.955 ;
        POLYGON 250.700 44.965 250.700 44.955 250.660 44.955 ;
        RECT 250.700 44.955 252.830 44.965 ;
        RECT 246.890 44.950 248.950 44.955 ;
        POLYGON 250.650 44.955 250.650 44.950 250.630 44.950 ;
        RECT 250.650 44.950 252.830 44.955 ;
        RECT 245.415 44.890 246.175 44.950 ;
        POLYGON 246.175 44.950 246.260 44.890 246.175 44.890 ;
        POLYGON 246.890 44.950 247.000 44.950 247.000 44.890 ;
        RECT 247.000 44.930 248.950 44.950 ;
        POLYGON 248.950 44.950 249.075 44.930 248.950 44.930 ;
        POLYGON 250.630 44.950 250.630 44.940 250.585 44.940 ;
        RECT 250.630 44.940 252.830 44.950 ;
        POLYGON 250.580 44.940 250.580 44.930 250.515 44.930 ;
        RECT 250.580 44.930 252.830 44.940 ;
        RECT 247.000 44.925 249.085 44.930 ;
        POLYGON 249.085 44.930 249.125 44.925 249.085 44.925 ;
        POLYGON 250.515 44.930 250.515 44.925 250.480 44.925 ;
        RECT 250.515 44.925 252.830 44.930 ;
        RECT 247.000 44.920 249.125 44.925 ;
        POLYGON 249.125 44.925 249.145 44.920 249.125 44.920 ;
        POLYGON 250.455 44.925 250.455 44.920 250.425 44.920 ;
        RECT 250.455 44.920 252.830 44.925 ;
        POLYGON 252.830 44.980 252.930 44.980 252.830 44.920 ;
        POLYGON 253.585 44.980 253.585 44.940 253.535 44.940 ;
        RECT 253.585 44.940 254.310 44.980 ;
        POLYGON 254.310 45.005 254.380 45.005 254.310 44.940 ;
        POLYGON 255.230 45.005 255.230 44.940 255.175 44.940 ;
        RECT 255.230 44.970 256.070 45.005 ;
        POLYGON 256.070 45.205 256.245 45.205 256.070 44.970 ;
        POLYGON 257.145 45.205 257.145 45.130 257.100 45.130 ;
        RECT 257.145 45.130 258.140 45.205 ;
        POLYGON 257.100 45.130 257.100 45.020 257.030 45.020 ;
        RECT 257.100 45.020 258.140 45.130 ;
        POLYGON 257.030 45.020 257.030 44.975 256.995 44.975 ;
        RECT 257.030 45.015 258.140 45.020 ;
        POLYGON 258.140 45.210 258.245 45.210 258.140 45.015 ;
        POLYGON 259.680 45.210 259.680 45.080 259.620 45.080 ;
        RECT 259.680 45.095 261.250 45.210 ;
        POLYGON 261.250 45.665 261.485 45.665 261.250 45.095 ;
        POLYGON 263.615 45.665 263.615 45.610 263.600 45.610 ;
        RECT 263.615 45.610 266.365 45.675 ;
        POLYGON 263.600 45.600 263.600 45.365 263.535 45.365 ;
        RECT 263.600 45.365 266.365 45.610 ;
        POLYGON 263.535 45.365 263.535 45.225 263.495 45.225 ;
        RECT 263.535 45.255 266.365 45.365 ;
        POLYGON 266.365 45.820 266.470 45.820 266.365 45.255 ;
        POLYGON 270.675 45.770 270.675 45.545 270.660 45.545 ;
        RECT 270.675 45.630 277.885 45.850 ;
        POLYGON 277.885 46.395 277.905 46.395 277.885 45.630 ;
        POLYGON 287.900 46.405 287.900 45.650 287.860 45.650 ;
        RECT 287.900 45.650 303.120 46.445 ;
        RECT 270.675 45.545 277.820 45.630 ;
        POLYGON 270.660 45.545 270.660 45.295 270.645 45.295 ;
        RECT 270.660 45.295 277.820 45.545 ;
        RECT 263.535 45.225 266.230 45.255 ;
        POLYGON 263.495 45.225 263.495 45.100 263.465 45.100 ;
        RECT 263.495 45.100 266.230 45.225 ;
        RECT 259.680 45.080 261.085 45.095 ;
        POLYGON 259.620 45.080 259.620 45.035 259.595 45.035 ;
        RECT 259.620 45.035 261.085 45.080 ;
        POLYGON 259.595 45.035 259.595 45.015 259.585 45.015 ;
        RECT 259.595 45.015 261.085 45.035 ;
        RECT 257.030 44.975 258.010 45.015 ;
        RECT 255.230 44.940 256.015 44.970 ;
        POLYGON 253.535 44.940 253.535 44.920 253.505 44.920 ;
        RECT 253.535 44.920 254.235 44.940 ;
        RECT 247.000 44.915 249.150 44.920 ;
        POLYGON 249.150 44.920 249.185 44.915 249.150 44.915 ;
        POLYGON 250.425 44.920 250.425 44.915 250.395 44.915 ;
        RECT 250.425 44.915 252.785 44.920 ;
        RECT 247.000 44.905 249.190 44.915 ;
        POLYGON 249.190 44.915 249.300 44.905 249.190 44.905 ;
        POLYGON 250.395 44.915 250.395 44.910 250.380 44.910 ;
        RECT 250.395 44.910 252.785 44.915 ;
        POLYGON 250.375 44.910 250.375 44.905 250.290 44.905 ;
        RECT 250.375 44.905 252.785 44.910 ;
        RECT 247.000 44.895 249.305 44.905 ;
        RECT 250.285 44.900 252.785 44.905 ;
        POLYGON 249.305 44.900 249.390 44.895 249.305 44.895 ;
        POLYGON 250.255 44.900 250.255 44.895 250.215 44.895 ;
        RECT 250.255 44.895 252.785 44.900 ;
        RECT 247.000 44.890 249.400 44.895 ;
        RECT 245.415 44.865 246.260 44.890 ;
        POLYGON 245.415 44.865 245.420 44.865 245.420 44.860 ;
        RECT 245.420 44.860 246.260 44.865 ;
        RECT 243.630 44.835 244.535 44.860 ;
        POLYGON 244.535 44.860 244.565 44.835 244.535 44.835 ;
        POLYGON 245.420 44.860 245.440 44.860 245.440 44.845 ;
        RECT 245.440 44.845 246.260 44.860 ;
        POLYGON 245.440 44.845 245.450 44.845 245.450 44.835 ;
        RECT 245.450 44.835 246.260 44.845 ;
        RECT 243.630 44.780 244.565 44.835 ;
        POLYGON 243.630 44.780 243.650 44.780 243.650 44.755 ;
        RECT 243.650 44.770 244.565 44.780 ;
        POLYGON 244.565 44.835 244.625 44.770 244.565 44.770 ;
        POLYGON 245.450 44.835 245.535 44.835 245.535 44.770 ;
        RECT 245.535 44.820 246.260 44.835 ;
        POLYGON 246.260 44.890 246.355 44.820 246.260 44.820 ;
        POLYGON 247.000 44.890 247.085 44.890 247.085 44.845 ;
        RECT 247.085 44.885 249.400 44.890 ;
        POLYGON 249.400 44.895 249.485 44.885 249.400 44.885 ;
        POLYGON 250.205 44.895 250.205 44.890 250.140 44.890 ;
        RECT 250.205 44.890 252.785 44.895 ;
        POLYGON 252.785 44.920 252.830 44.920 252.785 44.890 ;
        POLYGON 253.505 44.920 253.505 44.890 253.460 44.890 ;
        RECT 253.505 44.890 254.235 44.920 ;
        POLYGON 250.135 44.890 250.135 44.885 250.080 44.885 ;
        RECT 250.135 44.885 252.690 44.890 ;
        RECT 247.085 44.880 249.540 44.885 ;
        POLYGON 249.540 44.885 249.665 44.880 249.540 44.880 ;
        POLYGON 250.020 44.885 250.020 44.880 249.995 44.880 ;
        RECT 250.020 44.880 252.690 44.885 ;
        RECT 247.085 44.845 252.690 44.880 ;
        POLYGON 247.085 44.845 247.135 44.845 247.135 44.820 ;
        RECT 247.135 44.840 252.690 44.845 ;
        POLYGON 252.690 44.890 252.785 44.890 252.690 44.840 ;
        POLYGON 253.460 44.890 253.460 44.855 253.410 44.855 ;
        RECT 253.460 44.875 254.235 44.890 ;
        POLYGON 254.235 44.940 254.310 44.940 254.235 44.875 ;
        POLYGON 255.175 44.940 255.175 44.895 255.135 44.895 ;
        RECT 255.175 44.895 256.015 44.940 ;
        POLYGON 256.015 44.970 256.070 44.970 256.015 44.895 ;
        POLYGON 256.995 44.970 256.995 44.955 256.985 44.955 ;
        RECT 256.995 44.955 258.010 44.975 ;
        POLYGON 256.985 44.955 256.985 44.950 256.980 44.950 ;
        RECT 256.985 44.950 258.010 44.955 ;
        POLYGON 256.980 44.950 256.980 44.900 256.945 44.900 ;
        RECT 256.980 44.900 258.010 44.950 ;
        POLYGON 255.135 44.895 255.135 44.875 255.115 44.875 ;
        RECT 255.135 44.885 256.005 44.895 ;
        POLYGON 256.005 44.895 256.015 44.895 256.005 44.885 ;
        POLYGON 256.945 44.895 256.945 44.885 256.935 44.885 ;
        RECT 256.945 44.885 258.010 44.900 ;
        RECT 255.135 44.875 255.890 44.885 ;
        RECT 253.460 44.855 254.135 44.875 ;
        POLYGON 253.410 44.855 253.410 44.850 253.405 44.850 ;
        RECT 253.410 44.850 254.135 44.855 ;
        POLYGON 253.405 44.850 253.405 44.840 253.390 44.840 ;
        RECT 253.405 44.840 254.135 44.850 ;
        RECT 247.135 44.835 252.680 44.840 ;
        POLYGON 252.680 44.840 252.690 44.840 252.680 44.835 ;
        POLYGON 253.390 44.840 253.390 44.835 253.385 44.835 ;
        RECT 253.390 44.835 254.135 44.840 ;
        RECT 247.135 44.820 252.625 44.835 ;
        RECT 245.535 44.785 246.355 44.820 ;
        POLYGON 246.355 44.820 246.405 44.785 246.355 44.785 ;
        POLYGON 247.135 44.820 247.150 44.820 247.150 44.815 ;
        RECT 247.150 44.815 252.625 44.820 ;
        POLYGON 247.150 44.815 247.210 44.815 247.210 44.785 ;
        RECT 247.210 44.805 252.625 44.815 ;
        POLYGON 252.625 44.835 252.680 44.835 252.625 44.805 ;
        POLYGON 253.385 44.835 253.385 44.805 253.340 44.805 ;
        RECT 253.385 44.805 254.135 44.835 ;
        RECT 247.210 44.785 252.545 44.805 ;
        RECT 245.535 44.770 246.405 44.785 ;
        RECT 243.650 44.755 244.625 44.770 ;
        RECT 241.240 44.645 242.525 44.745 ;
        POLYGON 243.650 44.755 243.660 44.755 243.660 44.740 ;
        RECT 243.660 44.740 244.625 44.755 ;
        POLYGON 242.525 44.740 242.605 44.645 242.525 44.645 ;
        POLYGON 243.660 44.740 243.695 44.740 243.695 44.700 ;
        RECT 243.695 44.705 244.625 44.740 ;
        POLYGON 244.625 44.770 244.695 44.705 244.625 44.705 ;
        POLYGON 245.535 44.770 245.615 44.770 245.615 44.710 ;
        RECT 245.615 44.730 246.405 44.770 ;
        POLYGON 246.405 44.785 246.480 44.730 246.405 44.730 ;
        POLYGON 247.210 44.785 247.275 44.785 247.275 44.755 ;
        RECT 247.275 44.765 252.545 44.785 ;
        POLYGON 252.545 44.805 252.625 44.805 252.545 44.765 ;
        POLYGON 253.340 44.805 253.340 44.765 253.280 44.765 ;
        RECT 253.340 44.785 254.135 44.805 ;
        POLYGON 254.135 44.875 254.235 44.875 254.135 44.785 ;
        POLYGON 255.115 44.875 255.115 44.785 255.025 44.785 ;
        RECT 255.115 44.785 255.890 44.875 ;
        RECT 253.340 44.765 254.095 44.785 ;
        RECT 247.275 44.755 252.460 44.765 ;
        POLYGON 247.275 44.755 247.330 44.755 247.330 44.730 ;
        RECT 247.330 44.730 252.460 44.755 ;
        RECT 245.615 44.725 246.480 44.730 ;
        POLYGON 246.480 44.730 246.490 44.725 246.480 44.725 ;
        POLYGON 247.330 44.730 247.345 44.730 247.345 44.725 ;
        RECT 247.345 44.725 252.460 44.730 ;
        RECT 245.615 44.710 246.490 44.725 ;
        POLYGON 245.615 44.710 245.620 44.710 245.620 44.705 ;
        RECT 245.620 44.705 246.490 44.710 ;
        RECT 243.695 44.700 244.695 44.705 ;
        POLYGON 244.695 44.705 244.700 44.700 244.695 44.700 ;
        POLYGON 245.620 44.705 245.630 44.705 245.630 44.700 ;
        RECT 245.630 44.700 246.490 44.705 ;
        POLYGON 243.695 44.700 243.745 44.700 243.745 44.645 ;
        RECT 243.745 44.680 244.700 44.700 ;
        POLYGON 244.700 44.700 244.725 44.680 244.700 44.680 ;
        POLYGON 245.630 44.700 245.640 44.700 245.640 44.695 ;
        RECT 245.640 44.695 246.490 44.700 ;
        POLYGON 245.640 44.695 245.660 44.695 245.660 44.680 ;
        RECT 245.660 44.680 246.490 44.695 ;
        RECT 243.745 44.645 244.725 44.680 ;
        RECT 241.240 44.605 242.605 44.645 ;
        POLYGON 242.605 44.645 242.635 44.605 242.605 44.605 ;
        RECT 241.240 44.600 242.635 44.605 ;
        POLYGON 243.745 44.645 243.790 44.645 243.790 44.600 ;
        RECT 243.790 44.600 244.725 44.645 ;
        POLYGON 244.725 44.680 244.810 44.600 244.725 44.600 ;
        POLYGON 245.660 44.680 245.765 44.680 245.765 44.600 ;
        RECT 245.765 44.660 246.490 44.680 ;
        POLYGON 246.490 44.725 246.590 44.660 246.490 44.660 ;
        POLYGON 247.345 44.725 247.415 44.725 247.415 44.695 ;
        RECT 247.415 44.720 252.460 44.725 ;
        POLYGON 252.460 44.765 252.545 44.765 252.460 44.720 ;
        POLYGON 253.280 44.765 253.280 44.745 253.250 44.745 ;
        RECT 253.280 44.755 254.095 44.765 ;
        POLYGON 254.095 44.785 254.135 44.785 254.095 44.755 ;
        POLYGON 255.025 44.785 255.025 44.755 254.995 44.755 ;
        RECT 255.025 44.755 255.890 44.785 ;
        RECT 253.280 44.745 253.995 44.755 ;
        POLYGON 253.250 44.745 253.250 44.740 253.245 44.740 ;
        RECT 253.250 44.740 253.995 44.745 ;
        POLYGON 253.245 44.740 253.245 44.720 253.215 44.720 ;
        RECT 253.245 44.720 253.995 44.740 ;
        RECT 247.415 44.710 252.435 44.720 ;
        POLYGON 252.435 44.720 252.460 44.720 252.435 44.710 ;
        POLYGON 253.215 44.720 253.215 44.710 253.200 44.710 ;
        RECT 253.215 44.710 253.995 44.720 ;
        RECT 247.415 44.695 252.395 44.710 ;
        POLYGON 247.415 44.695 247.495 44.695 247.495 44.660 ;
        RECT 247.495 44.690 252.395 44.695 ;
        POLYGON 252.395 44.710 252.430 44.710 252.395 44.690 ;
        POLYGON 253.200 44.710 253.200 44.705 253.195 44.705 ;
        RECT 253.200 44.705 253.995 44.710 ;
        POLYGON 253.195 44.705 253.195 44.690 253.170 44.690 ;
        RECT 253.195 44.690 253.995 44.705 ;
        RECT 247.495 44.660 252.295 44.690 ;
        RECT 245.765 44.625 246.590 44.660 ;
        POLYGON 246.590 44.660 246.645 44.625 246.590 44.625 ;
        POLYGON 247.495 44.660 247.555 44.660 247.555 44.635 ;
        RECT 247.555 44.645 252.295 44.660 ;
        POLYGON 252.295 44.690 252.395 44.690 252.295 44.645 ;
        POLYGON 253.170 44.690 253.170 44.655 253.115 44.655 ;
        RECT 253.170 44.675 253.995 44.690 ;
        POLYGON 253.995 44.755 254.095 44.755 253.995 44.675 ;
        POLYGON 254.995 44.755 254.995 44.675 254.915 44.675 ;
        RECT 254.995 44.740 255.890 44.755 ;
        POLYGON 255.890 44.885 256.005 44.885 255.890 44.740 ;
        POLYGON 256.935 44.885 256.935 44.765 256.855 44.765 ;
        RECT 256.935 44.800 258.010 44.885 ;
        POLYGON 258.010 45.015 258.140 45.015 258.010 44.800 ;
        POLYGON 259.585 45.015 259.585 44.815 259.495 44.815 ;
        RECT 259.585 44.815 261.085 45.015 ;
        POLYGON 259.495 44.815 259.495 44.800 259.485 44.800 ;
        RECT 259.495 44.800 261.085 44.815 ;
        RECT 256.935 44.765 257.975 44.800 ;
        POLYGON 256.855 44.765 256.855 44.745 256.840 44.745 ;
        RECT 256.855 44.745 257.975 44.765 ;
        RECT 254.995 44.675 255.765 44.740 ;
        RECT 253.170 44.655 253.900 44.675 ;
        POLYGON 253.115 44.655 253.115 44.645 253.100 44.645 ;
        RECT 253.115 44.645 253.900 44.655 ;
        RECT 247.555 44.635 252.245 44.645 ;
        POLYGON 247.555 44.635 247.575 44.635 247.575 44.625 ;
        RECT 247.575 44.625 252.245 44.635 ;
        RECT 245.765 44.600 246.645 44.625 ;
        POLYGON 246.645 44.625 246.680 44.600 246.645 44.600 ;
        POLYGON 247.575 44.625 247.615 44.625 247.615 44.610 ;
        RECT 247.615 44.620 252.245 44.625 ;
        POLYGON 252.245 44.645 252.295 44.645 252.245 44.620 ;
        POLYGON 253.100 44.645 253.100 44.640 253.095 44.640 ;
        RECT 253.100 44.640 253.900 44.645 ;
        POLYGON 253.095 44.640 253.095 44.620 253.065 44.620 ;
        RECT 253.095 44.620 253.900 44.640 ;
        RECT 247.615 44.610 252.195 44.620 ;
        POLYGON 247.615 44.610 247.645 44.610 247.645 44.600 ;
        RECT 247.645 44.600 252.195 44.610 ;
        POLYGON 252.195 44.620 252.245 44.620 252.195 44.600 ;
        POLYGON 253.065 44.620 253.065 44.600 253.030 44.600 ;
        RECT 253.065 44.600 253.900 44.620 ;
        POLYGON 253.900 44.675 253.995 44.675 253.900 44.600 ;
        POLYGON 254.915 44.675 254.915 44.600 254.840 44.600 ;
        RECT 254.915 44.600 255.765 44.675 ;
        POLYGON 255.765 44.740 255.890 44.740 255.765 44.600 ;
        POLYGON 256.840 44.740 256.840 44.720 256.825 44.720 ;
        RECT 256.840 44.735 257.975 44.745 ;
        POLYGON 257.975 44.800 258.010 44.800 257.975 44.735 ;
        POLYGON 259.485 44.795 259.485 44.740 259.455 44.740 ;
        RECT 259.485 44.740 261.085 44.800 ;
        POLYGON 261.085 45.095 261.250 45.095 261.085 44.740 ;
        POLYGON 263.465 45.095 263.465 45.080 263.460 45.080 ;
        RECT 263.465 45.080 266.230 45.100 ;
        POLYGON 263.460 45.080 263.460 44.845 263.385 44.845 ;
        RECT 263.460 44.845 266.230 45.080 ;
        POLYGON 263.385 44.845 263.385 44.740 263.350 44.740 ;
        RECT 263.385 44.740 266.230 44.845 ;
        RECT 256.840 44.720 257.935 44.735 ;
        POLYGON 256.825 44.720 256.825 44.645 256.765 44.645 ;
        RECT 256.825 44.680 257.935 44.720 ;
        POLYGON 257.935 44.735 257.975 44.735 257.935 44.680 ;
        POLYGON 259.455 44.735 259.455 44.680 259.425 44.680 ;
        RECT 259.455 44.700 261.070 44.740 ;
        POLYGON 261.070 44.740 261.085 44.740 261.070 44.700 ;
        POLYGON 263.350 44.730 263.350 44.700 263.340 44.700 ;
        RECT 263.350 44.700 266.230 44.740 ;
        RECT 259.455 44.680 261.025 44.700 ;
        RECT 256.825 44.645 257.885 44.680 ;
        POLYGON 256.765 44.645 256.765 44.630 256.755 44.630 ;
        RECT 256.765 44.630 257.885 44.645 ;
        POLYGON 256.755 44.630 256.755 44.600 256.730 44.600 ;
        RECT 256.755 44.600 257.885 44.630 ;
        POLYGON 257.885 44.680 257.935 44.680 257.885 44.600 ;
        POLYGON 259.425 44.680 259.425 44.635 259.400 44.635 ;
        RECT 259.425 44.635 261.025 44.680 ;
        POLYGON 259.400 44.630 259.400 44.600 259.385 44.600 ;
        RECT 259.400 44.600 261.025 44.635 ;
        POLYGON 261.025 44.700 261.070 44.700 261.025 44.605 ;
        POLYGON 263.340 44.700 263.340 44.605 263.310 44.605 ;
        RECT 263.340 44.670 266.230 44.700 ;
        POLYGON 266.230 45.255 266.365 45.255 266.230 44.670 ;
        POLYGON 270.645 45.255 270.645 44.710 270.610 44.710 ;
        RECT 270.645 44.710 277.820 45.295 ;
        RECT 263.340 44.605 266.210 44.670 ;
        POLYGON 208.330 44.600 208.495 44.600 208.495 44.100 ;
        RECT 208.495 44.095 223.280 44.600 ;
        POLYGON 223.280 44.600 223.450 44.095 223.280 44.095 ;
        POLYGON 230.335 44.600 230.505 44.600 230.505 44.125 ;
        RECT 230.505 44.505 234.525 44.600 ;
        POLYGON 234.525 44.600 234.570 44.505 234.525 44.505 ;
        POLYGON 237.410 44.600 237.460 44.600 237.460 44.510 ;
        RECT 237.460 44.590 239.545 44.600 ;
        POLYGON 239.545 44.600 239.550 44.590 239.545 44.590 ;
        POLYGON 241.240 44.600 241.245 44.600 241.245 44.590 ;
        RECT 241.245 44.590 242.635 44.600 ;
        RECT 237.460 44.580 239.550 44.590 ;
        POLYGON 239.550 44.590 239.560 44.580 239.550 44.580 ;
        POLYGON 241.245 44.590 241.250 44.590 241.250 44.585 ;
        RECT 241.250 44.580 242.635 44.590 ;
        RECT 237.460 44.560 239.560 44.580 ;
        POLYGON 239.560 44.580 239.570 44.560 239.560 44.560 ;
        POLYGON 241.250 44.580 241.265 44.580 241.265 44.560 ;
        RECT 241.265 44.560 242.635 44.580 ;
        RECT 237.460 44.530 239.570 44.560 ;
        POLYGON 239.570 44.560 239.590 44.530 239.570 44.530 ;
        POLYGON 241.265 44.560 241.270 44.560 241.270 44.555 ;
        RECT 241.270 44.555 242.635 44.560 ;
        POLYGON 241.270 44.555 241.285 44.555 241.285 44.530 ;
        RECT 241.285 44.540 242.635 44.555 ;
        POLYGON 242.635 44.600 242.685 44.540 242.635 44.540 ;
        POLYGON 243.790 44.600 243.850 44.600 243.850 44.540 ;
        RECT 243.850 44.550 244.810 44.600 ;
        POLYGON 244.810 44.600 244.865 44.550 244.810 44.550 ;
        POLYGON 245.765 44.600 245.820 44.600 245.820 44.560 ;
        RECT 245.820 44.560 246.680 44.600 ;
        POLYGON 245.820 44.560 245.840 44.560 245.840 44.550 ;
        RECT 245.840 44.550 246.680 44.560 ;
        RECT 243.850 44.540 244.865 44.550 ;
        RECT 241.285 44.535 242.685 44.540 ;
        POLYGON 242.685 44.540 242.690 44.535 242.685 44.535 ;
        POLYGON 243.850 44.540 243.855 44.540 243.855 44.535 ;
        RECT 243.855 44.535 244.865 44.540 ;
        RECT 241.285 44.530 242.690 44.535 ;
        RECT 237.460 44.505 239.590 44.530 ;
        RECT 230.505 44.125 234.570 44.505 ;
        POLYGON 230.505 44.125 230.515 44.125 230.515 44.095 ;
        RECT 230.515 44.115 234.570 44.125 ;
        POLYGON 234.570 44.505 234.740 44.115 234.570 44.115 ;
        POLYGON 237.460 44.505 237.670 44.505 237.670 44.125 ;
        RECT 237.670 44.480 239.590 44.505 ;
        POLYGON 239.590 44.530 239.615 44.480 239.590 44.480 ;
        POLYGON 241.285 44.530 241.320 44.530 241.320 44.485 ;
        RECT 241.320 44.480 242.690 44.530 ;
        RECT 237.670 44.420 239.615 44.480 ;
        POLYGON 239.615 44.480 239.650 44.420 239.615 44.420 ;
        POLYGON 241.320 44.480 241.365 44.480 241.365 44.420 ;
        RECT 241.365 44.420 242.690 44.480 ;
        RECT 237.670 44.345 239.655 44.420 ;
        POLYGON 241.365 44.420 241.370 44.420 241.370 44.415 ;
        RECT 241.370 44.415 242.690 44.420 ;
        POLYGON 239.655 44.415 239.695 44.345 239.655 44.345 ;
        POLYGON 241.370 44.415 241.420 44.415 241.420 44.345 ;
        RECT 241.420 44.350 242.690 44.415 ;
        POLYGON 242.690 44.535 242.850 44.350 242.690 44.350 ;
        POLYGON 243.855 44.535 243.870 44.535 243.870 44.520 ;
        RECT 243.870 44.530 244.865 44.535 ;
        POLYGON 244.865 44.550 244.890 44.530 244.865 44.530 ;
        POLYGON 245.840 44.550 245.845 44.550 245.845 44.545 ;
        RECT 245.845 44.545 246.680 44.550 ;
        POLYGON 245.845 44.545 245.865 44.545 245.865 44.530 ;
        RECT 245.865 44.530 246.680 44.545 ;
        RECT 243.870 44.520 244.890 44.530 ;
        POLYGON 243.870 44.520 244.015 44.520 244.015 44.370 ;
        RECT 244.015 44.400 244.890 44.520 ;
        POLYGON 244.890 44.530 245.040 44.400 244.890 44.400 ;
        POLYGON 245.865 44.530 246.035 44.530 246.035 44.415 ;
        RECT 246.035 44.500 246.680 44.530 ;
        POLYGON 246.680 44.600 246.830 44.500 246.680 44.500 ;
        POLYGON 247.645 44.600 247.690 44.600 247.690 44.585 ;
        RECT 247.690 44.595 252.180 44.600 ;
        POLYGON 252.180 44.600 252.195 44.600 252.180 44.595 ;
        POLYGON 253.030 44.600 253.030 44.595 253.025 44.595 ;
        RECT 253.030 44.595 253.880 44.600 ;
        RECT 247.690 44.585 252.125 44.595 ;
        POLYGON 247.690 44.585 247.830 44.585 247.830 44.535 ;
        RECT 247.830 44.570 252.125 44.585 ;
        POLYGON 252.125 44.595 252.180 44.595 252.125 44.570 ;
        POLYGON 253.025 44.595 253.025 44.570 252.985 44.570 ;
        RECT 253.025 44.585 253.880 44.595 ;
        POLYGON 253.880 44.600 253.900 44.600 253.880 44.585 ;
        POLYGON 254.840 44.600 254.840 44.585 254.820 44.585 ;
        RECT 254.840 44.585 255.740 44.600 ;
        RECT 253.025 44.575 253.870 44.585 ;
        POLYGON 253.870 44.585 253.880 44.585 253.870 44.575 ;
        POLYGON 254.820 44.585 254.820 44.575 254.810 44.575 ;
        RECT 254.820 44.575 255.740 44.585 ;
        RECT 253.025 44.570 253.750 44.575 ;
        RECT 247.830 44.535 251.950 44.570 ;
        POLYGON 247.830 44.535 247.895 44.535 247.895 44.510 ;
        RECT 247.895 44.510 251.950 44.535 ;
        POLYGON 247.895 44.510 247.925 44.510 247.925 44.500 ;
        RECT 247.925 44.505 251.950 44.510 ;
        POLYGON 251.950 44.570 252.125 44.570 251.950 44.505 ;
        POLYGON 252.985 44.570 252.985 44.565 252.975 44.565 ;
        RECT 252.985 44.565 253.750 44.570 ;
        POLYGON 252.975 44.565 252.975 44.545 252.940 44.545 ;
        RECT 252.975 44.545 253.750 44.565 ;
        POLYGON 252.940 44.545 252.940 44.535 252.930 44.535 ;
        RECT 252.940 44.535 253.750 44.545 ;
        POLYGON 252.930 44.535 252.930 44.505 252.880 44.505 ;
        RECT 252.930 44.505 253.750 44.535 ;
        RECT 247.925 44.500 251.935 44.505 ;
        POLYGON 251.935 44.505 251.950 44.505 251.935 44.500 ;
        POLYGON 252.880 44.505 252.880 44.500 252.870 44.500 ;
        RECT 252.880 44.500 253.750 44.505 ;
        RECT 246.035 44.465 246.830 44.500 ;
        POLYGON 246.830 44.500 246.885 44.465 246.830 44.465 ;
        POLYGON 247.925 44.500 247.970 44.500 247.970 44.485 ;
        RECT 247.970 44.495 251.925 44.500 ;
        POLYGON 251.925 44.500 251.935 44.500 251.925 44.495 ;
        POLYGON 252.870 44.500 252.870 44.495 252.865 44.495 ;
        RECT 252.870 44.495 253.750 44.500 ;
        RECT 247.970 44.485 251.775 44.495 ;
        POLYGON 247.975 44.485 248.040 44.485 248.040 44.465 ;
        RECT 248.040 44.465 251.775 44.485 ;
        RECT 246.035 44.415 246.890 44.465 ;
        POLYGON 246.035 44.415 246.055 44.415 246.055 44.405 ;
        RECT 246.055 44.405 246.890 44.415 ;
        POLYGON 246.055 44.405 246.060 44.405 246.060 44.400 ;
        RECT 246.060 44.400 246.890 44.405 ;
        POLYGON 246.890 44.465 247.000 44.400 246.890 44.400 ;
        POLYGON 248.040 44.465 248.180 44.465 248.180 44.425 ;
        RECT 248.180 44.445 251.775 44.465 ;
        POLYGON 251.775 44.495 251.920 44.495 251.775 44.445 ;
        POLYGON 252.865 44.495 252.865 44.475 252.830 44.475 ;
        RECT 252.865 44.490 253.750 44.495 ;
        POLYGON 253.750 44.575 253.870 44.575 253.750 44.490 ;
        POLYGON 254.810 44.575 254.810 44.525 254.755 44.525 ;
        RECT 254.810 44.570 255.740 44.575 ;
        POLYGON 255.740 44.600 255.765 44.600 255.740 44.570 ;
        POLYGON 256.730 44.600 256.730 44.580 256.715 44.580 ;
        RECT 256.730 44.580 257.795 44.600 ;
        POLYGON 256.715 44.580 256.715 44.575 256.710 44.575 ;
        RECT 256.715 44.575 257.795 44.580 ;
        RECT 254.810 44.560 255.735 44.570 ;
        POLYGON 255.735 44.570 255.740 44.570 255.735 44.560 ;
        POLYGON 256.710 44.570 256.710 44.560 256.700 44.560 ;
        RECT 256.710 44.560 257.795 44.575 ;
        RECT 254.810 44.525 255.695 44.560 ;
        POLYGON 254.755 44.525 254.755 44.505 254.730 44.505 ;
        RECT 254.755 44.515 255.695 44.525 ;
        POLYGON 255.695 44.560 255.735 44.560 255.695 44.515 ;
        POLYGON 256.700 44.560 256.700 44.515 256.665 44.515 ;
        RECT 256.700 44.515 257.795 44.560 ;
        RECT 254.755 44.505 255.495 44.515 ;
        POLYGON 254.730 44.505 254.730 44.490 254.715 44.490 ;
        RECT 254.730 44.490 255.495 44.505 ;
        RECT 252.865 44.475 253.640 44.490 ;
        POLYGON 252.830 44.475 252.830 44.450 252.790 44.450 ;
        RECT 252.830 44.450 253.640 44.475 ;
        POLYGON 252.790 44.450 252.790 44.445 252.785 44.445 ;
        RECT 252.790 44.445 253.640 44.450 ;
        RECT 248.180 44.425 251.660 44.445 ;
        POLYGON 248.180 44.425 248.265 44.425 248.265 44.400 ;
        RECT 248.265 44.410 251.660 44.425 ;
        POLYGON 251.660 44.445 251.775 44.445 251.660 44.410 ;
        POLYGON 252.785 44.445 252.785 44.410 252.720 44.410 ;
        RECT 252.785 44.410 253.640 44.445 ;
        POLYGON 253.640 44.490 253.750 44.490 253.640 44.410 ;
        POLYGON 254.715 44.490 254.715 44.485 254.710 44.485 ;
        RECT 254.715 44.485 255.495 44.490 ;
        POLYGON 254.710 44.485 254.710 44.410 254.625 44.410 ;
        RECT 254.710 44.410 255.495 44.485 ;
        RECT 248.265 44.400 251.615 44.410 ;
        RECT 244.015 44.380 245.040 44.400 ;
        POLYGON 245.040 44.400 245.065 44.380 245.040 44.380 ;
        POLYGON 246.060 44.400 246.095 44.400 246.095 44.380 ;
        RECT 246.095 44.380 247.000 44.400 ;
        RECT 244.015 44.370 245.065 44.380 ;
        POLYGON 244.015 44.370 244.035 44.370 244.035 44.350 ;
        RECT 244.035 44.355 245.065 44.370 ;
        POLYGON 245.065 44.380 245.090 44.355 245.065 44.355 ;
        POLYGON 246.095 44.380 246.135 44.380 246.135 44.355 ;
        RECT 246.135 44.355 247.000 44.380 ;
        POLYGON 247.000 44.400 247.085 44.355 247.000 44.355 ;
        POLYGON 248.265 44.400 248.390 44.400 248.390 44.370 ;
        RECT 248.390 44.395 251.615 44.400 ;
        POLYGON 251.615 44.410 251.660 44.410 251.615 44.395 ;
        POLYGON 252.720 44.410 252.720 44.395 252.690 44.395 ;
        RECT 252.720 44.395 253.620 44.410 ;
        POLYGON 253.620 44.410 253.640 44.410 253.620 44.395 ;
        POLYGON 254.625 44.410 254.625 44.395 254.610 44.395 ;
        RECT 254.625 44.395 255.495 44.410 ;
        RECT 248.390 44.390 251.595 44.395 ;
        POLYGON 251.595 44.395 251.610 44.395 251.595 44.390 ;
        POLYGON 252.690 44.395 252.690 44.390 252.680 44.390 ;
        RECT 252.690 44.390 253.505 44.395 ;
        RECT 248.390 44.370 251.410 44.390 ;
        POLYGON 248.390 44.370 248.450 44.370 248.450 44.355 ;
        RECT 248.450 44.355 251.410 44.370 ;
        RECT 244.035 44.350 245.090 44.355 ;
        RECT 241.420 44.345 242.850 44.350 ;
        RECT 237.670 44.310 239.695 44.345 ;
        POLYGON 239.695 44.345 239.720 44.310 239.695 44.310 ;
        POLYGON 241.420 44.345 241.445 44.345 241.445 44.310 ;
        RECT 241.445 44.340 242.850 44.345 ;
        POLYGON 242.850 44.350 242.860 44.340 242.850 44.340 ;
        POLYGON 244.035 44.350 244.045 44.350 244.045 44.340 ;
        RECT 244.045 44.340 245.090 44.350 ;
        RECT 241.445 44.315 242.860 44.340 ;
        POLYGON 242.860 44.340 242.880 44.315 242.860 44.315 ;
        POLYGON 244.045 44.340 244.070 44.340 244.070 44.315 ;
        RECT 244.070 44.315 245.090 44.340 ;
        RECT 241.445 44.310 242.880 44.315 ;
        RECT 237.670 44.265 239.720 44.310 ;
        POLYGON 239.720 44.310 239.745 44.265 239.720 44.265 ;
        POLYGON 241.445 44.310 241.465 44.310 241.465 44.285 ;
        RECT 241.465 44.285 242.880 44.310 ;
        POLYGON 241.465 44.285 241.480 44.285 241.480 44.270 ;
        RECT 241.480 44.265 242.880 44.285 ;
        RECT 237.670 44.245 239.745 44.265 ;
        POLYGON 239.745 44.265 239.760 44.245 239.745 44.245 ;
        POLYGON 241.480 44.265 241.495 44.265 241.495 44.245 ;
        RECT 241.495 44.245 242.880 44.265 ;
        RECT 237.670 44.175 239.760 44.245 ;
        POLYGON 239.760 44.245 239.805 44.175 239.760 44.175 ;
        POLYGON 241.495 44.245 241.545 44.245 241.545 44.175 ;
        RECT 241.545 44.200 242.880 44.245 ;
        POLYGON 242.880 44.315 242.975 44.200 242.880 44.200 ;
        POLYGON 244.070 44.315 244.100 44.315 244.100 44.290 ;
        RECT 244.100 44.290 245.090 44.315 ;
        POLYGON 244.100 44.290 244.195 44.290 244.195 44.200 ;
        RECT 244.195 44.250 245.090 44.290 ;
        POLYGON 245.090 44.355 245.225 44.250 245.090 44.250 ;
        POLYGON 246.135 44.355 246.240 44.355 246.240 44.290 ;
        RECT 246.240 44.320 247.085 44.355 ;
        POLYGON 247.085 44.355 247.150 44.320 247.085 44.320 ;
        POLYGON 248.450 44.355 248.475 44.355 248.475 44.350 ;
        RECT 248.475 44.350 251.410 44.355 ;
        POLYGON 248.475 44.350 248.565 44.350 248.565 44.330 ;
        RECT 248.565 44.340 251.410 44.350 ;
        POLYGON 251.410 44.390 251.595 44.390 251.410 44.340 ;
        POLYGON 252.680 44.390 252.680 44.360 252.625 44.360 ;
        RECT 252.680 44.360 253.505 44.390 ;
        POLYGON 252.625 44.360 252.625 44.340 252.590 44.340 ;
        RECT 252.625 44.340 253.505 44.360 ;
        RECT 248.565 44.330 251.275 44.340 ;
        POLYGON 248.565 44.330 248.615 44.330 248.615 44.320 ;
        RECT 248.615 44.320 251.275 44.330 ;
        RECT 246.240 44.290 247.150 44.320 ;
        POLYGON 246.240 44.290 246.260 44.290 246.260 44.280 ;
        RECT 246.260 44.280 247.150 44.290 ;
        POLYGON 246.260 44.280 246.275 44.280 246.275 44.270 ;
        RECT 246.275 44.270 247.150 44.280 ;
        POLYGON 246.275 44.270 246.310 44.270 246.310 44.250 ;
        RECT 246.310 44.250 247.150 44.270 ;
        RECT 244.195 44.230 245.225 44.250 ;
        POLYGON 245.225 44.250 245.250 44.230 245.225 44.230 ;
        POLYGON 246.310 44.250 246.345 44.250 246.345 44.230 ;
        RECT 246.345 44.245 247.150 44.250 ;
        POLYGON 247.150 44.320 247.275 44.245 247.150 44.245 ;
        POLYGON 248.615 44.320 248.665 44.320 248.665 44.310 ;
        RECT 248.665 44.310 251.275 44.320 ;
        POLYGON 251.275 44.340 251.400 44.340 251.275 44.310 ;
        POLYGON 252.590 44.340 252.590 44.315 252.545 44.315 ;
        RECT 252.590 44.320 253.505 44.340 ;
        POLYGON 253.505 44.395 253.620 44.395 253.505 44.320 ;
        POLYGON 254.610 44.395 254.610 44.370 254.580 44.370 ;
        RECT 254.610 44.370 255.495 44.395 ;
        POLYGON 254.580 44.370 254.580 44.325 254.525 44.325 ;
        RECT 254.580 44.325 255.495 44.370 ;
        POLYGON 254.525 44.325 254.525 44.320 254.520 44.320 ;
        RECT 254.525 44.320 255.495 44.325 ;
        RECT 252.590 44.315 253.410 44.320 ;
        POLYGON 252.540 44.315 252.540 44.310 252.530 44.310 ;
        RECT 252.540 44.310 253.410 44.315 ;
        POLYGON 248.665 44.310 248.775 44.310 248.775 44.285 ;
        RECT 248.775 44.295 251.225 44.310 ;
        POLYGON 251.225 44.310 251.275 44.310 251.225 44.295 ;
        POLYGON 252.530 44.310 252.530 44.295 252.505 44.295 ;
        RECT 252.530 44.295 253.410 44.310 ;
        RECT 248.775 44.285 251.135 44.295 ;
        POLYGON 248.775 44.285 248.870 44.285 248.870 44.270 ;
        RECT 248.870 44.280 251.135 44.285 ;
        POLYGON 251.135 44.295 251.225 44.295 251.135 44.280 ;
        POLYGON 252.505 44.295 252.505 44.280 252.480 44.280 ;
        RECT 252.505 44.280 253.410 44.295 ;
        RECT 248.870 44.270 251.035 44.280 ;
        POLYGON 248.875 44.270 248.940 44.270 248.940 44.260 ;
        RECT 248.940 44.260 251.035 44.270 ;
        POLYGON 251.035 44.280 251.135 44.280 251.035 44.260 ;
        POLYGON 252.480 44.280 252.480 44.270 252.460 44.270 ;
        RECT 252.480 44.270 253.410 44.280 ;
        POLYGON 252.460 44.270 252.460 44.260 252.445 44.260 ;
        RECT 252.460 44.260 253.410 44.270 ;
        POLYGON 248.945 44.260 249.050 44.260 249.050 44.245 ;
        RECT 249.050 44.245 250.930 44.260 ;
        POLYGON 250.930 44.260 251.035 44.260 250.930 44.245 ;
        POLYGON 252.445 44.260 252.445 44.255 252.435 44.255 ;
        RECT 252.445 44.255 253.410 44.260 ;
        POLYGON 253.410 44.320 253.505 44.320 253.410 44.255 ;
        POLYGON 254.520 44.320 254.520 44.280 254.475 44.280 ;
        RECT 254.520 44.300 255.495 44.320 ;
        POLYGON 255.495 44.515 255.695 44.515 255.495 44.300 ;
        POLYGON 256.665 44.510 256.665 44.430 256.605 44.430 ;
        RECT 256.665 44.460 257.795 44.515 ;
        POLYGON 257.795 44.600 257.885 44.600 257.795 44.460 ;
        POLYGON 259.385 44.600 259.385 44.570 259.370 44.570 ;
        RECT 259.385 44.570 260.945 44.600 ;
        POLYGON 259.365 44.570 259.365 44.510 259.335 44.510 ;
        RECT 259.365 44.510 260.945 44.570 ;
        POLYGON 259.335 44.510 259.335 44.465 259.310 44.465 ;
        RECT 259.335 44.465 260.945 44.510 ;
        RECT 256.665 44.430 257.615 44.460 ;
        POLYGON 256.605 44.430 256.605 44.385 256.570 44.385 ;
        RECT 256.605 44.385 257.615 44.430 ;
        POLYGON 256.570 44.385 256.570 44.330 256.525 44.330 ;
        RECT 256.570 44.330 257.615 44.385 ;
        POLYGON 256.525 44.330 256.525 44.320 256.515 44.320 ;
        RECT 256.525 44.320 257.615 44.330 ;
        POLYGON 256.515 44.320 256.515 44.300 256.500 44.300 ;
        RECT 256.515 44.300 257.615 44.320 ;
        RECT 254.520 44.280 255.460 44.300 ;
        POLYGON 254.475 44.280 254.475 44.255 254.445 44.255 ;
        RECT 254.475 44.260 255.460 44.280 ;
        POLYGON 255.460 44.300 255.495 44.300 255.460 44.260 ;
        POLYGON 256.500 44.300 256.500 44.260 256.465 44.260 ;
        RECT 256.500 44.260 257.615 44.300 ;
        RECT 254.475 44.255 255.295 44.260 ;
        POLYGON 252.430 44.255 252.430 44.245 252.415 44.245 ;
        RECT 252.430 44.245 253.355 44.255 ;
        RECT 246.345 44.230 247.275 44.245 ;
        RECT 244.195 44.200 245.250 44.230 ;
        RECT 241.545 44.175 242.975 44.200 ;
        RECT 237.670 44.140 239.805 44.175 ;
        POLYGON 239.805 44.175 239.830 44.140 239.805 44.140 ;
        POLYGON 241.545 44.175 241.560 44.175 241.560 44.155 ;
        RECT 241.560 44.155 242.975 44.175 ;
        POLYGON 241.560 44.155 241.570 44.155 241.570 44.140 ;
        RECT 241.570 44.140 242.975 44.155 ;
        RECT 237.670 44.125 239.830 44.140 ;
        POLYGON 237.670 44.125 237.675 44.125 237.675 44.115 ;
        RECT 237.675 44.115 239.830 44.125 ;
        RECT 230.515 44.100 234.740 44.115 ;
        POLYGON 234.740 44.115 234.745 44.100 234.740 44.100 ;
        RECT 230.515 44.095 234.745 44.100 ;
        POLYGON 237.675 44.115 237.685 44.115 237.685 44.095 ;
        RECT 237.685 44.100 239.830 44.115 ;
        POLYGON 239.830 44.140 239.855 44.100 239.830 44.100 ;
        RECT 237.685 44.095 239.855 44.100 ;
        POLYGON 241.570 44.140 241.605 44.140 241.605 44.095 ;
        RECT 241.605 44.130 242.975 44.140 ;
        POLYGON 242.975 44.200 243.040 44.130 242.975 44.130 ;
        POLYGON 244.195 44.200 244.270 44.200 244.270 44.130 ;
        RECT 244.270 44.175 245.250 44.200 ;
        POLYGON 245.250 44.230 245.320 44.175 245.250 44.175 ;
        POLYGON 246.345 44.230 246.445 44.230 246.445 44.175 ;
        RECT 246.445 44.175 247.275 44.230 ;
        RECT 244.270 44.130 245.320 44.175 ;
        RECT 241.605 44.095 243.040 44.130 ;
        POLYGON 243.040 44.130 243.070 44.095 243.040 44.095 ;
        POLYGON 244.270 44.130 244.310 44.130 244.310 44.095 ;
        RECT 244.310 44.105 245.320 44.130 ;
        POLYGON 245.320 44.175 245.415 44.105 245.320 44.105 ;
        POLYGON 246.445 44.175 246.490 44.175 246.490 44.150 ;
        RECT 246.490 44.150 247.275 44.175 ;
        POLYGON 246.490 44.150 246.505 44.150 246.505 44.140 ;
        RECT 246.505 44.140 247.275 44.150 ;
        POLYGON 246.505 44.140 246.570 44.140 246.570 44.105 ;
        RECT 246.570 44.125 247.275 44.140 ;
        POLYGON 247.275 44.245 247.515 44.125 247.275 44.125 ;
        POLYGON 249.050 44.245 249.190 44.245 249.190 44.225 ;
        RECT 249.190 44.235 250.865 44.245 ;
        POLYGON 250.865 44.245 250.925 44.245 250.865 44.235 ;
        POLYGON 252.415 44.245 252.415 44.235 252.395 44.235 ;
        RECT 252.415 44.235 253.355 44.245 ;
        RECT 249.190 44.230 250.845 44.235 ;
        POLYGON 250.845 44.235 250.865 44.235 250.845 44.230 ;
        POLYGON 252.395 44.235 252.395 44.230 252.385 44.230 ;
        RECT 252.395 44.230 253.355 44.235 ;
        RECT 249.190 44.225 250.650 44.230 ;
        POLYGON 249.225 44.225 249.400 44.225 249.400 44.205 ;
        RECT 249.400 44.205 250.650 44.225 ;
        POLYGON 250.650 44.230 250.845 44.230 250.650 44.205 ;
        POLYGON 252.385 44.230 252.385 44.220 252.370 44.220 ;
        RECT 252.385 44.220 253.355 44.230 ;
        POLYGON 253.355 44.255 253.410 44.255 253.355 44.220 ;
        POLYGON 254.445 44.255 254.445 44.220 254.400 44.220 ;
        RECT 254.445 44.220 255.295 44.255 ;
        POLYGON 252.370 44.220 252.370 44.205 252.340 44.205 ;
        RECT 252.370 44.205 253.260 44.220 ;
        POLYGON 249.400 44.205 249.490 44.205 249.490 44.200 ;
        RECT 249.490 44.200 250.595 44.205 ;
        POLYGON 250.595 44.205 250.650 44.205 250.595 44.200 ;
        POLYGON 252.340 44.205 252.340 44.200 252.325 44.200 ;
        RECT 252.340 44.200 253.260 44.205 ;
        POLYGON 249.500 44.200 249.505 44.200 249.505 44.195 ;
        RECT 249.505 44.195 250.455 44.200 ;
        POLYGON 249.515 44.195 249.725 44.195 249.725 44.180 ;
        RECT 249.725 44.190 250.455 44.195 ;
        POLYGON 250.455 44.200 250.560 44.200 250.455 44.190 ;
        POLYGON 252.325 44.200 252.325 44.190 252.305 44.190 ;
        RECT 252.325 44.190 253.260 44.200 ;
        RECT 249.725 44.180 250.325 44.190 ;
        POLYGON 250.325 44.190 250.455 44.190 250.325 44.180 ;
        POLYGON 252.305 44.190 252.305 44.180 252.285 44.180 ;
        RECT 252.305 44.180 253.260 44.190 ;
        POLYGON 249.845 44.180 250.010 44.180 250.010 44.175 ;
        RECT 250.010 44.175 250.180 44.180 ;
        POLYGON 250.180 44.180 250.255 44.180 250.180 44.175 ;
        POLYGON 252.285 44.180 252.285 44.175 252.275 44.175 ;
        RECT 252.285 44.175 253.260 44.180 ;
        POLYGON 252.275 44.175 252.275 44.160 252.245 44.160 ;
        RECT 252.275 44.160 253.260 44.175 ;
        POLYGON 253.260 44.220 253.355 44.220 253.260 44.160 ;
        POLYGON 254.400 44.220 254.400 44.205 254.380 44.205 ;
        RECT 254.400 44.205 255.295 44.220 ;
        POLYGON 254.380 44.205 254.380 44.160 254.315 44.160 ;
        RECT 254.380 44.160 255.295 44.205 ;
        POLYGON 252.240 44.160 252.240 44.125 252.170 44.125 ;
        RECT 252.240 44.125 253.170 44.160 ;
        RECT 246.570 44.110 247.515 44.125 ;
        POLYGON 247.515 44.125 247.555 44.110 247.515 44.110 ;
        POLYGON 252.170 44.125 252.170 44.120 252.160 44.120 ;
        RECT 252.170 44.120 253.170 44.125 ;
        POLYGON 252.160 44.120 252.160 44.110 252.145 44.110 ;
        RECT 252.160 44.110 253.170 44.120 ;
        POLYGON 253.170 44.160 253.260 44.160 253.170 44.110 ;
        POLYGON 254.315 44.160 254.315 44.155 254.310 44.155 ;
        RECT 254.315 44.155 255.295 44.160 ;
        POLYGON 254.310 44.155 254.310 44.110 254.255 44.110 ;
        RECT 254.310 44.110 255.295 44.155 ;
        RECT 246.570 44.105 247.555 44.110 ;
        RECT 244.310 44.095 245.415 44.105 ;
        POLYGON 245.415 44.105 245.425 44.095 245.415 44.095 ;
        POLYGON 246.570 44.105 246.585 44.105 246.585 44.095 ;
        RECT 246.585 44.095 247.555 44.105 ;
        RECT 182.810 44.075 198.035 44.095 ;
        POLYGON 182.795 44.075 182.795 44.045 182.790 44.045 ;
        RECT 182.795 44.045 198.035 44.075 ;
        RECT 171.180 43.940 175.530 44.045 ;
        RECT 165.750 43.930 167.950 43.940 ;
        RECT 162.440 43.910 163.940 43.930 ;
        POLYGON 162.410 43.910 162.410 43.795 162.325 43.795 ;
        RECT 162.410 43.830 163.940 43.910 ;
        POLYGON 163.940 43.930 164.010 43.930 163.940 43.830 ;
        POLYGON 165.700 43.925 165.700 43.915 165.695 43.915 ;
        RECT 165.700 43.915 167.950 43.930 ;
        POLYGON 165.695 43.915 165.695 43.890 165.675 43.890 ;
        RECT 165.695 43.890 167.950 43.915 ;
        POLYGON 165.675 43.890 165.675 43.835 165.645 43.835 ;
        RECT 165.675 43.835 167.950 43.890 ;
        RECT 162.410 43.795 163.735 43.830 ;
        POLYGON 162.325 43.795 162.325 43.715 162.255 43.715 ;
        RECT 162.325 43.715 163.735 43.795 ;
        RECT 159.940 43.635 160.860 43.710 ;
        RECT 157.210 43.630 158.505 43.635 ;
        POLYGON 157.170 43.630 157.170 43.625 157.160 43.625 ;
        RECT 157.170 43.625 158.505 43.630 ;
        POLYGON 157.150 43.625 157.150 43.610 157.110 43.610 ;
        RECT 157.150 43.610 158.505 43.625 ;
        POLYGON 158.505 43.635 158.550 43.635 158.505 43.610 ;
        POLYGON 159.785 43.635 159.785 43.610 159.760 43.610 ;
        RECT 159.785 43.610 160.860 43.635 ;
        RECT 151.175 43.600 152.690 43.610 ;
        POLYGON 152.690 43.610 152.715 43.600 152.690 43.600 ;
        POLYGON 153.995 43.610 154.005 43.610 154.005 43.605 ;
        RECT 154.005 43.605 155.565 43.610 ;
        POLYGON 154.005 43.605 154.035 43.605 154.035 43.600 ;
        RECT 154.035 43.600 155.565 43.605 ;
        RECT 151.175 43.570 152.720 43.600 ;
        RECT 117.295 43.540 151.050 43.570 ;
        POLYGON 151.050 43.570 151.065 43.540 151.050 43.540 ;
        POLYGON 151.175 43.570 151.225 43.570 151.225 43.540 ;
        RECT 151.225 43.565 152.720 43.570 ;
        POLYGON 152.720 43.600 152.820 43.565 152.720 43.565 ;
        POLYGON 154.035 43.600 154.125 43.600 154.125 43.585 ;
        RECT 154.125 43.590 155.565 43.600 ;
        POLYGON 155.565 43.610 155.660 43.610 155.565 43.590 ;
        POLYGON 157.110 43.610 157.110 43.590 157.055 43.590 ;
        RECT 157.110 43.590 158.355 43.610 ;
        RECT 154.125 43.585 155.545 43.590 ;
        POLYGON 155.545 43.590 155.565 43.590 155.545 43.585 ;
        POLYGON 157.055 43.590 157.055 43.585 157.045 43.585 ;
        RECT 157.055 43.585 158.355 43.590 ;
        POLYGON 154.130 43.585 154.220 43.585 154.220 43.570 ;
        RECT 154.220 43.570 155.455 43.585 ;
        POLYGON 155.455 43.585 155.545 43.585 155.455 43.570 ;
        POLYGON 157.045 43.585 157.045 43.570 157.000 43.570 ;
        RECT 157.045 43.570 158.355 43.585 ;
        POLYGON 154.220 43.570 154.255 43.570 154.255 43.565 ;
        RECT 154.255 43.565 155.305 43.570 ;
        RECT 151.225 43.540 152.820 43.565 ;
        RECT 117.295 43.520 151.065 43.540 ;
        POLYGON 151.225 43.540 151.235 43.540 151.235 43.535 ;
        RECT 151.235 43.535 152.820 43.540 ;
        POLYGON 151.065 43.535 151.075 43.520 151.065 43.520 ;
        RECT 117.295 43.495 151.075 43.520 ;
        POLYGON 151.235 43.535 151.285 43.535 151.285 43.510 ;
        RECT 151.285 43.530 152.820 43.535 ;
        POLYGON 152.820 43.565 152.930 43.530 152.820 43.530 ;
        POLYGON 154.255 43.565 154.345 43.565 154.345 43.555 ;
        RECT 154.345 43.555 155.305 43.565 ;
        POLYGON 154.345 43.555 154.430 43.555 154.430 43.545 ;
        RECT 154.430 43.550 155.305 43.555 ;
        POLYGON 155.305 43.570 155.455 43.570 155.305 43.550 ;
        POLYGON 157.000 43.570 157.000 43.550 156.940 43.550 ;
        RECT 157.000 43.550 158.355 43.570 ;
        RECT 154.430 43.545 155.250 43.550 ;
        POLYGON 155.250 43.550 155.300 43.550 155.250 43.545 ;
        POLYGON 156.940 43.550 156.940 43.545 156.930 43.545 ;
        RECT 156.940 43.545 158.355 43.550 ;
        POLYGON 154.430 43.545 154.510 43.545 154.510 43.540 ;
        RECT 154.510 43.540 155.045 43.545 ;
        POLYGON 154.515 43.540 154.565 43.540 154.565 43.535 ;
        RECT 154.565 43.535 155.045 43.540 ;
        POLYGON 154.565 43.535 154.640 43.535 154.640 43.530 ;
        RECT 154.640 43.530 155.045 43.535 ;
        POLYGON 155.045 43.545 155.250 43.545 155.045 43.530 ;
        POLYGON 156.930 43.545 156.930 43.540 156.915 43.540 ;
        RECT 156.930 43.540 158.355 43.545 ;
        POLYGON 156.915 43.540 156.915 43.535 156.890 43.535 ;
        RECT 156.915 43.535 158.355 43.540 ;
        POLYGON 156.890 43.535 156.890 43.530 156.875 43.530 ;
        RECT 156.890 43.530 158.355 43.535 ;
        POLYGON 158.355 43.610 158.505 43.610 158.355 43.530 ;
        POLYGON 159.760 43.610 159.760 43.580 159.720 43.580 ;
        RECT 159.760 43.600 160.860 43.610 ;
        POLYGON 160.860 43.710 160.975 43.710 160.860 43.600 ;
        POLYGON 162.255 43.710 162.255 43.660 162.210 43.660 ;
        RECT 162.255 43.660 163.735 43.715 ;
        POLYGON 162.210 43.660 162.210 43.610 162.170 43.610 ;
        RECT 162.210 43.610 163.735 43.660 ;
        POLYGON 162.170 43.610 162.170 43.600 162.160 43.600 ;
        RECT 162.170 43.600 163.735 43.610 ;
        RECT 159.760 43.580 160.835 43.600 ;
        POLYGON 160.835 43.600 160.860 43.600 160.835 43.580 ;
        POLYGON 162.160 43.600 162.160 43.580 162.145 43.580 ;
        RECT 162.160 43.580 163.735 43.600 ;
        POLYGON 159.720 43.580 159.720 43.545 159.680 43.545 ;
        RECT 159.720 43.545 160.615 43.580 ;
        POLYGON 159.680 43.545 159.680 43.530 159.660 43.530 ;
        RECT 159.680 43.530 160.615 43.545 ;
        RECT 151.285 43.520 152.930 43.530 ;
        POLYGON 152.930 43.530 152.970 43.520 152.930 43.520 ;
        POLYGON 154.640 43.530 154.765 43.530 154.765 43.525 ;
        RECT 154.765 43.525 154.845 43.530 ;
        POLYGON 154.845 43.530 155.005 43.530 154.845 43.525 ;
        POLYGON 156.875 43.530 156.875 43.525 156.860 43.525 ;
        RECT 156.875 43.525 158.235 43.530 ;
        POLYGON 156.860 43.525 156.860 43.520 156.840 43.520 ;
        RECT 156.860 43.520 158.235 43.525 ;
        RECT 151.285 43.510 152.970 43.520 ;
        POLYGON 151.075 43.510 151.085 43.495 151.075 43.495 ;
        RECT 117.295 43.445 151.085 43.495 ;
        POLYGON 151.285 43.510 151.320 43.510 151.320 43.490 ;
        RECT 151.320 43.490 152.970 43.510 ;
        POLYGON 151.085 43.490 151.110 43.445 151.085 43.445 ;
        RECT 117.295 43.390 151.110 43.445 ;
        POLYGON 151.320 43.490 151.410 43.490 151.410 43.440 ;
        RECT 151.410 43.485 152.970 43.490 ;
        POLYGON 152.970 43.520 153.085 43.485 152.970 43.485 ;
        POLYGON 156.840 43.520 156.840 43.490 156.745 43.490 ;
        RECT 156.840 43.490 158.235 43.520 ;
        POLYGON 156.745 43.490 156.745 43.485 156.725 43.485 ;
        RECT 156.745 43.485 158.235 43.490 ;
        RECT 151.410 43.480 153.090 43.485 ;
        POLYGON 153.090 43.485 153.100 43.480 153.090 43.480 ;
        POLYGON 156.725 43.485 156.725 43.480 156.710 43.480 ;
        RECT 156.725 43.480 158.235 43.485 ;
        RECT 151.410 43.470 153.100 43.480 ;
        POLYGON 153.100 43.480 153.145 43.470 153.100 43.470 ;
        POLYGON 156.710 43.480 156.710 43.470 156.685 43.470 ;
        RECT 156.710 43.470 158.235 43.480 ;
        RECT 151.410 43.450 153.145 43.470 ;
        POLYGON 153.145 43.470 153.225 43.450 153.145 43.450 ;
        POLYGON 156.685 43.470 156.685 43.460 156.655 43.460 ;
        RECT 156.685 43.465 158.235 43.470 ;
        POLYGON 158.235 43.530 158.355 43.530 158.235 43.465 ;
        POLYGON 159.660 43.530 159.660 43.465 159.580 43.465 ;
        RECT 159.660 43.465 160.615 43.530 ;
        RECT 156.685 43.460 158.130 43.465 ;
        POLYGON 156.655 43.460 156.655 43.455 156.625 43.455 ;
        RECT 156.655 43.455 158.130 43.460 ;
        POLYGON 156.625 43.455 156.625 43.450 156.605 43.450 ;
        RECT 156.625 43.450 158.130 43.455 ;
        RECT 151.410 43.440 153.225 43.450 ;
        POLYGON 151.110 43.440 151.135 43.390 151.110 43.390 ;
        POLYGON 151.410 43.440 151.465 43.440 151.465 43.410 ;
        RECT 151.465 43.415 153.225 43.440 ;
        POLYGON 153.225 43.450 153.360 43.415 153.225 43.415 ;
        POLYGON 156.605 43.450 156.605 43.425 156.515 43.425 ;
        RECT 156.605 43.425 158.130 43.450 ;
        POLYGON 156.510 43.425 156.510 43.415 156.475 43.415 ;
        RECT 156.510 43.415 158.130 43.425 ;
        RECT 151.465 43.410 153.365 43.415 ;
        POLYGON 153.365 43.415 153.375 43.410 153.365 43.410 ;
        POLYGON 156.475 43.415 156.475 43.410 156.455 43.410 ;
        RECT 156.475 43.410 158.130 43.415 ;
        POLYGON 158.130 43.465 158.235 43.465 158.130 43.410 ;
        POLYGON 159.580 43.465 159.580 43.410 159.510 43.410 ;
        RECT 159.580 43.410 160.615 43.465 ;
        POLYGON 151.465 43.410 151.485 43.410 151.485 43.400 ;
        RECT 151.485 43.400 153.375 43.410 ;
        RECT 117.295 43.275 151.135 43.390 ;
        POLYGON 151.485 43.400 151.510 43.400 151.510 43.385 ;
        RECT 151.510 43.390 153.375 43.400 ;
        POLYGON 153.375 43.410 153.480 43.390 153.375 43.390 ;
        POLYGON 156.450 43.410 156.450 43.395 156.390 43.395 ;
        RECT 156.450 43.395 157.960 43.410 ;
        POLYGON 156.390 43.395 156.390 43.390 156.375 43.390 ;
        RECT 156.390 43.390 157.960 43.395 ;
        RECT 151.510 43.385 153.480 43.390 ;
        POLYGON 153.480 43.390 153.495 43.385 153.480 43.385 ;
        POLYGON 156.375 43.390 156.375 43.385 156.360 43.385 ;
        RECT 156.375 43.385 157.960 43.390 ;
        POLYGON 151.135 43.385 151.190 43.275 151.135 43.275 ;
        POLYGON 151.510 43.385 151.610 43.385 151.610 43.335 ;
        RECT 151.610 43.365 153.495 43.385 ;
        POLYGON 153.495 43.385 153.575 43.365 153.495 43.365 ;
        POLYGON 156.360 43.385 156.360 43.375 156.295 43.375 ;
        RECT 156.360 43.375 157.960 43.385 ;
        POLYGON 156.295 43.375 156.295 43.365 156.250 43.365 ;
        RECT 156.295 43.365 157.960 43.375 ;
        RECT 151.610 43.340 153.580 43.365 ;
        POLYGON 153.580 43.365 153.705 43.340 153.580 43.340 ;
        POLYGON 156.250 43.365 156.250 43.345 156.155 43.345 ;
        RECT 156.250 43.345 157.960 43.365 ;
        POLYGON 156.155 43.345 156.155 43.340 156.125 43.340 ;
        RECT 156.155 43.340 157.960 43.345 ;
        RECT 151.610 43.335 153.705 43.340 ;
        POLYGON 151.610 43.335 151.675 43.335 151.675 43.305 ;
        RECT 151.675 43.325 153.705 43.335 ;
        POLYGON 153.705 43.340 153.795 43.325 153.705 43.325 ;
        POLYGON 156.125 43.340 156.125 43.335 156.095 43.335 ;
        RECT 156.125 43.335 157.960 43.340 ;
        POLYGON 156.095 43.335 156.095 43.330 156.085 43.330 ;
        RECT 156.095 43.330 157.960 43.335 ;
        POLYGON 156.085 43.330 156.085 43.325 156.055 43.325 ;
        RECT 156.085 43.325 157.960 43.330 ;
        POLYGON 157.960 43.410 158.130 43.410 157.960 43.325 ;
        POLYGON 159.510 43.410 159.510 43.400 159.495 43.400 ;
        RECT 159.510 43.400 160.615 43.410 ;
        POLYGON 159.495 43.400 159.495 43.325 159.400 43.325 ;
        RECT 159.495 43.370 160.615 43.400 ;
        POLYGON 160.615 43.580 160.835 43.580 160.615 43.370 ;
        POLYGON 162.145 43.580 162.145 43.485 162.065 43.485 ;
        RECT 162.145 43.515 163.735 43.580 ;
        POLYGON 163.735 43.830 163.940 43.830 163.735 43.515 ;
        POLYGON 165.645 43.830 165.645 43.560 165.500 43.560 ;
        RECT 165.645 43.705 167.950 43.835 ;
        POLYGON 167.950 43.940 168.050 43.940 167.950 43.705 ;
        POLYGON 171.045 43.940 171.045 43.765 170.995 43.765 ;
        RECT 171.045 43.765 175.530 43.940 ;
        POLYGON 170.995 43.765 170.995 43.705 170.975 43.705 ;
        RECT 170.995 43.705 175.530 43.765 ;
        RECT 165.645 43.560 167.845 43.705 ;
        POLYGON 165.500 43.560 165.500 43.535 165.485 43.535 ;
        RECT 165.500 43.535 167.845 43.560 ;
        POLYGON 165.485 43.535 165.485 43.520 165.475 43.520 ;
        RECT 165.485 43.520 167.845 43.535 ;
        RECT 162.145 43.485 163.685 43.515 ;
        POLYGON 162.065 43.485 162.065 43.435 162.025 43.435 ;
        RECT 162.065 43.445 163.685 43.485 ;
        POLYGON 163.685 43.515 163.735 43.515 163.685 43.445 ;
        POLYGON 165.475 43.515 165.475 43.465 165.445 43.465 ;
        RECT 165.475 43.465 167.845 43.520 ;
        POLYGON 165.445 43.465 165.445 43.445 165.435 43.445 ;
        RECT 165.445 43.460 167.845 43.465 ;
        POLYGON 167.845 43.705 167.950 43.705 167.845 43.460 ;
        POLYGON 170.975 43.705 170.975 43.465 170.895 43.465 ;
        RECT 170.975 43.695 175.530 43.705 ;
        POLYGON 175.530 44.045 175.575 44.045 175.530 43.695 ;
        POLYGON 182.790 44.025 182.790 43.785 182.765 43.785 ;
        RECT 182.790 43.785 198.035 44.045 ;
        POLYGON 182.765 43.785 182.765 43.695 182.755 43.695 ;
        RECT 182.765 43.695 198.035 43.785 ;
        RECT 170.975 43.465 175.470 43.695 ;
        RECT 165.445 43.445 167.620 43.460 ;
        RECT 162.065 43.435 163.440 43.445 ;
        POLYGON 162.025 43.435 162.025 43.370 161.965 43.370 ;
        RECT 162.025 43.370 163.440 43.435 ;
        RECT 159.495 43.325 160.495 43.370 ;
        RECT 151.675 43.305 153.795 43.325 ;
        POLYGON 153.795 43.325 153.910 43.305 153.795 43.305 ;
        POLYGON 156.055 43.325 156.055 43.305 155.935 43.305 ;
        RECT 156.055 43.305 157.880 43.325 ;
        POLYGON 151.675 43.305 151.730 43.305 151.730 43.275 ;
        RECT 151.730 43.295 153.935 43.305 ;
        POLYGON 153.935 43.305 153.990 43.295 153.935 43.295 ;
        POLYGON 155.935 43.305 155.935 43.295 155.875 43.295 ;
        RECT 155.935 43.295 157.880 43.305 ;
        RECT 151.730 43.280 154.005 43.295 ;
        POLYGON 154.005 43.295 154.130 43.280 154.005 43.280 ;
        POLYGON 155.855 43.295 155.855 43.290 155.850 43.290 ;
        RECT 155.855 43.290 157.880 43.295 ;
        POLYGON 157.880 43.325 157.960 43.325 157.880 43.290 ;
        POLYGON 159.400 43.325 159.400 43.310 159.380 43.310 ;
        RECT 159.400 43.310 160.495 43.325 ;
        POLYGON 159.375 43.310 159.375 43.290 159.345 43.290 ;
        RECT 159.375 43.290 160.495 43.310 ;
        POLYGON 155.825 43.290 155.825 43.280 155.745 43.280 ;
        RECT 155.825 43.280 157.700 43.290 ;
        RECT 151.730 43.275 154.130 43.280 ;
        RECT 117.295 43.190 151.190 43.275 ;
        POLYGON 151.190 43.275 151.230 43.190 151.190 43.190 ;
        POLYGON 151.730 43.275 151.910 43.275 151.910 43.190 ;
        RECT 151.910 43.265 154.130 43.275 ;
        POLYGON 154.130 43.280 154.215 43.265 154.130 43.265 ;
        POLYGON 155.745 43.280 155.745 43.270 155.660 43.270 ;
        RECT 155.745 43.270 157.700 43.280 ;
        POLYGON 155.660 43.270 155.660 43.265 155.625 43.265 ;
        RECT 155.660 43.265 157.700 43.270 ;
        RECT 151.910 43.255 154.255 43.265 ;
        POLYGON 154.255 43.265 154.345 43.255 154.255 43.255 ;
        POLYGON 155.625 43.265 155.625 43.260 155.585 43.260 ;
        RECT 155.625 43.260 157.700 43.265 ;
        POLYGON 155.560 43.260 155.560 43.255 155.550 43.255 ;
        RECT 155.560 43.255 157.700 43.260 ;
        RECT 151.910 43.250 154.345 43.255 ;
        POLYGON 154.345 43.255 154.425 43.250 154.345 43.250 ;
        POLYGON 155.545 43.255 155.545 43.250 155.455 43.250 ;
        RECT 155.545 43.250 157.700 43.255 ;
        RECT 151.910 43.240 154.430 43.250 ;
        POLYGON 154.430 43.250 154.490 43.240 154.430 43.240 ;
        POLYGON 155.450 43.250 155.450 43.240 155.315 43.240 ;
        RECT 155.450 43.240 157.700 43.250 ;
        RECT 151.910 43.235 154.565 43.240 ;
        POLYGON 154.565 43.240 154.630 43.235 154.565 43.235 ;
        POLYGON 155.315 43.240 155.315 43.235 155.300 43.235 ;
        RECT 155.315 43.235 157.700 43.240 ;
        RECT 151.910 43.230 154.640 43.235 ;
        POLYGON 154.640 43.235 154.765 43.230 154.640 43.230 ;
        POLYGON 155.250 43.235 155.250 43.230 155.045 43.230 ;
        RECT 155.250 43.230 157.700 43.235 ;
        RECT 151.910 43.210 157.700 43.230 ;
        POLYGON 157.700 43.290 157.880 43.290 157.700 43.210 ;
        POLYGON 159.345 43.290 159.345 43.250 159.290 43.250 ;
        RECT 159.345 43.270 160.495 43.290 ;
        POLYGON 160.495 43.370 160.615 43.370 160.495 43.270 ;
        POLYGON 161.965 43.370 161.965 43.305 161.905 43.305 ;
        RECT 161.965 43.305 163.440 43.370 ;
        POLYGON 161.905 43.305 161.905 43.285 161.890 43.285 ;
        RECT 161.905 43.285 163.440 43.305 ;
        POLYGON 161.890 43.285 161.890 43.270 161.875 43.270 ;
        RECT 161.890 43.270 163.440 43.285 ;
        RECT 159.345 43.250 160.390 43.270 ;
        POLYGON 159.290 43.250 159.290 43.210 159.230 43.210 ;
        RECT 159.290 43.210 160.390 43.250 ;
        RECT 151.910 43.205 157.690 43.210 ;
        POLYGON 157.690 43.210 157.700 43.210 157.690 43.205 ;
        POLYGON 159.230 43.210 159.230 43.205 159.225 43.205 ;
        RECT 159.230 43.205 160.390 43.210 ;
        RECT 151.910 43.190 157.425 43.205 ;
        RECT 117.295 43.165 151.230 43.190 ;
        POLYGON 151.910 43.190 151.915 43.190 151.915 43.185 ;
        RECT 151.915 43.185 157.425 43.190 ;
        POLYGON 151.230 43.185 151.240 43.165 151.230 43.165 ;
        RECT 117.295 43.145 151.240 43.165 ;
        POLYGON 151.920 43.185 151.975 43.185 151.975 43.160 ;
        RECT 151.975 43.160 157.425 43.185 ;
        POLYGON 151.240 43.160 151.250 43.145 151.240 43.145 ;
        POLYGON 151.985 43.160 152.015 43.160 152.015 43.145 ;
        RECT 152.015 43.145 157.425 43.160 ;
        RECT 56.700 43.135 113.750 43.145 ;
        POLYGON 113.750 43.145 113.755 43.135 113.750 43.135 ;
        RECT 117.295 43.135 151.250 43.145 ;
        RECT 56.700 42.000 113.755 43.135 ;
        RECT 13.610 39.610 22.195 42.000 ;
        POLYGON 13.610 39.610 14.030 39.610 14.030 34.580 ;
        RECT 14.030 35.585 22.195 39.610 ;
        POLYGON 22.195 42.000 22.645 35.585 22.195 35.585 ;
        POLYGON 56.700 42.000 56.720 42.000 56.720 41.965 ;
        RECT 56.720 41.965 113.755 42.000 ;
        POLYGON 56.720 41.965 57.225 41.965 57.225 40.885 ;
        RECT 57.225 40.885 113.755 41.965 ;
        POLYGON 57.225 40.885 58.745 40.885 58.745 38.055 ;
        RECT 58.745 40.530 113.755 40.885 ;
        POLYGON 113.755 43.135 114.780 40.530 113.755 40.530 ;
        POLYGON 117.295 43.135 117.300 43.135 117.300 43.075 ;
        RECT 117.300 43.125 151.250 43.135 ;
        POLYGON 151.250 43.145 151.260 43.125 151.250 43.125 ;
        RECT 117.300 43.100 151.260 43.125 ;
        POLYGON 152.015 43.145 152.075 43.145 152.075 43.120 ;
        RECT 152.075 43.120 157.425 43.145 ;
        POLYGON 151.260 43.120 151.270 43.100 151.260 43.100 ;
        RECT 117.300 43.060 151.270 43.100 ;
        POLYGON 152.075 43.120 152.130 43.120 152.130 43.095 ;
        RECT 152.130 43.100 157.425 43.120 ;
        POLYGON 157.425 43.205 157.690 43.205 157.425 43.100 ;
        POLYGON 159.225 43.205 159.225 43.100 159.070 43.100 ;
        RECT 159.225 43.180 160.390 43.205 ;
        POLYGON 160.390 43.270 160.495 43.270 160.390 43.180 ;
        POLYGON 161.875 43.270 161.875 43.180 161.795 43.180 ;
        RECT 161.875 43.180 163.440 43.270 ;
        RECT 159.225 43.100 160.185 43.180 ;
        RECT 152.130 43.095 157.395 43.100 ;
        POLYGON 151.270 43.095 151.290 43.060 151.270 43.060 ;
        RECT 117.300 42.990 151.290 43.060 ;
        POLYGON 152.130 43.095 152.220 43.095 152.220 43.055 ;
        RECT 152.220 43.085 157.395 43.095 ;
        POLYGON 157.395 43.100 157.425 43.100 157.395 43.085 ;
        POLYGON 159.070 43.100 159.070 43.085 159.045 43.085 ;
        RECT 159.070 43.085 160.185 43.100 ;
        RECT 152.220 43.055 157.265 43.085 ;
        POLYGON 117.300 42.990 117.315 42.990 117.315 42.275 ;
        RECT 117.315 42.975 151.290 42.990 ;
        POLYGON 151.290 43.055 151.330 42.975 151.290 42.975 ;
        POLYGON 152.220 43.055 152.430 43.055 152.430 42.975 ;
        RECT 152.430 43.040 157.265 43.055 ;
        POLYGON 157.265 43.085 157.395 43.085 157.265 43.040 ;
        POLYGON 159.045 43.085 159.045 43.065 159.015 43.065 ;
        RECT 159.045 43.065 160.185 43.085 ;
        POLYGON 159.015 43.065 159.015 43.040 158.980 43.040 ;
        RECT 159.015 43.040 160.185 43.065 ;
        RECT 152.430 43.000 157.160 43.040 ;
        POLYGON 157.160 43.040 157.265 43.040 157.160 43.000 ;
        POLYGON 158.980 43.040 158.980 43.035 158.970 43.035 ;
        RECT 158.980 43.035 160.185 43.040 ;
        POLYGON 158.965 43.035 158.965 43.000 158.905 43.000 ;
        RECT 158.965 43.005 160.185 43.035 ;
        POLYGON 160.185 43.180 160.390 43.180 160.185 43.005 ;
        POLYGON 161.795 43.180 161.795 43.085 161.705 43.085 ;
        RECT 161.795 43.110 163.440 43.180 ;
        POLYGON 163.440 43.445 163.685 43.445 163.440 43.110 ;
        POLYGON 165.435 43.445 165.435 43.420 165.420 43.420 ;
        RECT 165.435 43.420 167.620 43.445 ;
        POLYGON 165.420 43.420 165.420 43.360 165.385 43.360 ;
        RECT 165.420 43.360 167.620 43.420 ;
        POLYGON 165.385 43.360 165.385 43.220 165.300 43.220 ;
        RECT 165.385 43.220 167.620 43.360 ;
        POLYGON 165.300 43.220 165.300 43.115 165.235 43.115 ;
        RECT 165.300 43.115 167.620 43.220 ;
        RECT 161.795 43.085 163.350 43.110 ;
        POLYGON 161.705 43.085 161.705 43.005 161.625 43.005 ;
        RECT 161.705 43.005 163.350 43.085 ;
        RECT 158.965 43.000 160.130 43.005 ;
        RECT 152.430 42.975 156.890 43.000 ;
        RECT 117.315 42.965 151.330 42.975 ;
        POLYGON 152.430 42.975 152.445 42.975 152.445 42.970 ;
        RECT 152.445 42.970 156.890 42.975 ;
        POLYGON 151.330 42.970 151.335 42.965 151.330 42.965 ;
        POLYGON 152.445 42.970 152.460 42.970 152.460 42.965 ;
        RECT 152.460 42.965 156.890 42.970 ;
        RECT 117.315 42.930 151.335 42.965 ;
        POLYGON 152.470 42.965 152.480 42.965 152.480 42.960 ;
        RECT 152.480 42.960 156.890 42.965 ;
        POLYGON 151.335 42.960 151.350 42.930 151.335 42.930 ;
        RECT 117.315 42.910 151.350 42.930 ;
        POLYGON 152.485 42.960 152.585 42.960 152.585 42.925 ;
        RECT 152.585 42.925 156.890 42.960 ;
        POLYGON 151.350 42.925 151.360 42.910 151.350 42.910 ;
        RECT 117.315 42.880 151.360 42.910 ;
        POLYGON 152.585 42.925 152.645 42.925 152.645 42.905 ;
        RECT 152.645 42.910 156.890 42.925 ;
        POLYGON 156.890 43.000 157.160 43.000 156.890 42.910 ;
        POLYGON 158.905 43.000 158.905 42.950 158.825 42.950 ;
        RECT 158.905 42.960 160.130 43.000 ;
        POLYGON 160.130 43.005 160.185 43.005 160.130 42.960 ;
        POLYGON 161.625 43.005 161.625 42.960 161.580 42.960 ;
        RECT 161.625 42.995 163.350 43.005 ;
        POLYGON 163.350 43.110 163.440 43.110 163.350 42.995 ;
        POLYGON 165.235 43.110 165.235 43.040 165.190 43.040 ;
        RECT 165.235 43.040 167.620 43.115 ;
        POLYGON 165.190 43.040 165.190 42.995 165.160 42.995 ;
        RECT 165.190 42.995 167.620 43.040 ;
        RECT 161.625 42.960 163.285 42.995 ;
        RECT 158.905 42.950 159.930 42.960 ;
        POLYGON 158.825 42.950 158.825 42.910 158.765 42.910 ;
        RECT 158.825 42.910 159.930 42.950 ;
        RECT 152.645 42.905 156.830 42.910 ;
        POLYGON 151.360 42.905 151.375 42.880 151.360 42.880 ;
        POLYGON 152.645 42.905 152.720 42.905 152.720 42.880 ;
        RECT 152.720 42.895 156.830 42.905 ;
        POLYGON 156.830 42.910 156.890 42.910 156.830 42.895 ;
        POLYGON 158.765 42.910 158.765 42.895 158.735 42.895 ;
        RECT 158.765 42.895 159.930 42.910 ;
        RECT 152.720 42.880 156.625 42.895 ;
        RECT 117.315 42.825 151.375 42.880 ;
        POLYGON 151.375 42.880 151.400 42.825 151.375 42.825 ;
        POLYGON 152.720 42.880 152.900 42.880 152.900 42.825 ;
        RECT 152.900 42.835 156.625 42.880 ;
        POLYGON 156.625 42.895 156.830 42.895 156.625 42.835 ;
        POLYGON 158.735 42.895 158.735 42.835 158.630 42.835 ;
        RECT 158.735 42.835 159.930 42.895 ;
        RECT 152.900 42.825 156.415 42.835 ;
        RECT 117.315 42.815 151.400 42.825 ;
        POLYGON 151.400 42.825 151.405 42.815 151.400 42.815 ;
        POLYGON 152.900 42.825 152.945 42.825 152.945 42.815 ;
        RECT 152.945 42.815 156.415 42.825 ;
        RECT 117.315 42.805 151.405 42.815 ;
        POLYGON 152.945 42.815 152.955 42.815 152.955 42.810 ;
        RECT 152.955 42.810 156.415 42.815 ;
        POLYGON 151.405 42.810 151.410 42.805 151.405 42.805 ;
        POLYGON 152.955 42.810 152.970 42.810 152.970 42.805 ;
        RECT 152.970 42.805 156.415 42.810 ;
        RECT 117.315 42.785 151.410 42.805 ;
        POLYGON 151.410 42.805 151.420 42.785 151.410 42.785 ;
        POLYGON 152.970 42.805 153.045 42.805 153.045 42.785 ;
        RECT 153.045 42.785 156.415 42.805 ;
        RECT 117.315 42.740 151.420 42.785 ;
        POLYGON 151.420 42.785 151.440 42.740 151.420 42.740 ;
        POLYGON 153.045 42.785 153.225 42.785 153.225 42.740 ;
        RECT 153.225 42.780 156.415 42.785 ;
        POLYGON 156.415 42.835 156.625 42.835 156.415 42.780 ;
        POLYGON 158.630 42.835 158.630 42.790 158.550 42.790 ;
        RECT 158.630 42.810 159.930 42.835 ;
        POLYGON 159.930 42.960 160.130 42.960 159.930 42.810 ;
        POLYGON 161.580 42.960 161.580 42.810 161.430 42.810 ;
        RECT 161.580 42.920 163.285 42.960 ;
        POLYGON 163.285 42.995 163.350 42.995 163.285 42.920 ;
        POLYGON 165.160 42.990 165.160 42.960 165.140 42.960 ;
        RECT 165.160 42.985 167.620 42.995 ;
        POLYGON 167.620 43.460 167.845 43.460 167.620 42.985 ;
        POLYGON 170.895 43.460 170.895 43.055 170.760 43.055 ;
        RECT 170.895 43.365 175.470 43.465 ;
        POLYGON 175.470 43.695 175.530 43.695 175.470 43.365 ;
        POLYGON 182.755 43.690 182.755 43.365 182.720 43.365 ;
        RECT 182.755 43.365 198.035 43.695 ;
        RECT 170.895 43.055 175.400 43.365 ;
        POLYGON 170.760 43.055 170.760 43.030 170.750 43.030 ;
        RECT 170.760 43.045 175.400 43.055 ;
        POLYGON 175.400 43.365 175.470 43.365 175.400 43.045 ;
        POLYGON 182.720 43.355 182.720 43.070 182.690 43.070 ;
        RECT 182.720 43.070 198.035 43.365 ;
        RECT 170.760 43.030 175.360 43.045 ;
        POLYGON 170.750 43.030 170.750 42.990 170.735 42.990 ;
        RECT 170.750 42.990 175.360 43.030 ;
        RECT 165.160 42.960 167.375 42.985 ;
        POLYGON 165.140 42.960 165.140 42.940 165.130 42.940 ;
        RECT 165.140 42.940 167.375 42.960 ;
        POLYGON 165.130 42.940 165.130 42.935 165.125 42.935 ;
        RECT 165.130 42.935 167.375 42.940 ;
        POLYGON 165.125 42.935 165.125 42.920 165.115 42.920 ;
        RECT 165.125 42.920 167.375 42.935 ;
        RECT 161.580 42.810 163.125 42.920 ;
        RECT 158.630 42.790 159.755 42.810 ;
        POLYGON 158.550 42.790 158.550 42.780 158.530 42.780 ;
        RECT 158.550 42.780 159.755 42.790 ;
        RECT 153.225 42.770 156.390 42.780 ;
        POLYGON 156.390 42.780 156.415 42.780 156.390 42.770 ;
        POLYGON 158.530 42.780 158.530 42.770 158.515 42.770 ;
        RECT 158.530 42.770 159.755 42.780 ;
        RECT 153.225 42.765 156.360 42.770 ;
        POLYGON 156.360 42.770 156.385 42.770 156.360 42.765 ;
        POLYGON 158.515 42.770 158.515 42.765 158.505 42.765 ;
        RECT 158.515 42.765 159.755 42.770 ;
        RECT 153.225 42.740 156.095 42.765 ;
        RECT 117.315 42.725 151.440 42.740 ;
        POLYGON 151.440 42.740 151.445 42.725 151.440 42.725 ;
        RECT 117.315 42.715 151.445 42.725 ;
        POLYGON 153.225 42.740 153.320 42.740 153.320 42.720 ;
        RECT 153.320 42.720 156.095 42.740 ;
        POLYGON 151.445 42.720 151.450 42.715 151.445 42.715 ;
        RECT 117.315 42.705 151.450 42.715 ;
        POLYGON 153.325 42.720 153.380 42.720 153.380 42.710 ;
        RECT 153.380 42.710 156.095 42.720 ;
        POLYGON 151.450 42.710 151.455 42.705 151.450 42.705 ;
        POLYGON 153.380 42.710 153.405 42.710 153.405 42.705 ;
        RECT 153.405 42.705 156.095 42.710 ;
        POLYGON 156.095 42.765 156.360 42.765 156.095 42.705 ;
        POLYGON 158.505 42.765 158.505 42.705 158.385 42.705 ;
        RECT 158.505 42.705 159.755 42.765 ;
        RECT 117.315 42.695 151.460 42.705 ;
        POLYGON 151.460 42.705 151.485 42.695 151.460 42.695 ;
        POLYGON 153.405 42.705 153.435 42.705 153.435 42.700 ;
        RECT 153.435 42.700 155.950 42.705 ;
        POLYGON 153.435 42.700 153.455 42.700 153.455 42.695 ;
        RECT 153.455 42.695 155.950 42.700 ;
        RECT 117.315 42.680 151.485 42.695 ;
        POLYGON 151.485 42.695 151.510 42.680 151.485 42.680 ;
        POLYGON 153.455 42.695 153.480 42.695 153.480 42.690 ;
        RECT 153.480 42.690 155.950 42.695 ;
        POLYGON 153.480 42.690 153.535 42.690 153.535 42.680 ;
        RECT 153.535 42.680 155.950 42.690 ;
        POLYGON 155.950 42.705 156.095 42.705 155.950 42.680 ;
        POLYGON 158.385 42.705 158.385 42.680 158.335 42.680 ;
        RECT 158.385 42.680 159.755 42.705 ;
        RECT 117.315 42.660 151.510 42.680 ;
        POLYGON 151.510 42.680 151.560 42.660 151.510 42.660 ;
        POLYGON 153.535 42.680 153.650 42.680 153.650 42.660 ;
        RECT 153.650 42.675 155.920 42.680 ;
        POLYGON 155.920 42.680 155.945 42.680 155.920 42.675 ;
        POLYGON 158.335 42.680 158.335 42.675 158.320 42.675 ;
        RECT 158.335 42.675 159.755 42.680 ;
        POLYGON 159.755 42.810 159.930 42.810 159.755 42.675 ;
        POLYGON 161.430 42.810 161.430 42.710 161.330 42.710 ;
        RECT 161.430 42.715 163.125 42.810 ;
        POLYGON 163.125 42.920 163.285 42.920 163.125 42.715 ;
        POLYGON 165.115 42.920 165.115 42.880 165.090 42.880 ;
        RECT 165.115 42.880 167.375 42.920 ;
        POLYGON 165.090 42.880 165.090 42.830 165.055 42.830 ;
        RECT 165.090 42.830 167.375 42.880 ;
        POLYGON 165.055 42.830 165.055 42.715 164.980 42.715 ;
        RECT 165.055 42.715 167.375 42.830 ;
        RECT 161.430 42.710 162.880 42.715 ;
        POLYGON 161.330 42.710 161.330 42.690 161.305 42.690 ;
        RECT 161.330 42.690 162.880 42.710 ;
        POLYGON 161.305 42.690 161.305 42.675 161.290 42.675 ;
        RECT 161.305 42.675 162.880 42.690 ;
        RECT 153.650 42.660 155.830 42.675 ;
        POLYGON 155.830 42.675 155.915 42.675 155.830 42.660 ;
        POLYGON 158.320 42.675 158.320 42.660 158.290 42.660 ;
        RECT 158.320 42.670 159.740 42.675 ;
        POLYGON 159.740 42.675 159.750 42.675 159.740 42.670 ;
        POLYGON 161.290 42.675 161.290 42.670 161.285 42.670 ;
        RECT 161.290 42.670 162.880 42.675 ;
        RECT 158.320 42.660 159.515 42.670 ;
        RECT 117.315 42.610 151.560 42.660 ;
        POLYGON 151.560 42.660 151.675 42.610 151.560 42.610 ;
        POLYGON 153.650 42.660 153.735 42.660 153.735 42.645 ;
        RECT 153.735 42.645 155.565 42.660 ;
        POLYGON 153.750 42.645 153.925 42.645 153.925 42.620 ;
        RECT 153.925 42.620 155.565 42.645 ;
        POLYGON 155.565 42.660 155.830 42.660 155.565 42.620 ;
        POLYGON 158.290 42.660 158.290 42.635 158.235 42.635 ;
        RECT 158.290 42.635 159.515 42.660 ;
        POLYGON 158.235 42.635 158.235 42.620 158.205 42.620 ;
        RECT 158.235 42.620 159.515 42.635 ;
        POLYGON 153.930 42.620 153.995 42.620 153.995 42.610 ;
        RECT 153.995 42.615 155.505 42.620 ;
        POLYGON 155.505 42.620 155.565 42.620 155.505 42.615 ;
        POLYGON 158.205 42.620 158.205 42.615 158.195 42.615 ;
        RECT 158.205 42.615 159.515 42.620 ;
        RECT 153.995 42.610 155.420 42.615 ;
        RECT 117.315 42.590 151.675 42.610 ;
        POLYGON 151.675 42.610 151.730 42.590 151.675 42.590 ;
        POLYGON 153.995 42.610 154.180 42.610 154.180 42.595 ;
        RECT 154.180 42.605 155.420 42.610 ;
        POLYGON 155.420 42.615 155.505 42.615 155.420 42.605 ;
        POLYGON 158.195 42.615 158.195 42.605 158.180 42.605 ;
        RECT 158.195 42.605 159.515 42.615 ;
        RECT 154.180 42.595 155.300 42.605 ;
        POLYGON 155.300 42.605 155.415 42.605 155.300 42.595 ;
        POLYGON 158.180 42.605 158.180 42.595 158.160 42.595 ;
        RECT 158.180 42.595 159.515 42.605 ;
        POLYGON 154.185 42.595 154.220 42.595 154.220 42.590 ;
        RECT 154.220 42.590 155.070 42.595 ;
        RECT 117.315 42.520 151.730 42.590 ;
        POLYGON 151.730 42.590 151.890 42.520 151.730 42.520 ;
        POLYGON 154.220 42.590 154.255 42.590 154.255 42.585 ;
        RECT 154.255 42.585 155.070 42.590 ;
        POLYGON 154.255 42.585 154.415 42.585 154.415 42.580 ;
        RECT 154.415 42.580 155.070 42.585 ;
        POLYGON 155.070 42.595 155.300 42.595 155.070 42.580 ;
        POLYGON 158.160 42.595 158.160 42.580 158.130 42.580 ;
        RECT 158.160 42.580 159.515 42.595 ;
        POLYGON 154.425 42.580 154.515 42.580 154.515 42.575 ;
        RECT 154.515 42.575 154.925 42.580 ;
        POLYGON 154.925 42.580 155.035 42.580 154.925 42.575 ;
        POLYGON 158.130 42.580 158.130 42.575 158.120 42.575 ;
        RECT 158.130 42.575 159.515 42.580 ;
        POLYGON 154.625 42.575 154.775 42.575 154.775 42.570 ;
        POLYGON 154.775 42.575 154.850 42.575 154.775 42.570 ;
        POLYGON 158.120 42.575 158.120 42.570 158.105 42.570 ;
        RECT 158.120 42.570 159.515 42.575 ;
        POLYGON 158.105 42.570 158.105 42.520 157.985 42.520 ;
        RECT 158.105 42.520 159.515 42.570 ;
        RECT 117.315 42.510 151.890 42.520 ;
        POLYGON 151.890 42.520 151.915 42.510 151.890 42.510 ;
        POLYGON 157.985 42.520 157.985 42.510 157.960 42.510 ;
        RECT 157.985 42.515 159.515 42.520 ;
        POLYGON 159.515 42.670 159.740 42.670 159.515 42.515 ;
        POLYGON 161.285 42.670 161.285 42.650 161.265 42.650 ;
        RECT 161.285 42.650 162.880 42.670 ;
        POLYGON 161.265 42.650 161.265 42.600 161.210 42.600 ;
        RECT 161.265 42.600 162.880 42.650 ;
        POLYGON 161.210 42.600 161.210 42.515 161.120 42.515 ;
        RECT 161.210 42.515 162.880 42.600 ;
        RECT 157.985 42.510 159.445 42.515 ;
        RECT 117.315 42.490 151.915 42.510 ;
        POLYGON 151.915 42.510 151.975 42.490 151.915 42.490 ;
        POLYGON 157.960 42.510 157.960 42.490 157.915 42.490 ;
        RECT 157.960 42.490 159.445 42.510 ;
        RECT 117.315 42.485 151.975 42.490 ;
        POLYGON 151.975 42.490 151.980 42.485 151.975 42.485 ;
        POLYGON 157.915 42.490 157.915 42.485 157.905 42.485 ;
        RECT 157.915 42.485 159.445 42.490 ;
        RECT 117.315 42.450 151.985 42.485 ;
        POLYGON 151.985 42.485 152.075 42.450 151.985 42.450 ;
        POLYGON 157.905 42.485 157.905 42.475 157.880 42.475 ;
        RECT 157.905 42.475 159.445 42.485 ;
        POLYGON 157.875 42.475 157.875 42.450 157.820 42.450 ;
        RECT 157.875 42.470 159.445 42.475 ;
        POLYGON 159.445 42.515 159.515 42.515 159.445 42.470 ;
        POLYGON 161.120 42.515 161.120 42.470 161.070 42.470 ;
        RECT 161.120 42.470 162.880 42.515 ;
        RECT 157.875 42.450 159.290 42.470 ;
        RECT 117.315 42.400 152.075 42.450 ;
        POLYGON 152.075 42.450 152.220 42.400 152.075 42.400 ;
        POLYGON 157.820 42.450 157.820 42.430 157.775 42.430 ;
        RECT 157.820 42.430 159.290 42.450 ;
        POLYGON 157.775 42.430 157.775 42.405 157.700 42.405 ;
        RECT 157.775 42.405 159.290 42.430 ;
        POLYGON 157.700 42.405 157.700 42.400 157.695 42.400 ;
        RECT 157.700 42.400 159.290 42.405 ;
        RECT 117.315 42.395 152.220 42.400 ;
        POLYGON 152.220 42.400 152.225 42.395 152.220 42.395 ;
        POLYGON 157.690 42.400 157.690 42.395 157.675 42.395 ;
        RECT 157.690 42.395 159.290 42.400 ;
        RECT 117.315 42.320 152.225 42.395 ;
        POLYGON 152.225 42.395 152.460 42.320 152.225 42.320 ;
        POLYGON 157.675 42.395 157.675 42.320 157.470 42.320 ;
        RECT 157.675 42.365 159.290 42.395 ;
        POLYGON 159.290 42.470 159.445 42.470 159.290 42.365 ;
        POLYGON 161.070 42.470 161.070 42.380 160.975 42.380 ;
        RECT 161.070 42.440 162.880 42.470 ;
        POLYGON 162.880 42.715 163.125 42.715 162.880 42.440 ;
        POLYGON 164.980 42.715 164.980 42.595 164.895 42.595 ;
        RECT 164.980 42.595 167.375 42.715 ;
        POLYGON 164.895 42.595 164.895 42.480 164.820 42.480 ;
        RECT 164.895 42.515 167.375 42.595 ;
        POLYGON 167.375 42.985 167.620 42.985 167.375 42.515 ;
        POLYGON 170.735 42.985 170.735 42.520 170.555 42.520 ;
        RECT 170.735 42.895 175.360 42.990 ;
        POLYGON 175.360 43.045 175.400 43.045 175.360 42.895 ;
        POLYGON 182.690 43.045 182.690 42.895 182.670 42.895 ;
        RECT 182.690 42.895 198.035 43.070 ;
        RECT 170.735 42.725 175.315 42.895 ;
        POLYGON 175.315 42.895 175.360 42.895 175.315 42.725 ;
        POLYGON 182.670 42.880 182.670 42.830 182.665 42.830 ;
        RECT 182.670 42.830 198.035 42.895 ;
        POLYGON 182.665 42.830 182.665 42.725 182.650 42.725 ;
        RECT 182.665 42.725 198.035 42.830 ;
        RECT 170.735 42.520 175.235 42.725 ;
        RECT 164.895 42.480 167.135 42.515 ;
        POLYGON 164.820 42.480 164.820 42.445 164.795 42.445 ;
        RECT 164.820 42.445 167.135 42.480 ;
        POLYGON 164.795 42.445 164.795 42.440 164.790 42.440 ;
        RECT 164.795 42.440 167.135 42.445 ;
        RECT 161.070 42.380 162.790 42.440 ;
        POLYGON 160.975 42.380 160.975 42.365 160.955 42.365 ;
        RECT 160.975 42.365 162.790 42.380 ;
        RECT 157.675 42.355 159.275 42.365 ;
        POLYGON 159.275 42.365 159.290 42.365 159.275 42.355 ;
        POLYGON 160.955 42.365 160.955 42.355 160.945 42.355 ;
        RECT 160.955 42.355 162.790 42.365 ;
        RECT 157.675 42.320 159.025 42.355 ;
        RECT 117.315 42.315 152.460 42.320 ;
        POLYGON 152.460 42.320 152.470 42.315 152.460 42.315 ;
        POLYGON 157.470 42.320 157.470 42.315 157.455 42.315 ;
        RECT 157.470 42.315 159.025 42.320 ;
        RECT 117.315 42.285 152.485 42.315 ;
        POLYGON 152.485 42.315 152.560 42.285 152.485 42.285 ;
        POLYGON 157.455 42.315 157.455 42.285 157.365 42.285 ;
        RECT 157.455 42.285 159.025 42.315 ;
        RECT 117.315 42.245 152.560 42.285 ;
        POLYGON 152.560 42.285 152.720 42.245 152.560 42.245 ;
        POLYGON 157.365 42.285 157.365 42.255 157.265 42.255 ;
        RECT 157.365 42.255 159.025 42.285 ;
        POLYGON 157.265 42.255 157.265 42.245 157.235 42.245 ;
        RECT 157.265 42.245 159.025 42.255 ;
        RECT 117.315 42.190 152.720 42.245 ;
        POLYGON 152.720 42.245 152.895 42.190 152.720 42.190 ;
        POLYGON 157.235 42.245 157.235 42.220 157.160 42.220 ;
        RECT 157.235 42.220 159.025 42.245 ;
        POLYGON 157.155 42.220 157.155 42.190 157.045 42.190 ;
        RECT 157.155 42.210 159.025 42.220 ;
        POLYGON 159.025 42.355 159.275 42.355 159.025 42.210 ;
        POLYGON 160.945 42.355 160.945 42.285 160.860 42.285 ;
        RECT 160.945 42.340 162.790 42.355 ;
        POLYGON 162.790 42.440 162.880 42.440 162.790 42.340 ;
        POLYGON 164.790 42.440 164.790 42.340 164.720 42.340 ;
        RECT 164.790 42.340 167.135 42.440 ;
        RECT 160.945 42.290 162.740 42.340 ;
        POLYGON 162.740 42.340 162.790 42.340 162.740 42.290 ;
        POLYGON 164.720 42.340 164.720 42.320 164.705 42.320 ;
        RECT 164.720 42.320 167.135 42.340 ;
        POLYGON 164.705 42.320 164.705 42.290 164.685 42.290 ;
        RECT 164.705 42.290 167.135 42.320 ;
        RECT 160.945 42.285 162.460 42.290 ;
        POLYGON 160.860 42.285 160.860 42.265 160.835 42.265 ;
        RECT 160.860 42.265 162.460 42.285 ;
        POLYGON 160.835 42.265 160.835 42.210 160.770 42.210 ;
        RECT 160.835 42.210 162.460 42.265 ;
        RECT 157.155 42.190 158.825 42.210 ;
        RECT 117.315 42.180 152.905 42.190 ;
        POLYGON 152.905 42.190 152.945 42.180 152.905 42.180 ;
        POLYGON 157.045 42.190 157.045 42.180 157.005 42.180 ;
        RECT 157.045 42.180 158.825 42.190 ;
        RECT 117.315 42.175 152.945 42.180 ;
        POLYGON 152.945 42.180 152.970 42.175 152.945 42.175 ;
        POLYGON 157.005 42.180 157.005 42.175 156.985 42.175 ;
        RECT 157.005 42.175 158.825 42.180 ;
        RECT 117.315 42.145 152.970 42.175 ;
        POLYGON 117.315 42.145 117.320 42.145 117.320 42.010 ;
        RECT 117.320 42.115 152.970 42.145 ;
        POLYGON 152.970 42.175 153.225 42.115 152.970 42.115 ;
        POLYGON 156.985 42.175 156.985 42.155 156.910 42.155 ;
        RECT 156.985 42.155 158.825 42.175 ;
        POLYGON 156.905 42.155 156.905 42.150 156.890 42.150 ;
        RECT 156.905 42.150 158.825 42.155 ;
        POLYGON 156.890 42.150 156.890 42.135 156.830 42.135 ;
        RECT 156.890 42.135 158.825 42.150 ;
        POLYGON 156.825 42.135 156.825 42.115 156.755 42.115 ;
        RECT 156.825 42.115 158.825 42.135 ;
        RECT 117.320 42.110 153.225 42.115 ;
        POLYGON 153.225 42.115 153.250 42.110 153.225 42.110 ;
        POLYGON 156.755 42.115 156.755 42.110 156.735 42.110 ;
        RECT 156.755 42.110 158.825 42.115 ;
        RECT 117.320 42.095 153.250 42.110 ;
        POLYGON 153.250 42.110 153.320 42.095 153.250 42.095 ;
        POLYGON 156.735 42.110 156.735 42.095 156.670 42.095 ;
        RECT 156.735 42.095 158.825 42.110 ;
        POLYGON 158.825 42.210 159.025 42.210 158.825 42.095 ;
        POLYGON 160.770 42.210 160.770 42.095 160.635 42.095 ;
        RECT 160.770 42.095 162.460 42.210 ;
        RECT 117.320 42.070 153.325 42.095 ;
        POLYGON 153.325 42.095 153.435 42.070 153.325 42.070 ;
        POLYGON 156.670 42.095 156.670 42.085 156.625 42.085 ;
        RECT 156.670 42.085 158.785 42.095 ;
        POLYGON 156.625 42.085 156.625 42.070 156.545 42.070 ;
        RECT 156.625 42.070 158.785 42.085 ;
        POLYGON 158.785 42.095 158.825 42.095 158.785 42.070 ;
        POLYGON 160.635 42.095 160.635 42.080 160.615 42.080 ;
        RECT 160.635 42.080 162.460 42.095 ;
        POLYGON 160.615 42.080 160.615 42.070 160.605 42.070 ;
        RECT 160.615 42.070 162.460 42.080 ;
        RECT 117.320 42.065 153.435 42.070 ;
        POLYGON 153.435 42.070 153.480 42.065 153.435 42.065 ;
        POLYGON 156.545 42.070 156.545 42.065 156.520 42.065 ;
        RECT 156.545 42.065 158.770 42.070 ;
        POLYGON 158.770 42.070 158.780 42.070 158.770 42.065 ;
        POLYGON 160.605 42.070 160.605 42.065 160.595 42.065 ;
        RECT 160.605 42.065 162.460 42.070 ;
        RECT 117.320 42.040 153.480 42.065 ;
        POLYGON 153.480 42.065 153.595 42.040 153.480 42.040 ;
        POLYGON 156.520 42.065 156.520 42.045 156.415 42.045 ;
        RECT 156.520 42.045 158.355 42.065 ;
        POLYGON 156.415 42.045 156.415 42.040 156.410 42.040 ;
        RECT 156.415 42.040 158.355 42.045 ;
        RECT 117.320 42.020 153.595 42.040 ;
        POLYGON 153.595 42.040 153.735 42.020 153.595 42.020 ;
        POLYGON 156.385 42.040 156.385 42.035 156.360 42.035 ;
        RECT 156.385 42.035 158.355 42.040 ;
        POLYGON 156.355 42.035 156.355 42.020 156.270 42.020 ;
        RECT 156.355 42.020 158.355 42.035 ;
        RECT 117.320 42.015 153.735 42.020 ;
        POLYGON 153.735 42.020 153.750 42.015 153.735 42.015 ;
        POLYGON 156.270 42.020 156.270 42.015 156.240 42.015 ;
        RECT 156.270 42.015 158.355 42.020 ;
        RECT 117.320 42.010 153.750 42.015 ;
        POLYGON 117.320 42.010 117.335 42.010 117.335 41.795 ;
        RECT 117.335 41.990 153.750 42.010 ;
        POLYGON 153.750 42.015 153.930 41.990 153.750 41.990 ;
        POLYGON 156.240 42.015 156.240 41.990 156.095 41.990 ;
        RECT 156.240 41.990 158.355 42.015 ;
        RECT 117.335 41.985 153.930 41.990 ;
        POLYGON 153.930 41.990 153.945 41.985 153.930 41.985 ;
        POLYGON 156.090 41.990 156.090 41.985 156.060 41.985 ;
        RECT 156.090 41.985 158.355 41.990 ;
        RECT 117.335 41.980 153.945 41.985 ;
        POLYGON 153.945 41.985 153.995 41.980 153.945 41.980 ;
        POLYGON 156.060 41.985 156.060 41.980 156.005 41.980 ;
        RECT 156.060 41.980 158.355 41.985 ;
        RECT 117.335 41.960 153.995 41.980 ;
        POLYGON 153.995 41.980 154.180 41.960 153.995 41.960 ;
        POLYGON 156.005 41.980 156.005 41.975 155.945 41.975 ;
        RECT 156.005 41.975 158.355 41.980 ;
        POLYGON 155.945 41.975 155.945 41.970 155.920 41.970 ;
        RECT 155.945 41.970 158.355 41.975 ;
        POLYGON 155.915 41.970 155.915 41.960 155.830 41.960 ;
        RECT 155.915 41.960 158.355 41.970 ;
        RECT 117.335 41.955 154.185 41.960 ;
        POLYGON 154.185 41.960 154.250 41.955 154.185 41.955 ;
        POLYGON 155.830 41.960 155.830 41.955 155.790 41.955 ;
        RECT 155.830 41.955 158.355 41.960 ;
        RECT 117.335 41.950 154.255 41.955 ;
        POLYGON 154.255 41.955 154.300 41.950 154.255 41.950 ;
        POLYGON 155.790 41.955 155.790 41.950 155.750 41.950 ;
        RECT 155.790 41.950 158.355 41.955 ;
        RECT 117.335 41.940 154.300 41.950 ;
        POLYGON 154.300 41.950 154.415 41.940 154.300 41.940 ;
        POLYGON 155.750 41.950 155.750 41.945 155.710 41.945 ;
        RECT 155.750 41.945 158.355 41.950 ;
        POLYGON 155.710 41.945 155.710 41.940 155.570 41.940 ;
        RECT 155.710 41.940 158.355 41.945 ;
        RECT 117.335 41.935 154.425 41.940 ;
        POLYGON 154.425 41.940 154.505 41.935 154.425 41.935 ;
        POLYGON 155.565 41.940 155.565 41.935 155.510 41.935 ;
        RECT 155.565 41.935 158.355 41.940 ;
        RECT 117.335 41.925 154.515 41.935 ;
        POLYGON 154.515 41.935 154.620 41.925 154.515 41.925 ;
        POLYGON 155.505 41.935 155.505 41.930 155.420 41.930 ;
        RECT 155.505 41.930 158.355 41.935 ;
        POLYGON 155.415 41.930 155.415 41.925 155.355 41.925 ;
        RECT 155.415 41.925 158.355 41.930 ;
        RECT 117.335 41.920 154.650 41.925 ;
        POLYGON 154.650 41.925 154.825 41.920 154.650 41.920 ;
        POLYGON 155.300 41.925 155.300 41.920 155.065 41.920 ;
        RECT 155.300 41.920 158.355 41.925 ;
        RECT 117.335 41.915 154.925 41.920 ;
        POLYGON 154.925 41.920 155.005 41.915 154.925 41.915 ;
        POLYGON 155.035 41.920 155.035 41.915 155.005 41.915 ;
        RECT 155.035 41.915 158.355 41.920 ;
        RECT 117.335 41.855 158.355 41.915 ;
        POLYGON 158.355 42.065 158.770 42.065 158.355 41.855 ;
        POLYGON 160.595 42.065 160.595 42.040 160.565 42.040 ;
        RECT 160.595 42.040 162.460 42.065 ;
        POLYGON 160.565 42.040 160.565 41.985 160.500 41.985 ;
        RECT 160.565 42.000 162.460 42.040 ;
        POLYGON 162.460 42.290 162.740 42.290 162.460 42.000 ;
        POLYGON 164.685 42.290 164.685 42.065 164.520 42.065 ;
        RECT 164.685 42.095 167.135 42.290 ;
        POLYGON 167.135 42.515 167.375 42.515 167.135 42.095 ;
        POLYGON 170.555 42.515 170.555 42.360 170.495 42.360 ;
        RECT 170.555 42.460 175.235 42.520 ;
        POLYGON 175.235 42.725 175.315 42.725 175.235 42.460 ;
        POLYGON 182.650 42.725 182.650 42.520 182.620 42.520 ;
        RECT 182.650 42.520 198.035 42.725 ;
        POLYGON 182.620 42.520 182.620 42.460 182.610 42.460 ;
        RECT 182.620 42.460 198.035 42.520 ;
        RECT 170.555 42.360 175.110 42.460 ;
        POLYGON 170.495 42.355 170.495 42.350 170.490 42.350 ;
        RECT 170.495 42.350 175.110 42.360 ;
        POLYGON 170.490 42.350 170.490 42.265 170.455 42.265 ;
        RECT 170.490 42.265 175.110 42.350 ;
        POLYGON 170.455 42.265 170.455 42.095 170.380 42.095 ;
        RECT 170.455 42.095 175.110 42.265 ;
        RECT 164.685 42.065 167.110 42.095 ;
        POLYGON 164.520 42.065 164.520 42.030 164.495 42.030 ;
        RECT 164.520 42.050 167.110 42.065 ;
        POLYGON 167.110 42.095 167.135 42.095 167.110 42.050 ;
        POLYGON 170.380 42.095 170.380 42.050 170.360 42.050 ;
        RECT 170.380 42.060 175.110 42.095 ;
        POLYGON 175.110 42.460 175.235 42.460 175.110 42.060 ;
        POLYGON 182.610 42.450 182.610 42.070 182.555 42.070 ;
        RECT 182.610 42.070 198.035 42.460 ;
        RECT 170.380 42.050 174.845 42.060 ;
        RECT 164.520 42.030 167.020 42.050 ;
        POLYGON 164.495 42.030 164.495 42.000 164.470 42.000 ;
        RECT 164.495 42.000 167.020 42.030 ;
        RECT 160.565 41.985 162.440 42.000 ;
        POLYGON 160.495 41.985 160.495 41.905 160.390 41.905 ;
        RECT 160.495 41.980 162.440 41.985 ;
        POLYGON 162.440 42.000 162.460 42.000 162.440 41.980 ;
        POLYGON 164.470 42.000 164.470 41.980 164.450 41.980 ;
        RECT 164.470 41.980 167.020 42.000 ;
        RECT 160.495 41.905 162.120 41.980 ;
        POLYGON 160.390 41.905 160.390 41.855 160.325 41.855 ;
        RECT 160.390 41.855 162.120 41.905 ;
        RECT 117.335 41.800 158.240 41.855 ;
        POLYGON 158.240 41.855 158.355 41.855 158.240 41.800 ;
        POLYGON 160.325 41.855 160.325 41.800 160.255 41.800 ;
        RECT 160.325 41.800 162.120 41.855 ;
        RECT 117.335 41.790 158.210 41.800 ;
        POLYGON 158.210 41.800 158.240 41.800 158.210 41.790 ;
        POLYGON 160.255 41.800 160.255 41.790 160.245 41.790 ;
        RECT 160.255 41.790 162.120 41.800 ;
        RECT 117.335 41.760 157.950 41.790 ;
        POLYGON 117.335 41.760 117.365 41.760 117.365 41.375 ;
        RECT 117.365 41.675 157.950 41.760 ;
        POLYGON 157.950 41.790 158.210 41.790 157.950 41.675 ;
        POLYGON 160.245 41.790 160.245 41.745 160.185 41.745 ;
        RECT 160.245 41.745 162.120 41.790 ;
        POLYGON 160.180 41.745 160.180 41.675 160.080 41.675 ;
        RECT 160.180 41.685 162.120 41.745 ;
        POLYGON 162.120 41.980 162.440 41.980 162.120 41.685 ;
        POLYGON 164.450 41.980 164.450 41.960 164.435 41.960 ;
        RECT 164.450 41.960 167.020 41.980 ;
        POLYGON 164.435 41.960 164.435 41.740 164.260 41.740 ;
        RECT 164.435 41.910 167.020 41.960 ;
        POLYGON 167.020 42.050 167.110 42.050 167.020 41.910 ;
        POLYGON 170.360 42.045 170.360 41.910 170.300 41.910 ;
        RECT 170.360 41.910 174.845 42.050 ;
        RECT 164.435 41.740 166.825 41.910 ;
        POLYGON 164.260 41.740 164.260 41.685 164.215 41.685 ;
        RECT 164.260 41.685 166.825 41.740 ;
        RECT 160.180 41.675 162.065 41.685 ;
        RECT 117.365 41.645 157.880 41.675 ;
        POLYGON 157.880 41.675 157.945 41.675 157.880 41.645 ;
        POLYGON 160.080 41.675 160.080 41.645 160.035 41.645 ;
        RECT 160.080 41.645 162.065 41.675 ;
        RECT 117.365 41.575 157.695 41.645 ;
        POLYGON 157.695 41.645 157.880 41.645 157.695 41.575 ;
        POLYGON 160.035 41.645 160.035 41.575 159.935 41.575 ;
        RECT 160.035 41.635 162.065 41.645 ;
        POLYGON 162.065 41.685 162.120 41.685 162.065 41.635 ;
        POLYGON 164.215 41.685 164.215 41.640 164.180 41.640 ;
        RECT 164.215 41.640 166.825 41.685 ;
        RECT 160.035 41.600 162.025 41.635 ;
        POLYGON 162.025 41.635 162.065 41.635 162.025 41.600 ;
        POLYGON 164.180 41.635 164.180 41.600 164.150 41.600 ;
        RECT 164.180 41.600 166.825 41.640 ;
        RECT 160.035 41.575 161.675 41.600 ;
        RECT 117.365 41.480 157.440 41.575 ;
        POLYGON 157.440 41.575 157.695 41.575 157.440 41.480 ;
        POLYGON 159.935 41.575 159.935 41.570 159.930 41.570 ;
        RECT 159.935 41.570 161.675 41.575 ;
        POLYGON 159.930 41.570 159.930 41.480 159.790 41.480 ;
        RECT 159.930 41.480 161.675 41.570 ;
        RECT 117.365 41.465 157.395 41.480 ;
        POLYGON 157.395 41.480 157.440 41.480 157.395 41.465 ;
        POLYGON 159.790 41.480 159.790 41.465 159.765 41.465 ;
        RECT 159.790 41.465 161.675 41.480 ;
        RECT 117.365 41.415 157.190 41.465 ;
        RECT 117.365 41.410 152.070 41.415 ;
        POLYGON 152.070 41.415 152.075 41.410 152.070 41.410 ;
        POLYGON 152.075 41.415 152.085 41.415 152.085 41.410 ;
        RECT 152.085 41.410 157.190 41.415 ;
        RECT 117.365 41.395 152.075 41.410 ;
        POLYGON 152.075 41.410 152.085 41.395 152.075 41.395 ;
        POLYGON 152.085 41.410 152.130 41.410 152.130 41.395 ;
        RECT 152.130 41.400 157.190 41.410 ;
        POLYGON 157.190 41.465 157.395 41.465 157.190 41.400 ;
        POLYGON 159.765 41.465 159.765 41.455 159.750 41.455 ;
        RECT 159.765 41.455 161.675 41.465 ;
        POLYGON 159.750 41.455 159.750 41.450 159.740 41.450 ;
        RECT 159.750 41.450 161.675 41.455 ;
        POLYGON 159.740 41.450 159.740 41.400 159.660 41.400 ;
        RECT 159.740 41.400 161.675 41.450 ;
        RECT 152.130 41.395 157.140 41.400 ;
        RECT 117.365 41.375 152.085 41.395 ;
        POLYGON 152.130 41.395 152.150 41.395 152.150 41.390 ;
        RECT 152.150 41.390 157.140 41.395 ;
        POLYGON 152.085 41.390 152.095 41.375 152.085 41.375 ;
        POLYGON 152.150 41.390 152.200 41.390 152.200 41.375 ;
        RECT 152.200 41.385 157.140 41.390 ;
        POLYGON 157.140 41.400 157.190 41.400 157.140 41.385 ;
        POLYGON 159.660 41.400 159.660 41.385 159.635 41.385 ;
        RECT 159.660 41.385 161.675 41.400 ;
        RECT 152.200 41.375 156.930 41.385 ;
        RECT 117.365 41.320 152.095 41.375 ;
        POLYGON 152.095 41.375 152.125 41.320 152.095 41.320 ;
        RECT 117.365 41.310 152.125 41.320 ;
        POLYGON 152.200 41.375 152.405 41.375 152.405 41.315 ;
        RECT 152.405 41.320 156.930 41.375 ;
        POLYGON 156.930 41.385 157.140 41.385 156.930 41.320 ;
        POLYGON 159.635 41.385 159.635 41.320 159.530 41.320 ;
        RECT 159.635 41.320 161.675 41.385 ;
        RECT 152.405 41.315 156.905 41.320 ;
        POLYGON 156.905 41.320 156.930 41.320 156.905 41.315 ;
        POLYGON 159.530 41.320 159.530 41.315 159.525 41.315 ;
        RECT 159.530 41.315 161.675 41.320 ;
        POLYGON 117.365 41.310 117.400 41.310 117.400 40.880 ;
        RECT 117.400 41.300 152.125 41.310 ;
        POLYGON 152.125 41.315 152.135 41.300 152.125 41.300 ;
        POLYGON 152.405 41.315 152.460 41.315 152.460 41.300 ;
        RECT 152.460 41.300 156.660 41.315 ;
        RECT 117.400 41.280 152.135 41.300 ;
        POLYGON 152.135 41.300 152.145 41.280 152.135 41.280 ;
        RECT 117.400 41.260 152.145 41.280 ;
        POLYGON 152.470 41.300 152.570 41.300 152.570 41.275 ;
        RECT 152.570 41.275 156.660 41.300 ;
        POLYGON 152.145 41.275 152.155 41.260 152.145 41.260 ;
        RECT 117.400 41.250 152.155 41.260 ;
        POLYGON 152.570 41.275 152.655 41.275 152.655 41.255 ;
        RECT 152.655 41.255 156.660 41.275 ;
        POLYGON 156.660 41.315 156.905 41.315 156.660 41.255 ;
        POLYGON 159.525 41.315 159.525 41.310 159.515 41.310 ;
        RECT 159.525 41.310 161.675 41.315 ;
        POLYGON 159.515 41.310 159.515 41.270 159.445 41.270 ;
        RECT 159.515 41.300 161.675 41.310 ;
        POLYGON 161.675 41.600 162.025 41.600 161.675 41.300 ;
        POLYGON 164.150 41.600 164.150 41.505 164.065 41.505 ;
        RECT 164.150 41.590 166.825 41.600 ;
        POLYGON 166.825 41.910 167.020 41.910 166.825 41.590 ;
        POLYGON 170.300 41.910 170.300 41.680 170.200 41.680 ;
        RECT 170.300 41.680 174.845 41.910 ;
        POLYGON 170.200 41.680 170.200 41.665 170.195 41.665 ;
        RECT 170.200 41.665 174.845 41.680 ;
        POLYGON 170.195 41.665 170.195 41.595 170.160 41.595 ;
        RECT 170.195 41.595 174.845 41.665 ;
        RECT 164.150 41.505 166.595 41.590 ;
        POLYGON 164.065 41.505 164.065 41.440 164.010 41.440 ;
        RECT 164.065 41.440 166.595 41.505 ;
        POLYGON 164.010 41.440 164.010 41.360 163.940 41.360 ;
        RECT 164.010 41.360 166.595 41.440 ;
        POLYGON 163.940 41.360 163.940 41.300 163.885 41.300 ;
        RECT 163.940 41.300 166.595 41.360 ;
        RECT 159.515 41.270 161.585 41.300 ;
        POLYGON 159.445 41.270 159.445 41.255 159.420 41.255 ;
        RECT 159.445 41.255 161.585 41.270 ;
        POLYGON 152.155 41.255 152.160 41.250 152.155 41.250 ;
        POLYGON 152.655 41.255 152.670 41.255 152.670 41.250 ;
        RECT 152.670 41.250 156.570 41.255 ;
        RECT 117.400 41.200 152.160 41.250 ;
        POLYGON 152.160 41.250 152.185 41.200 152.160 41.200 ;
        POLYGON 152.670 41.250 152.750 41.250 152.750 41.230 ;
        RECT 152.750 41.235 156.570 41.250 ;
        POLYGON 156.570 41.255 156.660 41.255 156.570 41.235 ;
        POLYGON 159.420 41.255 159.420 41.240 159.395 41.240 ;
        RECT 159.420 41.240 161.585 41.255 ;
        POLYGON 159.395 41.240 159.395 41.235 159.385 41.235 ;
        RECT 159.395 41.235 161.585 41.240 ;
        RECT 152.750 41.230 156.415 41.235 ;
        RECT 117.400 41.190 152.185 41.200 ;
        POLYGON 152.750 41.230 152.895 41.230 152.895 41.195 ;
        RECT 152.895 41.195 156.415 41.230 ;
        POLYGON 156.415 41.235 156.570 41.235 156.415 41.195 ;
        POLYGON 159.385 41.235 159.385 41.195 159.310 41.195 ;
        RECT 159.385 41.230 161.585 41.235 ;
        POLYGON 161.585 41.300 161.675 41.300 161.585 41.230 ;
        POLYGON 163.885 41.300 163.885 41.230 163.825 41.230 ;
        RECT 163.885 41.245 166.595 41.300 ;
        POLYGON 166.595 41.590 166.825 41.590 166.595 41.245 ;
        POLYGON 170.160 41.590 170.160 41.245 169.990 41.245 ;
        RECT 170.160 41.305 174.845 41.595 ;
        POLYGON 174.845 42.060 175.110 42.060 174.845 41.305 ;
        POLYGON 182.555 42.060 182.555 41.485 182.470 41.485 ;
        RECT 182.555 41.790 198.035 42.070 ;
        POLYGON 198.035 44.095 198.075 41.790 198.035 41.790 ;
        POLYGON 208.495 44.095 208.800 44.095 208.800 43.155 ;
        RECT 208.800 43.860 223.450 44.095 ;
        POLYGON 223.450 44.095 223.530 43.860 223.450 43.860 ;
        POLYGON 230.515 44.095 230.545 44.095 230.545 44.005 ;
        RECT 230.545 44.005 234.745 44.095 ;
        POLYGON 230.545 44.005 230.600 44.005 230.600 43.865 ;
        RECT 230.600 43.940 234.745 44.005 ;
        POLYGON 234.745 44.095 234.820 43.940 234.745 43.940 ;
        POLYGON 237.685 44.095 237.715 44.095 237.715 44.045 ;
        RECT 237.715 44.045 239.855 44.095 ;
        POLYGON 237.715 44.045 237.765 44.045 237.765 43.945 ;
        RECT 237.765 43.945 239.855 44.045 ;
        POLYGON 239.855 44.095 239.955 43.945 239.855 43.945 ;
        POLYGON 241.605 44.095 241.670 44.095 241.670 44.015 ;
        RECT 241.670 44.055 243.070 44.095 ;
        POLYGON 243.070 44.095 243.110 44.055 243.070 44.055 ;
        POLYGON 244.310 44.095 244.340 44.095 244.340 44.070 ;
        RECT 244.340 44.085 245.425 44.095 ;
        POLYGON 245.425 44.095 245.440 44.085 245.425 44.085 ;
        POLYGON 246.585 44.095 246.605 44.095 246.605 44.085 ;
        RECT 246.605 44.085 247.555 44.095 ;
        RECT 244.340 44.080 245.440 44.085 ;
        POLYGON 245.440 44.085 245.445 44.080 245.440 44.080 ;
        POLYGON 246.605 44.085 246.615 44.085 246.615 44.080 ;
        RECT 246.615 44.080 247.555 44.085 ;
        POLYGON 247.555 44.110 247.615 44.080 247.555 44.080 ;
        POLYGON 252.145 44.110 252.145 44.095 252.115 44.095 ;
        RECT 252.145 44.095 253.145 44.110 ;
        POLYGON 253.145 44.110 253.170 44.110 253.145 44.095 ;
        POLYGON 254.255 44.110 254.255 44.095 254.235 44.095 ;
        RECT 254.255 44.095 255.295 44.110 ;
        POLYGON 255.295 44.260 255.455 44.260 255.295 44.095 ;
        POLYGON 256.465 44.260 256.465 44.190 256.410 44.190 ;
        RECT 256.465 44.195 257.615 44.260 ;
        POLYGON 257.615 44.460 257.795 44.460 257.615 44.195 ;
        POLYGON 259.310 44.460 259.310 44.425 259.290 44.425 ;
        RECT 259.310 44.435 260.945 44.465 ;
        POLYGON 260.945 44.600 261.025 44.600 260.945 44.435 ;
        POLYGON 263.310 44.600 263.310 44.555 263.295 44.555 ;
        RECT 263.310 44.595 266.210 44.605 ;
        POLYGON 266.210 44.670 266.230 44.670 266.210 44.600 ;
        POLYGON 270.610 44.670 270.610 44.625 270.605 44.625 ;
        RECT 270.610 44.625 277.820 44.710 ;
        RECT 270.605 44.600 277.820 44.625 ;
        POLYGON 277.820 45.630 277.885 45.630 277.820 44.610 ;
        POLYGON 287.860 45.630 287.860 44.610 287.805 44.610 ;
        RECT 287.860 44.610 303.120 45.650 ;
        RECT 263.310 44.555 266.080 44.595 ;
        POLYGON 263.295 44.555 263.295 44.435 263.250 44.435 ;
        RECT 263.295 44.435 266.080 44.555 ;
        RECT 259.310 44.425 260.780 44.435 ;
        POLYGON 259.290 44.425 259.290 44.370 259.265 44.370 ;
        RECT 259.290 44.370 260.780 44.425 ;
        POLYGON 259.265 44.370 259.265 44.330 259.240 44.330 ;
        RECT 259.265 44.330 260.780 44.370 ;
        POLYGON 259.240 44.330 259.240 44.220 259.175 44.220 ;
        RECT 259.240 44.220 260.780 44.330 ;
        POLYGON 259.175 44.220 259.175 44.195 259.160 44.195 ;
        RECT 259.175 44.195 260.780 44.220 ;
        RECT 256.465 44.190 257.595 44.195 ;
        POLYGON 256.410 44.190 256.410 44.145 256.375 44.145 ;
        RECT 256.410 44.175 257.595 44.190 ;
        POLYGON 257.595 44.195 257.615 44.195 257.595 44.175 ;
        POLYGON 259.160 44.195 259.160 44.180 259.150 44.180 ;
        RECT 259.160 44.180 260.780 44.195 ;
        POLYGON 259.150 44.180 259.150 44.175 259.145 44.175 ;
        RECT 259.150 44.175 260.780 44.180 ;
        RECT 256.410 44.145 257.535 44.175 ;
        POLYGON 256.375 44.145 256.375 44.095 256.330 44.095 ;
        RECT 256.375 44.095 257.535 44.145 ;
        POLYGON 257.535 44.175 257.595 44.175 257.535 44.095 ;
        POLYGON 259.145 44.170 259.145 44.105 259.105 44.105 ;
        RECT 259.145 44.105 260.780 44.175 ;
        POLYGON 259.105 44.100 259.105 44.095 259.100 44.095 ;
        RECT 259.105 44.095 260.780 44.105 ;
        POLYGON 260.780 44.435 260.945 44.435 260.780 44.100 ;
        POLYGON 263.250 44.430 263.250 44.330 263.215 44.330 ;
        RECT 263.250 44.330 266.080 44.435 ;
        POLYGON 263.215 44.330 263.215 44.140 263.145 44.140 ;
        RECT 263.215 44.140 266.080 44.330 ;
        POLYGON 263.145 44.140 263.145 44.100 263.130 44.100 ;
        RECT 263.145 44.100 266.080 44.140 ;
        POLYGON 266.080 44.595 266.210 44.595 266.080 44.105 ;
        POLYGON 270.605 44.600 270.605 44.135 270.575 44.135 ;
        RECT 270.605 44.215 277.795 44.600 ;
        POLYGON 277.795 44.600 277.820 44.600 277.795 44.215 ;
        POLYGON 287.805 44.600 287.805 44.215 287.785 44.215 ;
        RECT 287.805 44.215 303.120 44.610 ;
        RECT 270.605 44.135 277.780 44.215 ;
        RECT 263.130 44.095 266.080 44.100 ;
        POLYGON 252.115 44.095 252.115 44.080 252.080 44.080 ;
        RECT 252.115 44.080 253.085 44.095 ;
        RECT 244.340 44.070 245.445 44.080 ;
        POLYGON 244.340 44.070 244.355 44.070 244.355 44.055 ;
        RECT 244.355 44.055 245.445 44.070 ;
        RECT 241.670 44.015 243.110 44.055 ;
        POLYGON 241.670 44.015 241.720 44.015 241.720 43.950 ;
        RECT 241.720 43.945 243.110 44.015 ;
        RECT 237.765 43.940 239.955 43.945 ;
        RECT 230.600 43.860 234.820 43.940 ;
        RECT 208.800 43.625 223.530 43.860 ;
        POLYGON 223.530 43.860 223.620 43.625 223.530 43.625 ;
        POLYGON 230.600 43.860 230.695 43.860 230.695 43.630 ;
        RECT 230.695 43.625 234.820 43.860 ;
        RECT 208.800 43.155 223.620 43.625 ;
        POLYGON 208.800 43.155 208.805 43.155 208.805 43.145 ;
        RECT 208.805 43.145 223.620 43.155 ;
        RECT 182.555 41.485 198.000 41.790 ;
        POLYGON 182.470 41.485 182.470 41.305 182.435 41.305 ;
        RECT 182.470 41.305 198.000 41.485 ;
        RECT 170.160 41.245 174.425 41.305 ;
        RECT 163.885 41.230 166.515 41.245 ;
        RECT 159.385 41.195 161.485 41.230 ;
        POLYGON 152.185 41.195 152.190 41.190 152.185 41.190 ;
        RECT 117.400 41.170 152.190 41.190 ;
        POLYGON 152.895 41.195 152.945 41.195 152.945 41.185 ;
        RECT 152.945 41.190 156.375 41.195 ;
        POLYGON 156.375 41.195 156.415 41.195 156.375 41.190 ;
        POLYGON 159.310 41.195 159.310 41.190 159.300 41.190 ;
        RECT 159.310 41.190 161.485 41.195 ;
        RECT 152.945 41.185 156.065 41.190 ;
        POLYGON 152.190 41.185 152.200 41.170 152.190 41.170 ;
        RECT 117.400 41.145 152.200 41.170 ;
        POLYGON 152.945 41.185 153.050 41.185 153.050 41.165 ;
        RECT 153.050 41.165 156.065 41.185 ;
        POLYGON 152.200 41.165 152.215 41.145 152.200 41.145 ;
        POLYGON 153.055 41.165 153.180 41.165 153.180 41.145 ;
        RECT 153.180 41.145 156.065 41.165 ;
        RECT 117.400 41.105 152.215 41.145 ;
        POLYGON 152.215 41.145 152.235 41.105 152.215 41.105 ;
        RECT 117.400 41.085 152.235 41.105 ;
        POLYGON 153.180 41.145 153.435 41.145 153.435 41.100 ;
        RECT 153.435 41.130 156.065 41.145 ;
        POLYGON 156.065 41.190 156.375 41.190 156.065 41.130 ;
        POLYGON 159.300 41.190 159.300 41.185 159.290 41.185 ;
        RECT 159.300 41.185 161.485 41.190 ;
        POLYGON 159.290 41.185 159.290 41.175 159.275 41.175 ;
        RECT 159.290 41.175 161.485 41.185 ;
        POLYGON 159.275 41.175 159.275 41.130 159.190 41.130 ;
        RECT 159.275 41.155 161.485 41.175 ;
        POLYGON 161.485 41.230 161.585 41.230 161.485 41.155 ;
        POLYGON 163.825 41.230 163.825 41.185 163.785 41.185 ;
        RECT 163.825 41.185 166.515 41.230 ;
        POLYGON 163.785 41.185 163.785 41.160 163.760 41.160 ;
        RECT 163.785 41.160 166.515 41.185 ;
        RECT 159.275 41.130 161.265 41.155 ;
        RECT 153.435 41.120 155.995 41.130 ;
        POLYGON 155.995 41.130 156.065 41.130 155.995 41.120 ;
        POLYGON 159.190 41.130 159.190 41.120 159.170 41.120 ;
        RECT 159.190 41.120 161.265 41.130 ;
        RECT 153.435 41.105 155.920 41.120 ;
        POLYGON 155.920 41.120 155.995 41.120 155.920 41.105 ;
        POLYGON 159.170 41.120 159.170 41.105 159.140 41.105 ;
        RECT 159.170 41.105 161.265 41.120 ;
        RECT 153.435 41.100 155.420 41.105 ;
        POLYGON 152.235 41.100 152.245 41.085 152.235 41.085 ;
        POLYGON 153.435 41.100 153.555 41.100 153.555 41.085 ;
        RECT 153.555 41.085 155.420 41.100 ;
        RECT 117.400 41.065 152.245 41.085 ;
        POLYGON 153.555 41.085 153.600 41.085 153.600 41.080 ;
        RECT 153.600 41.080 155.420 41.085 ;
        POLYGON 152.245 41.080 152.255 41.065 152.245 41.065 ;
        POLYGON 153.600 41.080 153.725 41.080 153.725 41.065 ;
        RECT 153.725 41.065 155.420 41.080 ;
        RECT 117.400 41.035 152.255 41.065 ;
        POLYGON 152.255 41.065 152.270 41.035 152.255 41.035 ;
        POLYGON 153.735 41.065 153.930 41.065 153.930 41.045 ;
        RECT 153.930 41.045 155.420 41.065 ;
        POLYGON 155.420 41.105 155.920 41.105 155.420 41.045 ;
        POLYGON 159.140 41.105 159.140 41.045 159.025 41.045 ;
        RECT 159.140 41.045 161.265 41.105 ;
        RECT 117.400 41.025 152.270 41.035 ;
        POLYGON 153.930 41.045 154.180 41.045 154.180 41.030 ;
        RECT 154.180 41.030 154.925 41.045 ;
        POLYGON 152.270 41.030 152.275 41.025 152.270 41.025 ;
        POLYGON 154.180 41.030 154.265 41.030 154.265 41.025 ;
        RECT 154.265 41.025 154.925 41.030 ;
        RECT 117.400 41.015 152.275 41.025 ;
        POLYGON 152.275 41.025 152.280 41.015 152.275 41.015 ;
        POLYGON 154.280 41.025 154.425 41.025 154.425 41.015 ;
        RECT 154.425 41.015 154.925 41.025 ;
        POLYGON 154.925 41.045 155.370 41.045 154.925 41.015 ;
        POLYGON 159.020 41.045 159.020 41.025 158.985 41.025 ;
        RECT 159.020 41.025 161.265 41.045 ;
        POLYGON 158.985 41.025 158.985 41.015 158.965 41.015 ;
        RECT 158.985 41.015 161.265 41.025 ;
        RECT 117.400 40.950 152.280 41.015 ;
        POLYGON 152.280 41.015 152.315 40.950 152.280 40.950 ;
        POLYGON 158.965 41.015 158.965 40.950 158.830 40.950 ;
        RECT 158.965 40.985 161.265 41.015 ;
        POLYGON 161.265 41.155 161.485 41.155 161.265 40.985 ;
        POLYGON 163.760 41.155 163.760 41.130 163.735 41.130 ;
        RECT 163.760 41.135 166.515 41.160 ;
        POLYGON 166.515 41.245 166.595 41.245 166.515 41.135 ;
        POLYGON 169.990 41.240 169.990 41.140 169.940 41.140 ;
        RECT 169.990 41.140 174.425 41.245 ;
        RECT 163.760 41.130 166.190 41.135 ;
        POLYGON 163.735 41.130 163.735 41.075 163.685 41.075 ;
        RECT 163.735 41.075 166.190 41.130 ;
        POLYGON 163.685 41.075 163.685 40.985 163.600 40.985 ;
        RECT 163.685 40.985 166.190 41.075 ;
        RECT 158.965 40.950 161.130 40.985 ;
        RECT 117.400 40.870 152.315 40.950 ;
        POLYGON 152.315 40.950 152.355 40.870 152.315 40.870 ;
        POLYGON 158.825 40.950 158.825 40.930 158.785 40.930 ;
        RECT 158.825 40.930 161.130 40.950 ;
        POLYGON 158.780 40.930 158.780 40.920 158.760 40.920 ;
        RECT 158.780 40.920 161.130 40.930 ;
        POLYGON 158.760 40.920 158.760 40.910 158.735 40.910 ;
        RECT 158.760 40.910 161.130 40.920 ;
        POLYGON 117.400 40.870 117.420 40.870 117.420 40.600 ;
        RECT 117.420 40.840 152.355 40.870 ;
        POLYGON 158.735 40.910 158.735 40.865 158.635 40.865 ;
        RECT 158.735 40.890 161.130 40.910 ;
        POLYGON 161.130 40.985 161.265 40.985 161.130 40.890 ;
        POLYGON 163.600 40.985 163.600 40.890 163.505 40.890 ;
        RECT 163.600 40.890 166.190 40.985 ;
        RECT 158.735 40.865 160.835 40.890 ;
        POLYGON 152.355 40.865 152.370 40.840 152.355 40.840 ;
        RECT 117.420 40.765 152.370 40.840 ;
        POLYGON 158.635 40.865 158.635 40.835 158.570 40.835 ;
        RECT 158.635 40.835 160.835 40.865 ;
        POLYGON 152.370 40.835 152.410 40.765 152.370 40.765 ;
        POLYGON 158.570 40.835 158.570 40.765 158.395 40.765 ;
        RECT 158.570 40.765 160.835 40.835 ;
        RECT 117.420 40.755 152.410 40.765 ;
        POLYGON 152.410 40.765 152.415 40.755 152.410 40.755 ;
        RECT 117.420 40.745 152.415 40.755 ;
        POLYGON 158.395 40.765 158.395 40.750 158.360 40.750 ;
        RECT 158.395 40.750 160.835 40.765 ;
        POLYGON 152.415 40.750 152.420 40.745 152.415 40.745 ;
        POLYGON 158.355 40.750 158.355 40.745 158.340 40.745 ;
        RECT 158.355 40.745 160.835 40.750 ;
        RECT 117.420 40.675 152.420 40.745 ;
        POLYGON 152.420 40.745 152.455 40.675 152.420 40.675 ;
        POLYGON 158.340 40.745 158.340 40.705 158.240 40.705 ;
        RECT 158.340 40.705 160.835 40.745 ;
        POLYGON 158.240 40.705 158.240 40.695 158.210 40.695 ;
        RECT 158.240 40.695 160.835 40.705 ;
        RECT 117.420 40.665 152.455 40.675 ;
        POLYGON 158.210 40.695 158.210 40.670 158.140 40.670 ;
        RECT 158.210 40.685 160.835 40.695 ;
        POLYGON 160.835 40.890 161.130 40.890 160.835 40.685 ;
        POLYGON 163.505 40.890 163.505 40.820 163.440 40.820 ;
        RECT 163.505 40.820 166.190 40.890 ;
        POLYGON 163.440 40.820 163.440 40.730 163.350 40.730 ;
        RECT 163.440 40.730 166.190 40.820 ;
        POLYGON 163.350 40.730 163.350 40.685 163.300 40.685 ;
        RECT 163.350 40.685 166.190 40.730 ;
        POLYGON 166.190 41.135 166.515 41.135 166.190 40.685 ;
        POLYGON 169.940 41.135 169.940 41.025 169.885 41.025 ;
        RECT 169.940 41.025 174.425 41.140 ;
        POLYGON 169.885 41.025 169.885 40.990 169.865 40.990 ;
        RECT 169.885 40.990 174.425 41.025 ;
        POLYGON 169.865 40.990 169.865 40.685 169.700 40.685 ;
        RECT 169.865 40.685 174.425 40.990 ;
        RECT 158.210 40.670 160.665 40.685 ;
        POLYGON 152.455 40.670 152.460 40.665 152.455 40.665 ;
        POLYGON 158.140 40.670 158.140 40.665 158.125 40.665 ;
        RECT 158.140 40.665 160.665 40.670 ;
        RECT 117.420 40.595 152.460 40.665 ;
        POLYGON 152.460 40.665 152.495 40.595 152.460 40.595 ;
        POLYGON 158.125 40.665 158.125 40.605 157.950 40.605 ;
        RECT 158.125 40.605 160.665 40.665 ;
        RECT 117.420 40.535 152.495 40.595 ;
        POLYGON 157.945 40.605 157.945 40.590 157.895 40.590 ;
        RECT 157.945 40.590 160.665 40.605 ;
        POLYGON 117.420 40.535 117.425 40.535 117.425 40.530 ;
        RECT 117.425 40.530 152.495 40.535 ;
        POLYGON 152.495 40.590 152.530 40.530 152.495 40.530 ;
        RECT 58.745 40.410 114.780 40.530 ;
        POLYGON 114.780 40.530 114.835 40.410 114.780 40.410 ;
        RECT 117.425 40.510 152.530 40.530 ;
        POLYGON 157.895 40.590 157.895 40.525 157.700 40.525 ;
        RECT 157.895 40.575 160.665 40.590 ;
        POLYGON 160.665 40.685 160.830 40.685 160.665 40.575 ;
        POLYGON 163.300 40.685 163.300 40.670 163.285 40.670 ;
        RECT 163.300 40.670 166.070 40.685 ;
        POLYGON 163.285 40.670 163.285 40.575 163.185 40.575 ;
        RECT 163.285 40.575 166.070 40.670 ;
        RECT 157.895 40.525 160.390 40.575 ;
        POLYGON 152.530 40.525 152.540 40.510 152.530 40.510 ;
        RECT 117.425 40.500 152.540 40.510 ;
        POLYGON 157.690 40.525 157.690 40.505 157.615 40.505 ;
        RECT 157.690 40.505 160.390 40.525 ;
        POLYGON 152.540 40.505 152.545 40.500 152.540 40.500 ;
        POLYGON 157.615 40.505 157.615 40.500 157.595 40.500 ;
        RECT 157.615 40.500 160.390 40.505 ;
        RECT 117.425 40.495 152.545 40.500 ;
        POLYGON 117.425 40.495 117.430 40.495 117.430 40.460 ;
        RECT 117.430 40.490 152.545 40.495 ;
        POLYGON 152.545 40.500 152.550 40.490 152.545 40.490 ;
        RECT 117.430 40.480 152.550 40.490 ;
        POLYGON 157.595 40.500 157.595 40.485 157.540 40.485 ;
        RECT 157.595 40.485 160.390 40.500 ;
        POLYGON 152.550 40.485 152.555 40.480 152.550 40.480 ;
        RECT 117.430 40.460 152.555 40.480 ;
        POLYGON 157.540 40.485 157.540 40.475 157.500 40.475 ;
        RECT 157.540 40.475 160.390 40.485 ;
        POLYGON 152.555 40.475 152.565 40.460 152.555 40.460 ;
        POLYGON 157.500 40.475 157.500 40.460 157.445 40.460 ;
        RECT 157.500 40.460 160.390 40.475 ;
        RECT 117.430 40.430 152.565 40.460 ;
        POLYGON 152.565 40.460 152.580 40.430 152.565 40.430 ;
        POLYGON 157.440 40.460 157.440 40.450 157.395 40.450 ;
        RECT 157.440 40.450 160.390 40.460 ;
        POLYGON 157.395 40.450 157.395 40.430 157.320 40.430 ;
        RECT 157.395 40.430 160.390 40.450 ;
        RECT 117.430 40.410 152.580 40.430 ;
        POLYGON 157.320 40.430 157.320 40.425 157.300 40.425 ;
        RECT 157.320 40.425 160.390 40.430 ;
        POLYGON 152.580 40.425 152.590 40.410 152.580 40.410 ;
        POLYGON 157.300 40.425 157.300 40.410 157.245 40.410 ;
        RECT 157.300 40.410 160.390 40.425 ;
        RECT 58.745 39.260 114.835 40.410 ;
        POLYGON 114.835 40.410 115.350 39.260 114.835 39.260 ;
        POLYGON 117.430 40.410 117.460 40.410 117.460 40.035 ;
        RECT 117.460 40.400 152.590 40.410 ;
        POLYGON 152.590 40.410 152.595 40.400 152.590 40.400 ;
        POLYGON 157.245 40.410 157.245 40.400 157.210 40.400 ;
        RECT 157.245 40.405 160.390 40.410 ;
        POLYGON 160.390 40.575 160.660 40.575 160.390 40.405 ;
        POLYGON 163.185 40.575 163.185 40.515 163.125 40.515 ;
        RECT 163.185 40.530 166.070 40.575 ;
        POLYGON 166.070 40.685 166.190 40.685 166.070 40.530 ;
        POLYGON 169.700 40.685 169.700 40.665 169.690 40.665 ;
        RECT 169.700 40.665 174.425 40.685 ;
        POLYGON 169.690 40.665 169.690 40.530 169.615 40.530 ;
        RECT 169.690 40.530 174.425 40.665 ;
        RECT 163.185 40.515 166.050 40.530 ;
        POLYGON 163.125 40.515 163.125 40.405 163.010 40.405 ;
        RECT 163.125 40.505 166.050 40.515 ;
        POLYGON 166.050 40.530 166.070 40.530 166.050 40.505 ;
        POLYGON 169.615 40.530 169.615 40.510 169.605 40.510 ;
        RECT 169.615 40.510 174.425 40.530 ;
        RECT 163.125 40.405 165.845 40.505 ;
        RECT 157.245 40.400 160.185 40.405 ;
        RECT 117.460 40.385 152.595 40.400 ;
        POLYGON 157.210 40.400 157.210 40.395 157.190 40.395 ;
        RECT 157.210 40.395 160.185 40.400 ;
        POLYGON 152.595 40.395 152.605 40.385 152.595 40.385 ;
        POLYGON 157.190 40.395 157.190 40.385 157.140 40.385 ;
        RECT 157.190 40.385 160.185 40.395 ;
        RECT 117.460 40.345 152.605 40.385 ;
        POLYGON 152.605 40.385 152.625 40.345 152.605 40.345 ;
        POLYGON 157.140 40.385 157.140 40.345 156.930 40.345 ;
        RECT 157.140 40.345 160.185 40.385 ;
        RECT 117.460 40.315 152.625 40.345 ;
        POLYGON 156.930 40.345 156.930 40.340 156.905 40.340 ;
        RECT 156.930 40.340 160.185 40.345 ;
        POLYGON 152.625 40.340 152.640 40.315 152.625 40.315 ;
        RECT 117.460 40.305 152.640 40.315 ;
        POLYGON 156.905 40.340 156.905 40.310 156.770 40.310 ;
        RECT 156.905 40.310 160.185 40.340 ;
        POLYGON 152.640 40.310 152.645 40.305 152.640 40.305 ;
        POLYGON 156.770 40.310 156.770 40.305 156.735 40.305 ;
        RECT 156.770 40.305 160.185 40.310 ;
        RECT 117.460 40.285 152.645 40.305 ;
        POLYGON 152.645 40.305 152.655 40.285 152.645 40.285 ;
        POLYGON 156.735 40.305 156.735 40.295 156.660 40.295 ;
        RECT 156.735 40.295 160.185 40.305 ;
        RECT 117.460 40.255 152.655 40.285 ;
        POLYGON 156.660 40.295 156.660 40.280 156.570 40.280 ;
        RECT 156.660 40.285 160.185 40.295 ;
        POLYGON 160.185 40.405 160.390 40.405 160.185 40.285 ;
        POLYGON 163.010 40.405 163.010 40.290 162.880 40.290 ;
        RECT 163.010 40.290 165.845 40.405 ;
        POLYGON 162.880 40.290 162.880 40.285 162.875 40.285 ;
        RECT 162.880 40.285 165.845 40.290 ;
        RECT 156.660 40.280 160.160 40.285 ;
        POLYGON 152.655 40.280 152.670 40.255 152.655 40.255 ;
        POLYGON 156.570 40.280 156.570 40.255 156.415 40.255 ;
        RECT 156.570 40.270 160.160 40.280 ;
        POLYGON 160.160 40.285 160.185 40.285 160.160 40.270 ;
        POLYGON 162.875 40.285 162.875 40.270 162.855 40.270 ;
        RECT 162.875 40.270 165.845 40.285 ;
        RECT 156.570 40.255 159.930 40.270 ;
        RECT 117.460 40.245 152.670 40.255 ;
        POLYGON 156.415 40.255 156.415 40.250 156.375 40.250 ;
        RECT 156.415 40.250 159.930 40.255 ;
        POLYGON 152.670 40.250 152.675 40.245 152.670 40.245 ;
        POLYGON 156.375 40.250 156.375 40.245 156.345 40.245 ;
        RECT 156.375 40.245 159.930 40.250 ;
        RECT 117.460 40.225 152.675 40.245 ;
        POLYGON 152.675 40.245 152.685 40.225 152.675 40.225 ;
        POLYGON 156.345 40.245 156.345 40.235 156.280 40.235 ;
        RECT 156.345 40.235 159.930 40.245 ;
        RECT 117.460 40.215 152.685 40.225 ;
        POLYGON 156.280 40.235 156.280 40.220 156.120 40.220 ;
        RECT 156.280 40.220 159.930 40.235 ;
        POLYGON 152.685 40.220 152.690 40.215 152.685 40.215 ;
        POLYGON 156.120 40.220 156.120 40.215 156.065 40.215 ;
        RECT 156.120 40.215 159.930 40.220 ;
        RECT 117.460 40.210 152.690 40.215 ;
        POLYGON 152.690 40.215 152.730 40.210 152.690 40.210 ;
        POLYGON 156.065 40.215 156.065 40.210 156.030 40.210 ;
        RECT 156.065 40.210 159.930 40.215 ;
        RECT 117.460 40.205 152.730 40.210 ;
        POLYGON 152.730 40.210 152.750 40.205 152.730 40.205 ;
        POLYGON 156.030 40.210 156.030 40.205 155.995 40.205 ;
        RECT 156.030 40.205 159.930 40.210 ;
        RECT 117.460 40.190 152.750 40.205 ;
        POLYGON 152.750 40.205 152.895 40.190 152.750 40.190 ;
        POLYGON 155.995 40.205 155.995 40.200 155.920 40.200 ;
        RECT 155.995 40.200 159.930 40.205 ;
        POLYGON 155.920 40.200 155.920 40.190 155.820 40.190 ;
        RECT 155.920 40.190 159.930 40.200 ;
        RECT 117.460 40.185 152.895 40.190 ;
        POLYGON 152.895 40.190 152.940 40.185 152.895 40.185 ;
        POLYGON 155.820 40.190 155.820 40.185 155.770 40.185 ;
        RECT 155.820 40.185 159.930 40.190 ;
        RECT 117.460 40.175 152.945 40.185 ;
        POLYGON 152.945 40.185 153.055 40.175 152.945 40.175 ;
        POLYGON 155.770 40.185 155.770 40.175 155.630 40.175 ;
        RECT 155.770 40.175 159.930 40.185 ;
        RECT 117.460 40.170 153.055 40.175 ;
        POLYGON 153.055 40.175 153.175 40.170 153.055 40.170 ;
        POLYGON 155.630 40.175 155.630 40.170 155.560 40.170 ;
        RECT 155.630 40.170 159.930 40.175 ;
        RECT 117.460 40.160 153.180 40.170 ;
        POLYGON 153.180 40.170 153.285 40.160 153.180 40.160 ;
        POLYGON 155.560 40.170 155.560 40.160 155.420 40.160 ;
        RECT 155.560 40.160 159.930 40.170 ;
        RECT 117.460 40.155 153.285 40.160 ;
        POLYGON 153.285 40.160 153.405 40.155 153.285 40.155 ;
        POLYGON 155.370 40.160 155.370 40.155 155.305 40.155 ;
        RECT 155.370 40.155 159.930 40.160 ;
        RECT 117.460 40.145 153.435 40.155 ;
        POLYGON 153.435 40.155 153.715 40.145 153.435 40.145 ;
        POLYGON 155.305 40.155 155.305 40.150 155.240 40.150 ;
        RECT 155.305 40.150 159.930 40.155 ;
        POLYGON 155.240 40.150 155.240 40.145 155.085 40.145 ;
        RECT 155.240 40.145 159.930 40.150 ;
        RECT 117.460 40.140 153.735 40.145 ;
        POLYGON 153.735 40.145 153.925 40.140 153.735 40.140 ;
        POLYGON 155.085 40.145 155.085 40.140 154.925 40.140 ;
        RECT 155.085 40.140 159.930 40.145 ;
        POLYGON 159.930 40.270 160.160 40.270 159.930 40.140 ;
        POLYGON 162.855 40.270 162.855 40.215 162.790 40.215 ;
        RECT 162.855 40.245 165.845 40.270 ;
        POLYGON 165.845 40.505 166.050 40.505 165.845 40.245 ;
        POLYGON 169.605 40.505 169.605 40.390 169.540 40.390 ;
        RECT 169.605 40.390 174.425 40.510 ;
        POLYGON 169.540 40.390 169.540 40.325 169.505 40.325 ;
        RECT 169.540 40.325 174.425 40.390 ;
        POLYGON 169.505 40.325 169.505 40.245 169.455 40.245 ;
        RECT 169.505 40.245 174.425 40.325 ;
        RECT 162.855 40.215 165.575 40.245 ;
        POLYGON 162.790 40.215 162.790 40.170 162.740 40.170 ;
        RECT 162.790 40.170 165.575 40.215 ;
        POLYGON 162.740 40.170 162.740 40.140 162.705 40.140 ;
        RECT 162.740 40.140 165.575 40.170 ;
        RECT 117.460 40.135 154.280 40.140 ;
        POLYGON 154.280 40.140 154.685 40.135 154.280 40.135 ;
        POLYGON 154.845 40.140 154.845 40.135 154.685 40.135 ;
        RECT 154.845 40.135 159.700 40.140 ;
        RECT 117.460 40.020 159.700 40.135 ;
        POLYGON 159.700 40.140 159.930 40.140 159.700 40.020 ;
        POLYGON 162.705 40.140 162.705 40.040 162.595 40.040 ;
        RECT 162.705 40.040 165.575 40.140 ;
        POLYGON 162.595 40.040 162.595 40.020 162.570 40.020 ;
        RECT 162.595 40.020 165.575 40.040 ;
        RECT 117.460 40.005 159.470 40.020 ;
        POLYGON 117.460 40.005 117.480 40.005 117.480 39.755 ;
        RECT 117.480 39.900 159.470 40.005 ;
        POLYGON 159.470 40.020 159.695 40.020 159.470 39.900 ;
        POLYGON 162.570 40.020 162.570 39.930 162.460 39.930 ;
        RECT 162.570 39.930 165.575 40.020 ;
        POLYGON 162.460 39.930 162.460 39.900 162.420 39.900 ;
        RECT 162.460 39.925 165.575 39.930 ;
        POLYGON 165.575 40.245 165.845 40.245 165.575 39.925 ;
        POLYGON 169.455 40.245 169.455 40.115 169.375 40.115 ;
        RECT 169.455 40.240 174.425 40.245 ;
        POLYGON 174.425 41.305 174.845 41.305 174.425 40.240 ;
        POLYGON 182.435 41.305 182.435 41.000 182.375 41.000 ;
        RECT 182.435 41.000 198.000 41.305 ;
        POLYGON 182.375 41.000 182.375 40.240 182.230 40.240 ;
        RECT 182.375 40.240 198.000 41.000 ;
        RECT 169.455 40.115 174.025 40.240 ;
        POLYGON 169.375 40.115 169.375 39.930 169.260 39.930 ;
        RECT 169.375 39.930 174.025 40.115 ;
        RECT 162.460 39.900 165.475 39.925 ;
        RECT 117.480 39.890 159.445 39.900 ;
        POLYGON 159.445 39.900 159.470 39.900 159.445 39.890 ;
        POLYGON 162.420 39.900 162.420 39.890 162.410 39.890 ;
        RECT 162.420 39.890 165.475 39.900 ;
        RECT 117.480 39.770 159.200 39.890 ;
        POLYGON 159.200 39.890 159.445 39.890 159.200 39.770 ;
        POLYGON 162.410 39.890 162.410 39.770 162.255 39.770 ;
        RECT 162.410 39.810 165.475 39.890 ;
        POLYGON 165.475 39.925 165.575 39.925 165.475 39.810 ;
        POLYGON 169.260 39.925 169.260 39.815 169.190 39.815 ;
        RECT 169.260 39.815 174.025 39.930 ;
        RECT 162.410 39.770 165.115 39.810 ;
        RECT 117.480 39.700 158.785 39.770 ;
        POLYGON 117.480 39.700 117.510 39.700 117.510 39.330 ;
        RECT 117.510 39.570 158.785 39.700 ;
        POLYGON 158.785 39.770 159.200 39.770 158.785 39.570 ;
        POLYGON 162.255 39.770 162.255 39.695 162.160 39.695 ;
        RECT 162.255 39.695 165.115 39.770 ;
        POLYGON 162.160 39.695 162.160 39.665 162.120 39.665 ;
        RECT 162.160 39.665 165.115 39.695 ;
        POLYGON 162.120 39.665 162.120 39.625 162.065 39.625 ;
        RECT 162.120 39.625 165.115 39.665 ;
        POLYGON 162.065 39.625 162.065 39.595 162.025 39.595 ;
        RECT 162.065 39.595 165.115 39.625 ;
        POLYGON 162.025 39.595 162.025 39.570 161.990 39.570 ;
        RECT 162.025 39.570 165.115 39.595 ;
        RECT 117.510 39.555 158.755 39.570 ;
        POLYGON 158.755 39.570 158.785 39.570 158.755 39.555 ;
        POLYGON 161.990 39.570 161.990 39.555 161.970 39.555 ;
        RECT 161.990 39.555 165.115 39.570 ;
        RECT 117.510 39.530 158.690 39.555 ;
        POLYGON 158.690 39.555 158.755 39.555 158.690 39.530 ;
        POLYGON 161.970 39.555 161.970 39.530 161.935 39.530 ;
        RECT 161.970 39.530 165.115 39.555 ;
        RECT 117.510 39.320 158.210 39.530 ;
        POLYGON 158.210 39.530 158.690 39.530 158.210 39.320 ;
        POLYGON 161.935 39.530 161.935 39.365 161.715 39.365 ;
        RECT 161.935 39.410 165.115 39.530 ;
        POLYGON 165.115 39.810 165.475 39.810 165.115 39.410 ;
        POLYGON 169.190 39.810 169.190 39.765 169.160 39.765 ;
        RECT 169.190 39.765 174.025 39.815 ;
        POLYGON 169.160 39.765 169.160 39.670 169.105 39.670 ;
        RECT 169.160 39.670 174.025 39.765 ;
        POLYGON 169.105 39.670 169.105 39.640 169.085 39.640 ;
        RECT 169.105 39.640 174.025 39.670 ;
        POLYGON 169.085 39.640 169.085 39.635 169.080 39.635 ;
        RECT 169.085 39.635 174.025 39.640 ;
        POLYGON 169.080 39.635 169.080 39.600 169.060 39.600 ;
        RECT 169.080 39.600 174.025 39.635 ;
        POLYGON 169.060 39.600 169.060 39.545 169.020 39.545 ;
        RECT 169.060 39.545 174.025 39.600 ;
        POLYGON 169.020 39.545 169.020 39.460 168.965 39.460 ;
        RECT 169.020 39.460 174.025 39.545 ;
        POLYGON 168.965 39.460 168.965 39.410 168.930 39.410 ;
        RECT 168.965 39.410 174.025 39.460 ;
        RECT 161.935 39.380 165.090 39.410 ;
        POLYGON 165.090 39.410 165.115 39.410 165.090 39.380 ;
        POLYGON 168.930 39.405 168.930 39.385 168.915 39.385 ;
        RECT 168.930 39.385 174.025 39.410 ;
        RECT 161.935 39.365 165.045 39.380 ;
        POLYGON 161.715 39.365 161.715 39.340 161.675 39.340 ;
        RECT 161.715 39.340 165.045 39.365 ;
        POLYGON 161.675 39.340 161.675 39.320 161.645 39.320 ;
        RECT 161.675 39.335 165.045 39.340 ;
        POLYGON 165.045 39.380 165.090 39.380 165.045 39.335 ;
        POLYGON 168.915 39.380 168.915 39.345 168.890 39.345 ;
        RECT 168.915 39.345 174.025 39.385 ;
        POLYGON 168.890 39.345 168.890 39.340 168.885 39.340 ;
        RECT 168.890 39.340 174.025 39.345 ;
        RECT 168.885 39.335 174.025 39.340 ;
        POLYGON 174.025 40.240 174.425 40.240 174.025 39.335 ;
        POLYGON 182.230 40.230 182.230 40.175 182.220 40.175 ;
        RECT 182.230 40.175 198.000 40.240 ;
        POLYGON 182.220 40.175 182.220 39.525 182.060 39.525 ;
        RECT 182.220 39.525 198.000 40.175 ;
        POLYGON 182.060 39.525 182.060 39.335 182.015 39.335 ;
        RECT 182.060 39.495 198.000 39.525 ;
        POLYGON 198.000 41.790 198.075 41.790 198.000 39.495 ;
        POLYGON 208.805 43.145 209.390 43.145 209.390 41.645 ;
        RECT 209.390 43.000 223.620 43.145 ;
        POLYGON 223.620 43.625 223.855 43.000 223.620 43.000 ;
        POLYGON 230.695 43.625 230.745 43.625 230.745 43.505 ;
        RECT 230.745 43.505 234.820 43.625 ;
        POLYGON 230.745 43.505 230.795 43.505 230.795 43.380 ;
        RECT 230.795 43.380 234.820 43.505 ;
        POLYGON 230.795 43.380 230.955 43.380 230.955 43.005 ;
        RECT 230.955 43.310 234.820 43.380 ;
        POLYGON 234.820 43.940 235.135 43.310 234.820 43.310 ;
        POLYGON 237.765 43.940 237.780 43.940 237.780 43.915 ;
        RECT 237.780 43.915 239.955 43.940 ;
        POLYGON 237.780 43.915 238.135 43.915 238.135 43.335 ;
        RECT 238.135 43.880 239.955 43.915 ;
        POLYGON 239.955 43.945 239.995 43.880 239.955 43.880 ;
        POLYGON 241.720 43.945 241.775 43.945 241.775 43.880 ;
        RECT 241.775 43.920 243.110 43.945 ;
        POLYGON 243.110 44.055 243.235 43.920 243.110 43.920 ;
        POLYGON 244.355 44.055 244.425 44.055 244.425 43.995 ;
        RECT 244.425 44.000 245.445 44.055 ;
        POLYGON 245.445 44.080 245.550 44.000 245.445 44.000 ;
        POLYGON 246.615 44.080 246.725 44.080 246.725 44.025 ;
        RECT 246.725 44.045 247.615 44.080 ;
        POLYGON 247.615 44.080 247.690 44.045 247.615 44.045 ;
        POLYGON 252.080 44.080 252.080 44.045 252.005 44.045 ;
        RECT 252.080 44.060 253.085 44.080 ;
        POLYGON 253.085 44.095 253.145 44.095 253.085 44.060 ;
        POLYGON 254.235 44.095 254.235 44.075 254.215 44.075 ;
        RECT 254.235 44.090 255.290 44.095 ;
        POLYGON 255.290 44.095 255.295 44.095 255.290 44.090 ;
        POLYGON 256.330 44.095 256.330 44.090 256.325 44.090 ;
        RECT 256.330 44.090 257.535 44.095 ;
        RECT 254.235 44.075 255.165 44.090 ;
        POLYGON 254.215 44.075 254.215 44.060 254.195 44.060 ;
        RECT 254.215 44.060 255.165 44.075 ;
        RECT 252.080 44.045 253.010 44.060 ;
        RECT 246.725 44.025 247.690 44.045 ;
        POLYGON 247.690 44.045 247.730 44.025 247.690 44.025 ;
        POLYGON 252.005 44.045 252.005 44.025 251.960 44.025 ;
        RECT 252.005 44.025 253.010 44.045 ;
        POLYGON 246.725 44.025 246.740 44.025 246.740 44.015 ;
        RECT 246.740 44.015 247.730 44.025 ;
        POLYGON 246.740 44.015 246.770 44.015 246.770 44.000 ;
        RECT 246.770 44.000 247.730 44.015 ;
        RECT 244.425 43.995 245.550 44.000 ;
        POLYGON 244.425 43.995 244.510 43.995 244.510 43.920 ;
        RECT 244.510 43.960 245.550 43.995 ;
        POLYGON 245.550 44.000 245.615 43.960 245.550 43.960 ;
        POLYGON 246.770 44.000 246.855 44.000 246.855 43.960 ;
        RECT 246.855 43.985 247.730 44.000 ;
        POLYGON 247.730 44.025 247.830 43.985 247.730 43.985 ;
        POLYGON 251.960 44.025 251.960 44.020 251.950 44.020 ;
        RECT 251.960 44.020 253.010 44.025 ;
        POLYGON 253.010 44.060 253.085 44.060 253.010 44.020 ;
        POLYGON 254.195 44.060 254.195 44.020 254.135 44.020 ;
        RECT 254.195 44.020 255.165 44.060 ;
        POLYGON 251.950 44.020 251.950 44.010 251.920 44.010 ;
        RECT 251.950 44.010 252.930 44.020 ;
        POLYGON 251.920 44.010 251.920 43.985 251.860 43.985 ;
        RECT 251.920 43.985 252.930 44.010 ;
        RECT 246.855 43.960 247.830 43.985 ;
        POLYGON 247.830 43.985 247.895 43.960 247.830 43.960 ;
        POLYGON 251.860 43.985 251.860 43.960 251.800 43.960 ;
        RECT 251.860 43.975 252.930 43.985 ;
        POLYGON 252.930 44.020 253.010 44.020 252.930 43.975 ;
        POLYGON 254.135 44.020 254.135 43.975 254.075 43.975 ;
        RECT 254.135 43.975 255.165 44.020 ;
        POLYGON 255.165 44.090 255.290 44.090 255.165 43.980 ;
        POLYGON 256.325 44.090 256.325 44.030 256.275 44.030 ;
        RECT 256.325 44.030 257.410 44.090 ;
        POLYGON 256.275 44.030 256.275 44.020 256.265 44.020 ;
        RECT 256.275 44.020 257.410 44.030 ;
        POLYGON 256.265 44.020 256.265 43.995 256.245 43.995 ;
        RECT 256.265 43.995 257.410 44.020 ;
        POLYGON 256.245 43.995 256.245 43.980 256.230 43.980 ;
        RECT 256.245 43.980 257.410 43.995 ;
        RECT 251.860 43.960 252.680 43.975 ;
        RECT 244.510 43.940 245.615 43.960 ;
        POLYGON 245.615 43.960 245.640 43.940 245.615 43.940 ;
        POLYGON 246.855 43.960 246.895 43.960 246.895 43.940 ;
        RECT 246.895 43.940 247.895 43.960 ;
        RECT 244.510 43.920 245.640 43.940 ;
        RECT 241.775 43.905 243.235 43.920 ;
        POLYGON 243.235 43.920 243.245 43.905 243.235 43.905 ;
        POLYGON 244.510 43.920 244.530 43.920 244.530 43.905 ;
        RECT 244.530 43.905 245.640 43.920 ;
        RECT 241.775 43.880 243.245 43.905 ;
        RECT 238.135 43.865 239.995 43.880 ;
        POLYGON 239.995 43.880 240.005 43.865 239.995 43.865 ;
        POLYGON 241.775 43.880 241.785 43.880 241.785 43.865 ;
        RECT 241.785 43.865 243.245 43.880 ;
        RECT 238.135 43.740 240.005 43.865 ;
        POLYGON 240.005 43.865 240.095 43.740 240.005 43.740 ;
        POLYGON 241.785 43.865 241.865 43.865 241.865 43.765 ;
        RECT 241.865 43.765 243.245 43.865 ;
        POLYGON 241.865 43.765 241.880 43.765 241.880 43.745 ;
        RECT 241.880 43.755 243.245 43.765 ;
        POLYGON 243.245 43.905 243.395 43.755 243.245 43.755 ;
        POLYGON 244.530 43.905 244.585 43.905 244.585 43.860 ;
        RECT 244.585 43.860 245.640 43.905 ;
        POLYGON 244.590 43.860 244.700 43.860 244.700 43.765 ;
        RECT 244.700 43.835 245.640 43.860 ;
        POLYGON 245.640 43.940 245.785 43.835 245.640 43.835 ;
        POLYGON 246.895 43.940 246.985 43.940 246.985 43.900 ;
        RECT 246.985 43.935 247.895 43.940 ;
        POLYGON 247.895 43.960 247.945 43.935 247.895 43.935 ;
        POLYGON 251.800 43.960 251.800 43.950 251.775 43.950 ;
        RECT 251.800 43.950 252.680 43.960 ;
        POLYGON 251.775 43.950 251.775 43.935 251.735 43.935 ;
        RECT 251.775 43.935 252.680 43.950 ;
        RECT 246.985 43.925 247.945 43.935 ;
        POLYGON 247.945 43.935 247.975 43.925 247.945 43.925 ;
        POLYGON 251.735 43.935 251.735 43.925 251.710 43.925 ;
        RECT 251.735 43.925 252.680 43.935 ;
        RECT 246.985 43.900 247.975 43.925 ;
        POLYGON 246.985 43.900 247.000 43.900 247.000 43.895 ;
        RECT 247.000 43.895 247.975 43.900 ;
        POLYGON 247.000 43.895 247.075 43.895 247.075 43.860 ;
        RECT 247.075 43.875 247.975 43.895 ;
        POLYGON 247.975 43.925 248.110 43.875 247.975 43.875 ;
        POLYGON 251.710 43.925 251.710 43.905 251.665 43.905 ;
        RECT 251.710 43.905 252.680 43.925 ;
        POLYGON 251.660 43.905 251.660 43.890 251.610 43.890 ;
        RECT 251.660 43.890 252.680 43.905 ;
        POLYGON 251.610 43.890 251.610 43.880 251.595 43.880 ;
        RECT 251.610 43.880 252.680 43.890 ;
        POLYGON 251.595 43.880 251.595 43.875 251.580 43.875 ;
        RECT 251.595 43.875 252.680 43.880 ;
        RECT 247.075 43.860 248.110 43.875 ;
        POLYGON 247.075 43.860 247.130 43.860 247.130 43.835 ;
        RECT 247.130 43.855 248.110 43.860 ;
        POLYGON 248.110 43.875 248.160 43.855 248.110 43.855 ;
        POLYGON 251.580 43.875 251.580 43.855 251.520 43.855 ;
        RECT 251.580 43.855 252.680 43.875 ;
        RECT 247.130 43.850 248.160 43.855 ;
        POLYGON 248.160 43.855 248.175 43.850 248.160 43.850 ;
        POLYGON 251.520 43.855 251.520 43.850 251.505 43.850 ;
        RECT 251.520 43.850 252.680 43.855 ;
        POLYGON 252.680 43.975 252.930 43.975 252.680 43.850 ;
        POLYGON 254.075 43.975 254.075 43.940 254.020 43.940 ;
        RECT 254.075 43.940 255.070 43.975 ;
        POLYGON 254.020 43.940 254.020 43.920 253.995 43.920 ;
        RECT 254.020 43.920 255.070 43.940 ;
        POLYGON 253.995 43.920 253.995 43.850 253.890 43.850 ;
        RECT 253.995 43.890 255.070 43.920 ;
        POLYGON 255.070 43.975 255.165 43.975 255.070 43.890 ;
        POLYGON 256.230 43.980 256.230 43.895 256.155 43.895 ;
        RECT 256.230 43.920 257.410 43.980 ;
        POLYGON 257.410 44.090 257.535 44.090 257.410 43.920 ;
        POLYGON 259.100 44.090 259.100 43.955 259.020 43.955 ;
        RECT 259.100 43.955 260.695 44.095 ;
        POLYGON 259.020 43.955 259.020 43.940 259.010 43.940 ;
        RECT 259.020 43.940 260.695 43.955 ;
        POLYGON 259.010 43.940 259.010 43.920 258.995 43.920 ;
        RECT 259.010 43.925 260.695 43.940 ;
        POLYGON 260.695 44.095 260.780 44.095 260.695 43.925 ;
        POLYGON 263.130 44.095 263.130 44.030 263.110 44.030 ;
        RECT 263.130 44.085 266.075 44.095 ;
        POLYGON 266.075 44.095 266.080 44.095 266.075 44.085 ;
        POLYGON 270.575 44.095 270.575 44.085 270.570 44.085 ;
        RECT 270.575 44.085 277.780 44.135 ;
        POLYGON 277.780 44.215 277.795 44.215 277.780 44.095 ;
        POLYGON 287.785 44.210 287.785 44.110 287.780 44.110 ;
        RECT 287.785 44.110 303.120 44.215 ;
        RECT 263.130 44.030 265.950 44.085 ;
        POLYGON 263.110 44.030 263.110 43.930 263.070 43.930 ;
        RECT 263.110 43.930 265.950 44.030 ;
        RECT 259.010 43.920 260.420 43.925 ;
        RECT 256.230 43.895 257.275 43.920 ;
        RECT 253.995 43.850 254.865 43.890 ;
        RECT 247.130 43.835 248.180 43.850 ;
        RECT 244.700 43.815 245.785 43.835 ;
        POLYGON 245.785 43.835 245.820 43.815 245.785 43.815 ;
        POLYGON 247.130 43.835 247.180 43.835 247.180 43.815 ;
        RECT 247.180 43.820 248.180 43.835 ;
        POLYGON 248.180 43.850 248.265 43.820 248.180 43.820 ;
        POLYGON 251.505 43.850 251.505 43.820 251.425 43.820 ;
        RECT 251.505 43.820 252.525 43.850 ;
        RECT 247.180 43.815 248.265 43.820 ;
        RECT 244.700 43.805 245.820 43.815 ;
        POLYGON 245.820 43.815 245.840 43.805 245.820 43.805 ;
        POLYGON 247.180 43.815 247.200 43.815 247.200 43.805 ;
        RECT 247.200 43.805 248.265 43.815 ;
        RECT 244.700 43.800 245.840 43.805 ;
        POLYGON 245.840 43.805 245.845 43.800 245.840 43.800 ;
        POLYGON 247.200 43.805 247.215 43.805 247.215 43.800 ;
        RECT 247.215 43.800 248.265 43.805 ;
        RECT 244.700 43.765 245.845 43.800 ;
        POLYGON 244.700 43.765 244.710 43.765 244.710 43.755 ;
        RECT 244.710 43.755 245.845 43.765 ;
        RECT 241.880 43.740 243.395 43.755 ;
        RECT 238.135 43.680 240.095 43.740 ;
        POLYGON 240.095 43.740 240.140 43.680 240.095 43.680 ;
        POLYGON 241.880 43.740 241.935 43.740 241.935 43.680 ;
        RECT 241.935 43.710 243.395 43.740 ;
        POLYGON 243.395 43.755 243.435 43.710 243.395 43.710 ;
        POLYGON 244.710 43.755 244.770 43.755 244.770 43.710 ;
        RECT 244.770 43.710 245.845 43.755 ;
        RECT 241.935 43.680 243.435 43.710 ;
        RECT 238.135 43.585 240.140 43.680 ;
        POLYGON 240.140 43.680 240.210 43.585 240.140 43.585 ;
        POLYGON 241.935 43.680 242.015 43.680 242.015 43.585 ;
        RECT 242.015 43.585 243.435 43.680 ;
        RECT 238.135 43.560 240.210 43.585 ;
        POLYGON 240.210 43.585 240.225 43.560 240.210 43.560 ;
        POLYGON 242.015 43.585 242.040 43.585 242.040 43.560 ;
        RECT 242.040 43.560 243.435 43.585 ;
        POLYGON 243.435 43.710 243.585 43.560 243.435 43.560 ;
        POLYGON 244.770 43.710 244.840 43.710 244.840 43.660 ;
        RECT 244.840 43.685 245.845 43.710 ;
        POLYGON 245.845 43.800 246.020 43.685 245.845 43.685 ;
        POLYGON 247.215 43.800 247.250 43.800 247.250 43.785 ;
        RECT 247.250 43.785 248.265 43.800 ;
        POLYGON 247.250 43.785 247.275 43.785 247.275 43.775 ;
        RECT 247.275 43.780 248.265 43.785 ;
        POLYGON 248.265 43.820 248.375 43.780 248.265 43.780 ;
        POLYGON 251.425 43.820 251.425 43.815 251.410 43.815 ;
        RECT 251.425 43.815 252.525 43.820 ;
        POLYGON 251.410 43.815 251.410 43.810 251.400 43.810 ;
        RECT 251.410 43.810 252.525 43.815 ;
        POLYGON 251.400 43.810 251.400 43.780 251.305 43.780 ;
        RECT 251.400 43.780 252.525 43.810 ;
        POLYGON 252.525 43.850 252.680 43.850 252.525 43.780 ;
        POLYGON 253.890 43.850 253.890 43.840 253.870 43.840 ;
        RECT 253.890 43.840 254.865 43.850 ;
        POLYGON 253.870 43.840 253.870 43.805 253.820 43.805 ;
        RECT 253.870 43.805 254.865 43.840 ;
        POLYGON 253.820 43.805 253.820 43.780 253.775 43.780 ;
        RECT 253.820 43.780 254.865 43.805 ;
        RECT 247.275 43.775 248.375 43.780 ;
        POLYGON 248.375 43.780 248.390 43.775 248.375 43.775 ;
        POLYGON 251.305 43.780 251.305 43.775 251.290 43.775 ;
        RECT 251.305 43.775 252.510 43.780 ;
        POLYGON 252.510 43.780 252.525 43.780 252.510 43.775 ;
        POLYGON 253.775 43.780 253.775 43.775 253.770 43.775 ;
        RECT 253.775 43.775 254.865 43.780 ;
        POLYGON 247.275 43.775 247.510 43.775 247.510 43.685 ;
        RECT 247.510 43.750 248.390 43.775 ;
        POLYGON 248.390 43.775 248.470 43.750 248.390 43.750 ;
        POLYGON 251.290 43.775 251.290 43.770 251.275 43.770 ;
        RECT 251.290 43.770 252.435 43.775 ;
        POLYGON 251.275 43.770 251.275 43.755 251.225 43.755 ;
        RECT 251.275 43.755 252.435 43.770 ;
        POLYGON 251.225 43.755 251.225 43.750 251.205 43.750 ;
        RECT 251.225 43.750 252.435 43.755 ;
        RECT 247.510 43.725 248.475 43.750 ;
        POLYGON 248.475 43.750 248.565 43.725 248.475 43.725 ;
        POLYGON 251.205 43.750 251.205 43.730 251.135 43.730 ;
        RECT 251.205 43.740 252.435 43.750 ;
        POLYGON 252.435 43.775 252.510 43.775 252.435 43.740 ;
        POLYGON 253.770 43.775 253.770 43.765 253.750 43.765 ;
        RECT 253.770 43.765 254.865 43.775 ;
        POLYGON 253.750 43.765 253.750 43.740 253.715 43.740 ;
        RECT 253.750 43.740 254.865 43.765 ;
        RECT 251.205 43.730 252.255 43.740 ;
        POLYGON 251.135 43.730 251.135 43.725 251.120 43.725 ;
        RECT 251.135 43.725 252.255 43.730 ;
        RECT 247.510 43.715 248.565 43.725 ;
        POLYGON 248.565 43.725 248.590 43.715 248.565 43.715 ;
        POLYGON 251.120 43.725 251.120 43.715 251.095 43.715 ;
        RECT 251.120 43.715 252.255 43.725 ;
        RECT 247.510 43.695 248.590 43.715 ;
        POLYGON 248.590 43.715 248.665 43.695 248.590 43.695 ;
        POLYGON 251.095 43.715 251.095 43.695 251.015 43.695 ;
        RECT 251.095 43.695 252.255 43.715 ;
        RECT 247.510 43.685 248.665 43.695 ;
        RECT 244.840 43.675 246.020 43.685 ;
        POLYGON 246.020 43.685 246.035 43.675 246.020 43.675 ;
        POLYGON 247.515 43.685 247.540 43.685 247.540 43.675 ;
        RECT 247.540 43.675 248.665 43.685 ;
        RECT 244.840 43.665 246.035 43.675 ;
        POLYGON 246.035 43.675 246.055 43.665 246.035 43.665 ;
        POLYGON 247.540 43.675 247.555 43.675 247.555 43.670 ;
        RECT 247.555 43.670 248.665 43.675 ;
        POLYGON 248.665 43.695 248.775 43.670 248.665 43.670 ;
        POLYGON 251.015 43.695 251.015 43.670 250.925 43.670 ;
        RECT 251.015 43.670 252.255 43.695 ;
        POLYGON 252.255 43.740 252.435 43.740 252.255 43.670 ;
        POLYGON 253.715 43.740 253.715 43.695 253.645 43.695 ;
        RECT 253.715 43.710 254.865 43.740 ;
        POLYGON 254.865 43.890 255.070 43.890 254.865 43.710 ;
        POLYGON 256.155 43.890 256.155 43.805 256.070 43.805 ;
        RECT 256.155 43.805 257.275 43.895 ;
        POLYGON 256.070 43.805 256.070 43.740 256.015 43.740 ;
        RECT 256.070 43.755 257.275 43.805 ;
        POLYGON 257.275 43.920 257.410 43.920 257.275 43.755 ;
        POLYGON 258.995 43.915 258.995 43.810 258.925 43.810 ;
        RECT 258.995 43.810 260.420 43.920 ;
        POLYGON 258.925 43.810 258.925 43.755 258.890 43.755 ;
        RECT 258.925 43.755 260.420 43.810 ;
        RECT 256.070 43.740 257.200 43.755 ;
        POLYGON 256.015 43.740 256.015 43.735 256.005 43.735 ;
        RECT 256.015 43.735 257.200 43.740 ;
        POLYGON 256.005 43.735 256.005 43.710 255.980 43.710 ;
        RECT 256.005 43.710 257.200 43.735 ;
        RECT 253.715 43.700 254.850 43.710 ;
        POLYGON 254.850 43.710 254.860 43.710 254.850 43.700 ;
        POLYGON 255.980 43.710 255.980 43.700 255.975 43.700 ;
        RECT 255.980 43.700 257.200 43.710 ;
        RECT 253.715 43.695 254.615 43.700 ;
        POLYGON 253.640 43.695 253.640 43.680 253.620 43.680 ;
        RECT 253.640 43.680 254.615 43.695 ;
        POLYGON 253.615 43.680 253.615 43.670 253.600 43.670 ;
        RECT 253.615 43.670 254.615 43.680 ;
        POLYGON 247.555 43.670 247.565 43.670 247.565 43.665 ;
        RECT 247.565 43.665 248.775 43.670 ;
        RECT 244.840 43.660 246.055 43.665 ;
        POLYGON 244.845 43.660 244.970 43.660 244.970 43.560 ;
        RECT 244.970 43.560 246.055 43.660 ;
        RECT 238.135 43.440 240.225 43.560 ;
        POLYGON 240.225 43.560 240.315 43.440 240.225 43.440 ;
        POLYGON 242.040 43.560 242.105 43.560 242.105 43.485 ;
        RECT 242.105 43.520 243.585 43.560 ;
        POLYGON 243.585 43.560 243.630 43.520 243.585 43.520 ;
        POLYGON 244.970 43.560 245.025 43.560 245.025 43.520 ;
        RECT 245.025 43.550 246.055 43.560 ;
        POLYGON 246.055 43.665 246.240 43.550 246.055 43.550 ;
        POLYGON 247.565 43.665 247.785 43.665 247.785 43.590 ;
        RECT 247.785 43.660 248.775 43.665 ;
        POLYGON 248.775 43.670 248.805 43.660 248.775 43.660 ;
        POLYGON 250.925 43.670 250.925 43.660 250.880 43.660 ;
        RECT 250.925 43.660 252.180 43.670 ;
        RECT 247.785 43.630 248.805 43.660 ;
        POLYGON 248.805 43.660 248.945 43.630 248.805 43.630 ;
        RECT 250.865 43.655 252.180 43.660 ;
        POLYGON 250.845 43.655 250.845 43.630 250.735 43.630 ;
        RECT 250.845 43.640 252.180 43.655 ;
        POLYGON 252.180 43.670 252.255 43.670 252.180 43.640 ;
        POLYGON 253.600 43.670 253.600 43.640 253.545 43.640 ;
        RECT 253.600 43.640 254.615 43.670 ;
        RECT 250.845 43.630 252.065 43.640 ;
        RECT 247.785 43.615 248.945 43.630 ;
        POLYGON 248.945 43.630 249.020 43.615 248.945 43.615 ;
        POLYGON 250.735 43.630 250.735 43.615 250.670 43.615 ;
        RECT 250.735 43.615 252.065 43.630 ;
        RECT 247.785 43.605 249.020 43.615 ;
        POLYGON 249.020 43.615 249.085 43.605 249.020 43.605 ;
        POLYGON 250.650 43.615 250.650 43.605 250.600 43.605 ;
        RECT 250.650 43.605 252.065 43.615 ;
        RECT 247.785 43.590 249.085 43.605 ;
        POLYGON 247.785 43.590 247.830 43.590 247.830 43.575 ;
        RECT 247.830 43.585 249.085 43.590 ;
        POLYGON 249.085 43.605 249.190 43.585 249.085 43.585 ;
        RECT 250.595 43.600 252.065 43.605 ;
        POLYGON 252.065 43.640 252.180 43.640 252.065 43.600 ;
        POLYGON 253.545 43.640 253.545 43.615 253.505 43.615 ;
        RECT 253.545 43.615 254.615 43.640 ;
        POLYGON 253.505 43.615 253.505 43.600 253.480 43.600 ;
        RECT 253.505 43.600 254.615 43.615 ;
        POLYGON 250.590 43.600 250.590 43.595 250.560 43.595 ;
        RECT 250.590 43.595 252.000 43.600 ;
        POLYGON 250.560 43.595 250.560 43.585 250.495 43.585 ;
        RECT 250.560 43.585 252.000 43.595 ;
        RECT 247.830 43.580 249.190 43.585 ;
        POLYGON 249.190 43.585 249.220 43.580 249.190 43.580 ;
        POLYGON 250.495 43.585 250.495 43.580 250.465 43.580 ;
        RECT 250.495 43.580 252.000 43.585 ;
        RECT 247.830 43.575 249.230 43.580 ;
        POLYGON 247.830 43.575 247.910 43.575 247.910 43.550 ;
        RECT 247.910 43.560 249.230 43.575 ;
        POLYGON 249.230 43.580 249.400 43.560 249.230 43.560 ;
        POLYGON 250.455 43.580 250.455 43.560 250.325 43.560 ;
        RECT 250.455 43.575 252.000 43.580 ;
        POLYGON 252.000 43.600 252.065 43.600 252.000 43.575 ;
        POLYGON 253.480 43.600 253.480 43.575 253.435 43.575 ;
        RECT 253.480 43.575 254.615 43.600 ;
        RECT 250.455 43.560 251.920 43.575 ;
        RECT 247.910 43.555 249.400 43.560 ;
        POLYGON 249.400 43.560 249.440 43.555 249.400 43.555 ;
        POLYGON 250.315 43.560 250.315 43.555 250.260 43.555 ;
        RECT 250.315 43.555 251.920 43.560 ;
        RECT 247.910 43.550 249.440 43.555 ;
        POLYGON 249.440 43.555 249.495 43.550 249.440 43.550 ;
        POLYGON 250.255 43.555 250.255 43.550 250.205 43.550 ;
        RECT 250.255 43.550 251.920 43.555 ;
        POLYGON 251.920 43.575 252.000 43.575 251.920 43.550 ;
        POLYGON 253.435 43.575 253.435 43.560 253.410 43.560 ;
        RECT 253.435 43.560 254.615 43.575 ;
        POLYGON 253.405 43.560 253.405 43.550 253.390 43.550 ;
        RECT 253.405 43.550 254.615 43.560 ;
        RECT 245.025 43.540 246.240 43.550 ;
        POLYGON 246.240 43.550 246.255 43.540 246.240 43.540 ;
        POLYGON 247.910 43.550 247.945 43.550 247.945 43.540 ;
        RECT 247.945 43.540 249.515 43.550 ;
        RECT 245.025 43.530 246.260 43.540 ;
        POLYGON 246.260 43.540 246.275 43.530 246.260 43.530 ;
        POLYGON 247.945 43.540 247.975 43.540 247.975 43.530 ;
        RECT 247.975 43.535 249.515 43.540 ;
        POLYGON 249.515 43.550 249.650 43.535 249.515 43.535 ;
        POLYGON 250.205 43.550 250.205 43.535 250.055 43.535 ;
        RECT 250.205 43.535 251.745 43.550 ;
        RECT 247.975 43.530 249.845 43.535 ;
        POLYGON 249.845 43.535 249.860 43.530 249.845 43.530 ;
        POLYGON 250.050 43.535 250.050 43.530 249.860 43.530 ;
        RECT 250.050 43.530 251.745 43.535 ;
        RECT 245.025 43.520 246.275 43.530 ;
        RECT 242.105 43.485 243.630 43.520 ;
        POLYGON 242.105 43.485 242.140 43.485 242.140 43.440 ;
        RECT 242.140 43.455 243.630 43.485 ;
        POLYGON 243.630 43.520 243.695 43.455 243.630 43.455 ;
        POLYGON 245.025 43.520 245.065 43.520 245.065 43.490 ;
        RECT 245.065 43.490 246.275 43.520 ;
        POLYGON 245.065 43.490 245.110 43.490 245.110 43.465 ;
        RECT 245.110 43.465 246.275 43.490 ;
        POLYGON 245.110 43.465 245.120 43.465 245.120 43.455 ;
        RECT 245.120 43.455 246.275 43.465 ;
        RECT 242.140 43.440 243.695 43.455 ;
        RECT 238.135 43.425 240.315 43.440 ;
        POLYGON 240.315 43.440 240.325 43.425 240.315 43.425 ;
        POLYGON 242.140 43.440 242.155 43.440 242.155 43.425 ;
        RECT 242.155 43.425 243.695 43.440 ;
        RECT 238.135 43.420 240.325 43.425 ;
        POLYGON 240.325 43.425 240.330 43.420 240.325 43.420 ;
        POLYGON 242.155 43.425 242.160 43.425 242.160 43.420 ;
        RECT 242.160 43.420 243.695 43.425 ;
        RECT 238.135 43.335 240.330 43.420 ;
        POLYGON 238.135 43.335 238.150 43.335 238.150 43.310 ;
        RECT 238.150 43.310 240.330 43.335 ;
        RECT 230.955 43.265 235.135 43.310 ;
        POLYGON 235.135 43.310 235.160 43.265 235.135 43.265 ;
        POLYGON 238.150 43.310 238.180 43.310 238.180 43.265 ;
        RECT 238.180 43.265 240.330 43.310 ;
        RECT 230.955 43.235 235.160 43.265 ;
        POLYGON 235.160 43.265 235.175 43.235 235.160 43.235 ;
        POLYGON 238.180 43.265 238.200 43.265 238.200 43.235 ;
        RECT 238.200 43.255 240.330 43.265 ;
        POLYGON 240.330 43.420 240.460 43.255 240.330 43.255 ;
        POLYGON 242.160 43.420 242.185 43.420 242.185 43.390 ;
        RECT 242.185 43.390 243.695 43.420 ;
        POLYGON 242.185 43.390 242.315 43.390 242.315 43.255 ;
        RECT 242.315 43.290 243.695 43.390 ;
        POLYGON 243.695 43.455 243.870 43.290 243.695 43.290 ;
        POLYGON 245.120 43.455 245.265 43.455 245.265 43.360 ;
        RECT 245.265 43.415 246.275 43.455 ;
        POLYGON 246.275 43.530 246.490 43.415 246.275 43.415 ;
        POLYGON 247.975 43.530 248.050 43.530 248.050 43.505 ;
        RECT 248.050 43.505 251.745 43.530 ;
        POLYGON 248.050 43.505 248.110 43.505 248.110 43.490 ;
        RECT 248.110 43.495 251.745 43.505 ;
        POLYGON 251.745 43.550 251.920 43.550 251.745 43.495 ;
        POLYGON 253.390 43.550 253.390 43.530 253.355 43.530 ;
        RECT 253.390 43.530 254.615 43.550 ;
        POLYGON 253.355 43.530 253.355 43.495 253.290 43.495 ;
        RECT 253.355 43.515 254.615 43.530 ;
        POLYGON 254.615 43.700 254.850 43.700 254.615 43.515 ;
        POLYGON 255.975 43.700 255.975 43.610 255.890 43.610 ;
        RECT 255.975 43.660 257.200 43.700 ;
        POLYGON 257.200 43.755 257.275 43.755 257.200 43.660 ;
        POLYGON 258.890 43.755 258.890 43.665 258.830 43.665 ;
        RECT 258.890 43.665 260.420 43.755 ;
        POLYGON 258.830 43.665 258.830 43.660 258.825 43.660 ;
        RECT 258.830 43.660 260.420 43.665 ;
        RECT 255.975 43.620 257.165 43.660 ;
        POLYGON 257.165 43.660 257.200 43.660 257.165 43.620 ;
        POLYGON 258.825 43.660 258.825 43.650 258.820 43.650 ;
        RECT 258.825 43.650 260.420 43.660 ;
        POLYGON 258.820 43.650 258.820 43.620 258.800 43.620 ;
        RECT 258.820 43.620 260.420 43.650 ;
        RECT 255.975 43.610 256.985 43.620 ;
        POLYGON 255.890 43.610 255.890 43.605 255.885 43.605 ;
        RECT 255.890 43.605 256.985 43.610 ;
        POLYGON 255.885 43.605 255.885 43.515 255.790 43.515 ;
        RECT 255.885 43.515 256.985 43.605 ;
        RECT 253.355 43.495 254.550 43.515 ;
        RECT 248.110 43.490 251.660 43.495 ;
        POLYGON 248.110 43.490 248.320 43.490 248.320 43.435 ;
        RECT 248.320 43.470 251.660 43.490 ;
        POLYGON 251.660 43.495 251.745 43.495 251.660 43.470 ;
        POLYGON 253.290 43.495 253.290 43.470 253.240 43.470 ;
        RECT 253.290 43.470 254.550 43.495 ;
        RECT 248.320 43.455 251.605 43.470 ;
        POLYGON 251.605 43.470 251.660 43.470 251.605 43.455 ;
        POLYGON 253.240 43.470 253.240 43.455 253.210 43.455 ;
        RECT 253.240 43.465 254.550 43.470 ;
        POLYGON 254.550 43.515 254.615 43.515 254.550 43.465 ;
        POLYGON 255.790 43.515 255.790 43.465 255.740 43.465 ;
        RECT 255.790 43.465 256.985 43.515 ;
        RECT 253.240 43.460 254.545 43.465 ;
        POLYGON 254.545 43.465 254.550 43.465 254.545 43.460 ;
        POLYGON 255.740 43.465 255.740 43.460 255.735 43.460 ;
        RECT 255.740 43.460 256.985 43.465 ;
        RECT 253.240 43.455 254.380 43.460 ;
        RECT 248.320 43.435 251.485 43.455 ;
        POLYGON 248.320 43.435 248.390 43.435 248.390 43.420 ;
        RECT 248.390 43.425 251.485 43.435 ;
        POLYGON 251.485 43.455 251.605 43.455 251.485 43.425 ;
        POLYGON 253.210 43.455 253.210 43.425 253.150 43.425 ;
        RECT 253.210 43.425 254.380 43.455 ;
        RECT 248.390 43.420 251.400 43.425 ;
        POLYGON 248.390 43.420 248.410 43.420 248.410 43.415 ;
        RECT 248.410 43.415 251.400 43.420 ;
        RECT 245.265 43.405 246.490 43.415 ;
        POLYGON 246.490 43.415 246.500 43.405 246.490 43.405 ;
        POLYGON 248.410 43.415 248.455 43.415 248.455 43.405 ;
        RECT 248.455 43.405 251.400 43.415 ;
        RECT 245.265 43.360 246.505 43.405 ;
        POLYGON 245.265 43.360 245.365 43.360 245.365 43.290 ;
        RECT 245.365 43.295 246.505 43.360 ;
        POLYGON 246.505 43.405 246.725 43.295 246.505 43.295 ;
        POLYGON 248.455 43.405 248.585 43.405 248.585 43.375 ;
        RECT 248.585 43.400 251.400 43.405 ;
        POLYGON 251.400 43.425 251.485 43.425 251.400 43.400 ;
        POLYGON 253.150 43.425 253.150 43.400 253.095 43.400 ;
        RECT 253.150 43.400 254.380 43.425 ;
        RECT 248.585 43.375 251.230 43.400 ;
        POLYGON 248.585 43.375 248.665 43.375 248.665 43.360 ;
        RECT 248.665 43.365 251.230 43.375 ;
        POLYGON 251.230 43.400 251.400 43.400 251.230 43.365 ;
        POLYGON 253.095 43.400 253.095 43.395 253.085 43.395 ;
        RECT 253.095 43.395 254.380 43.400 ;
        POLYGON 253.085 43.395 253.085 43.365 253.030 43.365 ;
        RECT 253.085 43.365 254.380 43.395 ;
        RECT 248.665 43.360 251.145 43.365 ;
        POLYGON 248.665 43.360 248.840 43.360 248.840 43.330 ;
        RECT 248.840 43.350 251.145 43.360 ;
        POLYGON 251.145 43.365 251.225 43.365 251.145 43.350 ;
        POLYGON 253.030 43.365 253.030 43.350 253.000 43.350 ;
        RECT 253.030 43.350 254.380 43.365 ;
        RECT 248.840 43.345 251.135 43.350 ;
        POLYGON 251.135 43.350 251.145 43.350 251.135 43.345 ;
        POLYGON 253.000 43.350 253.000 43.345 252.990 43.345 ;
        RECT 253.000 43.345 254.380 43.350 ;
        RECT 248.840 43.330 250.965 43.345 ;
        POLYGON 248.850 43.330 248.945 43.330 248.945 43.310 ;
        RECT 248.945 43.320 250.965 43.330 ;
        POLYGON 250.965 43.345 251.135 43.345 250.965 43.320 ;
        POLYGON 252.990 43.345 252.990 43.335 252.965 43.335 ;
        RECT 252.990 43.340 254.380 43.345 ;
        POLYGON 254.380 43.460 254.545 43.460 254.380 43.340 ;
        POLYGON 255.735 43.460 255.735 43.425 255.695 43.425 ;
        RECT 255.735 43.425 256.985 43.460 ;
        POLYGON 255.695 43.425 255.695 43.340 255.610 43.340 ;
        RECT 255.695 43.405 256.985 43.425 ;
        POLYGON 256.985 43.620 257.165 43.620 256.985 43.405 ;
        POLYGON 258.800 43.615 258.800 43.600 258.790 43.600 ;
        RECT 258.800 43.600 260.420 43.620 ;
        POLYGON 258.790 43.600 258.790 43.520 258.735 43.520 ;
        RECT 258.790 43.520 260.420 43.600 ;
        POLYGON 258.735 43.520 258.735 43.475 258.705 43.475 ;
        RECT 258.735 43.475 260.420 43.520 ;
        POLYGON 258.705 43.475 258.705 43.405 258.655 43.405 ;
        RECT 258.705 43.430 260.420 43.475 ;
        POLYGON 260.420 43.925 260.695 43.925 260.420 43.430 ;
        POLYGON 263.070 43.925 263.070 43.820 263.025 43.820 ;
        RECT 263.070 43.820 265.950 43.930 ;
        POLYGON 263.025 43.820 263.025 43.805 263.020 43.805 ;
        RECT 263.025 43.805 265.950 43.820 ;
        POLYGON 263.020 43.805 263.020 43.510 262.900 43.510 ;
        RECT 263.020 43.675 265.950 43.805 ;
        POLYGON 265.950 44.085 266.075 44.085 265.950 43.675 ;
        RECT 270.570 44.075 277.780 44.085 ;
        POLYGON 270.570 44.055 270.570 43.705 270.520 43.705 ;
        RECT 270.570 43.705 277.650 44.075 ;
        POLYGON 270.520 43.705 270.520 43.680 270.515 43.680 ;
        RECT 270.520 43.680 277.650 43.705 ;
        RECT 263.020 43.510 265.900 43.675 ;
        POLYGON 262.900 43.510 262.900 43.430 262.865 43.430 ;
        RECT 262.900 43.505 265.900 43.510 ;
        POLYGON 265.900 43.675 265.950 43.675 265.900 43.505 ;
        POLYGON 270.515 43.675 270.515 43.600 270.500 43.600 ;
        RECT 270.515 43.600 277.650 43.680 ;
        POLYGON 270.500 43.600 270.500 43.515 270.485 43.515 ;
        RECT 270.500 43.515 277.650 43.600 ;
        RECT 262.900 43.430 265.850 43.505 ;
        RECT 258.705 43.405 260.385 43.430 ;
        RECT 255.695 43.345 256.930 43.405 ;
        POLYGON 256.930 43.405 256.985 43.405 256.930 43.345 ;
        POLYGON 258.655 43.405 258.655 43.345 258.610 43.345 ;
        RECT 258.655 43.365 260.385 43.405 ;
        POLYGON 260.385 43.430 260.420 43.430 260.385 43.365 ;
        POLYGON 262.865 43.430 262.865 43.365 262.835 43.365 ;
        RECT 262.865 43.365 265.850 43.430 ;
        POLYGON 265.850 43.505 265.900 43.505 265.850 43.365 ;
        POLYGON 270.485 43.505 270.485 43.375 270.460 43.375 ;
        RECT 270.485 43.375 277.650 43.515 ;
        RECT 258.655 43.345 260.145 43.365 ;
        RECT 255.695 43.340 256.755 43.345 ;
        RECT 252.990 43.335 254.230 43.340 ;
        POLYGON 252.965 43.335 252.965 43.320 252.930 43.320 ;
        RECT 252.965 43.320 254.230 43.335 ;
        RECT 248.945 43.310 250.865 43.320 ;
        POLYGON 248.945 43.310 249.070 43.310 249.070 43.295 ;
        RECT 249.070 43.300 250.865 43.310 ;
        POLYGON 250.865 43.320 250.965 43.320 250.865 43.300 ;
        POLYGON 252.930 43.320 252.930 43.300 252.885 43.300 ;
        RECT 252.930 43.300 254.230 43.320 ;
        RECT 249.070 43.295 250.710 43.300 ;
        RECT 245.365 43.290 246.725 43.295 ;
        RECT 242.315 43.260 243.870 43.290 ;
        POLYGON 243.870 43.290 243.900 43.260 243.870 43.260 ;
        POLYGON 245.365 43.290 245.380 43.290 245.380 43.280 ;
        RECT 245.380 43.285 246.725 43.290 ;
        POLYGON 246.725 43.295 246.740 43.285 246.725 43.285 ;
        POLYGON 249.070 43.295 249.115 43.295 249.115 43.290 ;
        RECT 249.115 43.290 250.710 43.295 ;
        POLYGON 249.120 43.290 249.155 43.290 249.155 43.285 ;
        RECT 249.155 43.285 250.710 43.290 ;
        RECT 245.380 43.280 246.745 43.285 ;
        POLYGON 245.380 43.280 245.405 43.280 245.405 43.260 ;
        RECT 245.405 43.260 246.745 43.280 ;
        RECT 242.315 43.255 243.900 43.260 ;
        RECT 238.200 43.235 240.460 43.255 ;
        RECT 230.955 43.200 235.175 43.235 ;
        POLYGON 235.175 43.235 235.190 43.200 235.175 43.200 ;
        POLYGON 238.200 43.235 238.225 43.235 238.225 43.200 ;
        RECT 238.225 43.200 240.460 43.235 ;
        RECT 230.955 43.000 235.190 43.200 ;
        RECT 209.390 42.355 223.855 43.000 ;
        POLYGON 223.855 43.000 224.120 42.355 223.855 42.355 ;
        POLYGON 230.955 43.000 231.005 43.000 231.005 42.890 ;
        RECT 231.005 42.890 235.190 43.000 ;
        POLYGON 231.005 42.890 231.060 42.890 231.060 42.760 ;
        RECT 231.060 42.760 235.190 42.890 ;
        POLYGON 231.060 42.760 231.140 42.760 231.140 42.590 ;
        RECT 231.140 42.590 235.190 42.760 ;
        POLYGON 231.140 42.590 231.245 42.590 231.245 42.365 ;
        RECT 231.245 42.525 235.190 42.590 ;
        POLYGON 235.190 43.200 235.575 42.525 235.190 42.525 ;
        POLYGON 238.225 43.200 238.320 43.200 238.320 43.065 ;
        RECT 238.320 43.165 240.460 43.200 ;
        POLYGON 240.460 43.255 240.530 43.165 240.460 43.165 ;
        POLYGON 242.315 43.255 242.340 43.255 242.340 43.230 ;
        RECT 242.340 43.230 243.900 43.255 ;
        POLYGON 242.340 43.230 242.400 43.230 242.400 43.165 ;
        RECT 242.400 43.165 243.900 43.230 ;
        RECT 238.320 43.070 240.530 43.165 ;
        POLYGON 240.530 43.165 240.600 43.070 240.530 43.070 ;
        POLYGON 242.400 43.165 242.490 43.165 242.490 43.070 ;
        RECT 242.490 43.160 243.900 43.165 ;
        POLYGON 243.900 43.260 244.015 43.160 243.900 43.160 ;
        POLYGON 245.405 43.260 245.445 43.260 245.445 43.235 ;
        RECT 245.445 43.235 246.745 43.260 ;
        POLYGON 245.445 43.235 245.570 43.235 245.570 43.160 ;
        RECT 245.570 43.170 246.745 43.235 ;
        POLYGON 246.745 43.285 246.985 43.170 246.745 43.170 ;
        POLYGON 249.155 43.285 249.225 43.285 249.225 43.275 ;
        RECT 249.225 43.280 250.710 43.285 ;
        POLYGON 250.710 43.300 250.865 43.300 250.710 43.280 ;
        POLYGON 252.885 43.300 252.885 43.280 252.845 43.280 ;
        RECT 252.885 43.280 254.230 43.300 ;
        RECT 249.225 43.275 250.595 43.280 ;
        POLYGON 249.225 43.275 249.290 43.275 249.290 43.270 ;
        RECT 249.290 43.270 250.595 43.275 ;
        POLYGON 250.595 43.280 250.675 43.280 250.595 43.270 ;
        POLYGON 252.845 43.280 252.845 43.270 252.820 43.270 ;
        RECT 252.845 43.270 254.230 43.280 ;
        POLYGON 249.300 43.270 249.380 43.270 249.380 43.260 ;
        RECT 249.380 43.260 250.445 43.270 ;
        POLYGON 249.385 43.260 249.500 43.260 249.500 43.250 ;
        RECT 249.500 43.255 250.445 43.260 ;
        POLYGON 250.445 43.270 250.595 43.270 250.445 43.255 ;
        POLYGON 252.820 43.270 252.820 43.265 252.810 43.265 ;
        RECT 252.820 43.265 254.230 43.270 ;
        POLYGON 252.810 43.265 252.810 43.255 252.785 43.255 ;
        RECT 252.810 43.255 254.230 43.265 ;
        RECT 249.500 43.250 250.325 43.255 ;
        POLYGON 249.500 43.250 249.640 43.250 249.640 43.245 ;
        RECT 249.640 43.245 250.325 43.250 ;
        POLYGON 250.325 43.255 250.440 43.255 250.325 43.245 ;
        POLYGON 252.785 43.255 252.785 43.245 252.760 43.245 ;
        RECT 252.785 43.245 254.230 43.255 ;
        POLYGON 249.650 43.245 249.755 43.245 249.755 43.240 ;
        RECT 249.755 43.240 250.180 43.245 ;
        POLYGON 250.180 43.245 250.220 43.245 250.180 43.240 ;
        POLYGON 252.760 43.245 252.760 43.240 252.750 43.240 ;
        RECT 252.760 43.240 254.230 43.245 ;
        POLYGON 249.775 43.240 249.915 43.240 249.915 43.235 ;
        RECT 249.915 43.235 250.050 43.240 ;
        POLYGON 250.050 43.240 250.175 43.240 250.050 43.235 ;
        POLYGON 252.750 43.240 252.750 43.235 252.740 43.235 ;
        RECT 252.750 43.235 254.230 43.240 ;
        POLYGON 254.230 43.340 254.380 43.340 254.230 43.235 ;
        POLYGON 255.610 43.340 255.610 43.240 255.495 43.240 ;
        RECT 255.610 43.240 256.755 43.340 ;
        POLYGON 255.495 43.240 255.495 43.235 255.490 43.235 ;
        RECT 255.495 43.235 256.755 43.240 ;
        POLYGON 252.740 43.235 252.740 43.215 252.700 43.215 ;
        RECT 252.740 43.230 254.220 43.235 ;
        POLYGON 254.220 43.235 254.230 43.235 254.220 43.230 ;
        POLYGON 255.490 43.235 255.490 43.230 255.485 43.230 ;
        RECT 255.490 43.230 256.755 43.235 ;
        RECT 252.740 43.215 254.135 43.230 ;
        POLYGON 252.700 43.215 252.700 43.210 252.680 43.210 ;
        RECT 252.700 43.210 254.135 43.215 ;
        POLYGON 252.680 43.210 252.680 43.170 252.585 43.170 ;
        RECT 252.680 43.170 254.135 43.210 ;
        POLYGON 254.135 43.230 254.220 43.230 254.135 43.170 ;
        POLYGON 255.485 43.230 255.485 43.200 255.455 43.200 ;
        RECT 255.485 43.200 256.755 43.230 ;
        POLYGON 255.455 43.200 255.455 43.170 255.420 43.170 ;
        RECT 255.455 43.170 256.755 43.200 ;
        RECT 245.570 43.165 246.985 43.170 ;
        POLYGON 246.985 43.170 247.000 43.165 246.985 43.165 ;
        POLYGON 252.585 43.170 252.585 43.165 252.575 43.165 ;
        RECT 252.585 43.165 254.015 43.170 ;
        RECT 245.570 43.160 247.000 43.165 ;
        RECT 242.490 43.155 244.015 43.160 ;
        POLYGON 244.015 43.160 244.020 43.155 244.015 43.155 ;
        POLYGON 245.570 43.160 245.580 43.160 245.580 43.155 ;
        RECT 245.580 43.155 247.000 43.160 ;
        RECT 242.490 43.085 244.020 43.155 ;
        POLYGON 244.020 43.155 244.100 43.085 244.020 43.085 ;
        POLYGON 245.580 43.155 245.660 43.155 245.660 43.110 ;
        RECT 245.660 43.130 247.000 43.155 ;
        POLYGON 247.000 43.165 247.075 43.130 247.000 43.130 ;
        POLYGON 252.575 43.165 252.575 43.145 252.525 43.145 ;
        RECT 252.575 43.145 254.015 43.165 ;
        POLYGON 252.525 43.145 252.525 43.140 252.510 43.140 ;
        RECT 252.525 43.140 254.015 43.145 ;
        POLYGON 252.510 43.140 252.510 43.130 252.490 43.130 ;
        RECT 252.510 43.130 254.015 43.140 ;
        RECT 245.660 43.110 247.075 43.130 ;
        POLYGON 245.660 43.110 245.700 43.110 245.700 43.085 ;
        RECT 245.700 43.085 247.075 43.110 ;
        RECT 242.490 43.070 244.100 43.085 ;
        RECT 238.320 43.065 240.600 43.070 ;
        POLYGON 238.320 43.065 238.605 43.065 238.605 42.650 ;
        RECT 238.605 43.020 240.600 43.065 ;
        POLYGON 240.600 43.070 240.640 43.020 240.600 43.020 ;
        POLYGON 242.490 43.070 242.540 43.070 242.540 43.020 ;
        RECT 242.540 43.020 244.100 43.070 ;
        RECT 238.605 42.890 240.640 43.020 ;
        POLYGON 240.640 43.020 240.755 42.890 240.640 42.890 ;
        POLYGON 242.540 43.020 242.585 43.020 242.585 42.980 ;
        RECT 242.585 42.980 244.100 43.020 ;
        POLYGON 242.585 42.980 242.675 42.980 242.675 42.890 ;
        RECT 242.675 42.975 244.100 42.980 ;
        POLYGON 244.100 43.085 244.220 42.975 244.100 42.975 ;
        POLYGON 245.700 43.085 245.815 43.085 245.815 43.015 ;
        RECT 245.815 43.065 247.075 43.085 ;
        POLYGON 247.075 43.130 247.235 43.065 247.075 43.065 ;
        POLYGON 252.490 43.130 252.490 43.105 252.435 43.105 ;
        RECT 252.490 43.105 254.015 43.130 ;
        POLYGON 252.435 43.105 252.435 43.065 252.325 43.065 ;
        RECT 252.435 43.095 254.015 43.105 ;
        POLYGON 254.015 43.170 254.135 43.170 254.015 43.095 ;
        POLYGON 255.420 43.170 255.420 43.105 255.350 43.105 ;
        RECT 255.420 43.155 256.755 43.170 ;
        POLYGON 256.755 43.345 256.930 43.345 256.755 43.155 ;
        POLYGON 258.610 43.345 258.610 43.305 258.580 43.305 ;
        RECT 258.610 43.305 260.145 43.345 ;
        POLYGON 258.580 43.305 258.580 43.260 258.545 43.260 ;
        RECT 258.580 43.260 260.145 43.305 ;
        POLYGON 258.545 43.260 258.545 43.155 258.470 43.155 ;
        RECT 258.545 43.155 260.145 43.260 ;
        RECT 255.420 43.115 256.720 43.155 ;
        POLYGON 256.720 43.155 256.755 43.155 256.720 43.115 ;
        POLYGON 258.470 43.155 258.470 43.120 258.445 43.120 ;
        RECT 258.470 43.120 260.145 43.155 ;
        POLYGON 258.445 43.120 258.445 43.115 258.440 43.115 ;
        RECT 258.445 43.115 260.145 43.120 ;
        RECT 255.420 43.105 256.515 43.115 ;
        POLYGON 255.350 43.105 255.350 43.095 255.340 43.095 ;
        RECT 255.350 43.095 256.515 43.105 ;
        RECT 252.435 43.065 253.900 43.095 ;
        RECT 245.815 43.060 247.235 43.065 ;
        POLYGON 247.235 43.065 247.250 43.060 247.235 43.060 ;
        POLYGON 252.325 43.065 252.325 43.060 252.310 43.060 ;
        RECT 252.325 43.060 253.900 43.065 ;
        RECT 245.815 43.050 247.250 43.060 ;
        POLYGON 247.250 43.060 247.275 43.050 247.250 43.050 ;
        POLYGON 252.310 43.060 252.310 43.050 252.285 43.050 ;
        RECT 252.310 43.050 253.900 43.060 ;
        RECT 245.815 43.015 247.275 43.050 ;
        POLYGON 245.815 43.015 245.840 43.015 245.840 43.000 ;
        RECT 245.840 43.000 247.275 43.015 ;
        POLYGON 245.840 43.000 245.885 43.000 245.885 42.975 ;
        RECT 245.885 42.975 247.275 43.000 ;
        RECT 242.675 42.890 244.220 42.975 ;
        RECT 238.605 42.800 240.755 42.890 ;
        POLYGON 240.755 42.890 240.830 42.800 240.755 42.800 ;
        POLYGON 242.675 42.890 242.765 42.890 242.765 42.800 ;
        RECT 242.765 42.880 244.220 42.890 ;
        POLYGON 244.220 42.975 244.340 42.880 244.220 42.880 ;
        POLYGON 245.885 42.975 245.945 42.975 245.945 42.945 ;
        RECT 245.945 42.970 247.275 42.975 ;
        POLYGON 247.275 43.050 247.480 42.970 247.275 42.970 ;
        POLYGON 252.285 43.050 252.285 43.010 252.165 43.010 ;
        RECT 252.285 43.025 253.900 43.050 ;
        POLYGON 253.900 43.095 254.015 43.095 253.900 43.025 ;
        POLYGON 255.340 43.095 255.340 43.055 255.290 43.055 ;
        RECT 255.340 43.055 256.515 43.095 ;
        POLYGON 255.290 43.055 255.290 43.025 255.255 43.025 ;
        RECT 255.290 43.025 256.515 43.055 ;
        RECT 252.285 43.015 253.880 43.025 ;
        POLYGON 253.880 43.025 253.900 43.025 253.880 43.015 ;
        POLYGON 255.255 43.025 255.255 43.015 255.240 43.015 ;
        RECT 255.255 43.015 256.515 43.025 ;
        RECT 252.285 43.010 253.800 43.015 ;
        POLYGON 252.165 43.010 252.165 42.975 252.065 42.975 ;
        RECT 252.165 42.975 253.800 43.010 ;
        POLYGON 252.065 42.975 252.065 42.970 252.050 42.970 ;
        RECT 252.065 42.970 253.800 42.975 ;
        RECT 245.945 42.965 247.480 42.970 ;
        POLYGON 247.480 42.970 247.505 42.965 247.480 42.965 ;
        POLYGON 252.050 42.970 252.050 42.965 252.035 42.965 ;
        RECT 252.050 42.965 253.800 42.970 ;
        POLYGON 253.800 43.015 253.880 43.015 253.800 42.965 ;
        POLYGON 255.240 43.015 255.240 42.965 255.185 42.965 ;
        RECT 255.240 42.965 256.515 43.015 ;
        RECT 245.945 42.960 247.510 42.965 ;
        POLYGON 247.510 42.965 247.515 42.960 247.510 42.960 ;
        POLYGON 252.035 42.965 252.035 42.960 252.015 42.960 ;
        RECT 252.035 42.960 253.620 42.965 ;
        RECT 245.945 42.950 247.515 42.960 ;
        POLYGON 247.515 42.960 247.555 42.950 247.515 42.950 ;
        POLYGON 252.015 42.960 252.015 42.950 251.985 42.950 ;
        RECT 252.015 42.950 253.620 42.960 ;
        RECT 245.945 42.945 247.555 42.950 ;
        POLYGON 245.945 42.945 246.065 42.945 246.065 42.880 ;
        RECT 246.065 42.890 247.555 42.945 ;
        POLYGON 247.555 42.950 247.730 42.890 247.555 42.890 ;
        POLYGON 251.985 42.950 251.985 42.925 251.920 42.925 ;
        RECT 251.985 42.925 253.620 42.950 ;
        POLYGON 251.920 42.925 251.920 42.920 251.900 42.920 ;
        RECT 251.920 42.920 253.620 42.925 ;
        POLYGON 251.900 42.920 251.900 42.890 251.795 42.890 ;
        RECT 251.900 42.890 253.620 42.920 ;
        RECT 246.065 42.880 247.730 42.890 ;
        RECT 242.765 42.870 244.340 42.880 ;
        POLYGON 244.340 42.880 244.350 42.870 244.340 42.870 ;
        POLYGON 246.065 42.880 246.085 42.880 246.085 42.870 ;
        RECT 246.085 42.875 247.730 42.880 ;
        POLYGON 247.730 42.890 247.785 42.875 247.730 42.875 ;
        POLYGON 251.795 42.890 251.795 42.875 251.745 42.875 ;
        RECT 251.795 42.875 253.620 42.890 ;
        RECT 246.085 42.870 247.785 42.875 ;
        RECT 242.765 42.810 244.350 42.870 ;
        POLYGON 244.350 42.870 244.425 42.810 244.350 42.810 ;
        POLYGON 246.085 42.870 246.200 42.870 246.200 42.810 ;
        RECT 246.200 42.860 247.785 42.870 ;
        POLYGON 247.785 42.875 247.830 42.860 247.785 42.860 ;
        POLYGON 251.745 42.875 251.745 42.860 251.695 42.860 ;
        RECT 251.745 42.865 253.620 42.875 ;
        POLYGON 253.620 42.965 253.800 42.965 253.620 42.865 ;
        POLYGON 255.185 42.965 255.185 42.950 255.165 42.950 ;
        RECT 255.185 42.950 256.515 42.965 ;
        POLYGON 255.165 42.950 255.165 42.875 255.070 42.875 ;
        RECT 255.165 42.910 256.515 42.950 ;
        POLYGON 256.515 43.115 256.720 43.115 256.515 42.910 ;
        POLYGON 258.440 43.115 258.440 43.075 258.410 43.075 ;
        RECT 258.440 43.075 260.145 43.115 ;
        POLYGON 258.410 43.075 258.410 42.935 258.295 42.935 ;
        RECT 258.410 42.975 260.145 43.075 ;
        POLYGON 260.145 43.365 260.385 43.365 260.145 42.975 ;
        POLYGON 262.835 43.360 262.835 43.315 262.815 43.315 ;
        RECT 262.835 43.315 265.705 43.365 ;
        POLYGON 262.815 43.315 262.815 43.215 262.770 43.215 ;
        RECT 262.815 43.215 265.705 43.315 ;
        POLYGON 262.770 43.215 262.770 43.000 262.675 43.000 ;
        RECT 262.770 43.000 265.705 43.215 ;
        POLYGON 262.675 43.000 262.675 42.980 262.665 42.980 ;
        RECT 262.675 42.980 265.705 43.000 ;
        RECT 258.410 42.950 260.130 42.975 ;
        POLYGON 260.130 42.975 260.145 42.975 260.130 42.950 ;
        POLYGON 262.665 42.975 262.665 42.950 262.650 42.950 ;
        RECT 262.665 42.950 265.705 42.980 ;
        RECT 258.410 42.935 259.820 42.950 ;
        POLYGON 258.295 42.935 258.295 42.910 258.275 42.910 ;
        RECT 258.295 42.910 259.820 42.935 ;
        RECT 255.165 42.875 256.265 42.910 ;
        POLYGON 255.070 42.875 255.070 42.865 255.060 42.865 ;
        RECT 255.070 42.865 256.265 42.875 ;
        RECT 251.745 42.860 253.580 42.865 ;
        RECT 246.200 42.825 247.830 42.860 ;
        POLYGON 247.830 42.860 247.945 42.825 247.830 42.825 ;
        POLYGON 251.695 42.860 251.695 42.850 251.660 42.850 ;
        RECT 251.695 42.850 253.580 42.860 ;
        POLYGON 251.660 42.850 251.660 42.840 251.635 42.840 ;
        RECT 251.660 42.845 253.580 42.850 ;
        POLYGON 253.580 42.865 253.620 42.865 253.580 42.845 ;
        POLYGON 255.060 42.865 255.060 42.845 255.035 42.845 ;
        RECT 255.060 42.845 256.265 42.865 ;
        RECT 251.660 42.840 253.420 42.845 ;
        POLYGON 251.635 42.840 251.635 42.835 251.605 42.835 ;
        RECT 251.635 42.835 253.420 42.840 ;
        POLYGON 251.605 42.835 251.605 42.825 251.565 42.825 ;
        RECT 251.605 42.825 253.420 42.835 ;
        RECT 246.200 42.815 247.945 42.825 ;
        POLYGON 247.945 42.825 247.985 42.815 247.945 42.815 ;
        POLYGON 251.565 42.825 251.565 42.815 251.525 42.815 ;
        RECT 251.565 42.815 253.420 42.825 ;
        RECT 246.200 42.810 247.985 42.815 ;
        RECT 242.765 42.800 244.425 42.810 ;
        RECT 238.605 42.705 240.830 42.800 ;
        POLYGON 240.830 42.800 240.915 42.705 240.830 42.705 ;
        POLYGON 242.765 42.800 242.840 42.800 242.840 42.730 ;
        RECT 242.840 42.730 244.425 42.800 ;
        POLYGON 242.840 42.730 242.865 42.730 242.865 42.705 ;
        RECT 242.865 42.710 244.425 42.730 ;
        POLYGON 244.425 42.810 244.545 42.710 244.425 42.710 ;
        POLYGON 246.200 42.810 246.240 42.810 246.240 42.790 ;
        RECT 246.240 42.800 247.985 42.810 ;
        POLYGON 247.985 42.815 248.050 42.800 247.985 42.800 ;
        POLYGON 251.525 42.815 251.525 42.805 251.485 42.805 ;
        RECT 251.525 42.805 253.420 42.815 ;
        POLYGON 251.485 42.805 251.485 42.800 251.470 42.800 ;
        RECT 251.485 42.800 253.420 42.805 ;
        RECT 246.240 42.790 248.050 42.800 ;
        POLYGON 246.240 42.790 246.310 42.790 246.310 42.760 ;
        RECT 246.310 42.785 248.050 42.790 ;
        POLYGON 248.050 42.800 248.105 42.785 248.050 42.785 ;
        POLYGON 251.470 42.800 251.470 42.785 251.415 42.785 ;
        RECT 251.470 42.785 253.420 42.800 ;
        RECT 246.310 42.760 248.110 42.785 ;
        POLYGON 246.310 42.760 246.410 42.760 246.410 42.710 ;
        RECT 246.410 42.750 248.110 42.760 ;
        POLYGON 248.110 42.785 248.235 42.750 248.110 42.750 ;
        POLYGON 251.415 42.785 251.415 42.780 251.400 42.780 ;
        RECT 251.415 42.780 253.420 42.785 ;
        POLYGON 251.400 42.780 251.400 42.775 251.370 42.775 ;
        RECT 251.400 42.775 253.420 42.780 ;
        POLYGON 251.370 42.775 251.370 42.750 251.250 42.750 ;
        RECT 251.370 42.760 253.420 42.775 ;
        POLYGON 253.420 42.845 253.580 42.845 253.420 42.760 ;
        POLYGON 255.035 42.845 255.035 42.760 254.925 42.760 ;
        RECT 255.035 42.760 256.265 42.845 ;
        RECT 251.370 42.750 253.355 42.760 ;
        RECT 246.410 42.735 248.235 42.750 ;
        POLYGON 248.235 42.750 248.320 42.735 248.235 42.735 ;
        POLYGON 251.250 42.750 251.250 42.745 251.225 42.745 ;
        RECT 251.250 42.745 253.355 42.750 ;
        POLYGON 251.225 42.745 251.225 42.735 251.185 42.735 ;
        RECT 251.225 42.735 253.355 42.745 ;
        RECT 246.410 42.720 248.320 42.735 ;
        POLYGON 248.320 42.735 248.385 42.720 248.320 42.720 ;
        POLYGON 251.185 42.735 251.185 42.725 251.145 42.725 ;
        RECT 251.185 42.725 253.355 42.735 ;
        POLYGON 253.355 42.760 253.420 42.760 253.355 42.725 ;
        POLYGON 254.925 42.760 254.925 42.725 254.880 42.725 ;
        RECT 254.925 42.725 256.265 42.760 ;
        POLYGON 251.135 42.725 251.135 42.720 251.120 42.720 ;
        RECT 251.135 42.720 253.085 42.725 ;
        RECT 246.410 42.710 248.390 42.720 ;
        RECT 242.865 42.705 244.545 42.710 ;
        RECT 238.605 42.650 240.915 42.705 ;
        POLYGON 238.605 42.650 238.640 42.650 238.640 42.600 ;
        RECT 238.640 42.620 240.915 42.650 ;
        POLYGON 240.915 42.705 240.990 42.620 240.915 42.620 ;
        POLYGON 242.865 42.705 242.885 42.705 242.885 42.685 ;
        RECT 242.885 42.685 244.545 42.705 ;
        POLYGON 242.885 42.685 242.955 42.685 242.955 42.620 ;
        RECT 242.955 42.680 244.545 42.685 ;
        POLYGON 244.545 42.710 244.590 42.680 244.545 42.680 ;
        POLYGON 246.410 42.710 246.475 42.710 246.475 42.680 ;
        RECT 246.475 42.695 248.390 42.710 ;
        POLYGON 248.390 42.720 248.490 42.695 248.390 42.695 ;
        POLYGON 251.120 42.720 251.120 42.715 251.100 42.715 ;
        RECT 251.120 42.715 253.085 42.720 ;
        POLYGON 251.100 42.715 251.100 42.695 250.990 42.695 ;
        RECT 251.100 42.695 253.085 42.715 ;
        RECT 246.475 42.680 248.490 42.695 ;
        POLYGON 248.490 42.695 248.585 42.680 248.490 42.680 ;
        POLYGON 250.990 42.695 250.990 42.690 250.965 42.690 ;
        RECT 250.990 42.690 253.085 42.695 ;
        POLYGON 250.965 42.690 250.965 42.680 250.900 42.680 ;
        RECT 250.965 42.680 253.085 42.690 ;
        RECT 242.955 42.620 244.590 42.680 ;
        RECT 238.640 42.605 240.990 42.620 ;
        POLYGON 240.990 42.620 241.005 42.605 240.990 42.605 ;
        POLYGON 242.955 42.620 242.975 42.620 242.975 42.605 ;
        RECT 242.975 42.605 244.590 42.620 ;
        RECT 238.640 42.600 241.005 42.605 ;
        POLYGON 238.640 42.600 238.695 42.600 238.695 42.525 ;
        RECT 238.695 42.525 241.005 42.600 ;
        RECT 231.245 42.485 235.575 42.525 ;
        POLYGON 235.575 42.525 235.595 42.485 235.575 42.485 ;
        POLYGON 238.695 42.525 238.730 42.525 238.730 42.485 ;
        RECT 238.730 42.515 241.005 42.525 ;
        POLYGON 241.005 42.605 241.090 42.515 241.005 42.515 ;
        POLYGON 242.975 42.605 243.075 42.605 243.075 42.515 ;
        RECT 243.075 42.590 244.590 42.605 ;
        POLYGON 244.590 42.680 244.700 42.590 244.590 42.590 ;
        POLYGON 246.475 42.680 246.540 42.680 246.540 42.650 ;
        RECT 246.540 42.665 248.585 42.680 ;
        POLYGON 248.585 42.680 248.665 42.665 248.585 42.665 ;
        POLYGON 250.900 42.680 250.900 42.675 250.865 42.675 ;
        RECT 250.900 42.675 253.085 42.680 ;
        POLYGON 250.865 42.675 250.865 42.670 250.840 42.670 ;
        RECT 250.865 42.670 253.085 42.675 ;
        POLYGON 250.840 42.670 250.840 42.665 250.805 42.665 ;
        RECT 250.840 42.665 253.085 42.670 ;
        RECT 246.540 42.655 248.665 42.665 ;
        POLYGON 248.665 42.665 248.750 42.655 248.665 42.655 ;
        POLYGON 250.805 42.665 250.805 42.655 250.740 42.655 ;
        RECT 250.805 42.655 253.085 42.665 ;
        RECT 246.540 42.650 248.750 42.655 ;
        POLYGON 246.545 42.650 246.655 42.650 246.655 42.600 ;
        RECT 246.655 42.640 248.750 42.650 ;
        POLYGON 248.750 42.655 248.840 42.640 248.750 42.640 ;
        POLYGON 250.740 42.655 250.740 42.650 250.705 42.650 ;
        RECT 250.740 42.650 253.085 42.655 ;
        POLYGON 250.700 42.650 250.700 42.645 250.680 42.645 ;
        RECT 250.700 42.645 253.085 42.650 ;
        POLYGON 250.675 42.645 250.675 42.640 250.635 42.640 ;
        RECT 250.675 42.640 253.085 42.645 ;
        RECT 246.655 42.630 248.850 42.640 ;
        POLYGON 248.850 42.640 248.945 42.630 248.850 42.630 ;
        POLYGON 250.635 42.640 250.635 42.635 250.595 42.635 ;
        RECT 250.635 42.635 253.085 42.640 ;
        POLYGON 250.595 42.635 250.595 42.630 250.575 42.630 ;
        RECT 250.595 42.630 253.085 42.635 ;
        RECT 246.655 42.620 248.945 42.630 ;
        POLYGON 248.945 42.630 249.005 42.620 248.945 42.620 ;
        POLYGON 250.575 42.630 250.575 42.620 250.445 42.620 ;
        RECT 250.575 42.620 253.085 42.630 ;
        RECT 246.655 42.610 249.005 42.620 ;
        POLYGON 249.005 42.620 249.115 42.610 249.005 42.610 ;
        POLYGON 250.440 42.620 250.440 42.610 250.365 42.610 ;
        RECT 250.440 42.610 253.085 42.620 ;
        RECT 246.655 42.600 249.120 42.610 ;
        POLYGON 249.120 42.610 249.220 42.600 249.120 42.600 ;
        POLYGON 250.365 42.610 250.365 42.605 250.330 42.605 ;
        RECT 250.365 42.605 253.085 42.610 ;
        POLYGON 250.310 42.605 250.310 42.600 250.220 42.600 ;
        RECT 250.310 42.600 253.085 42.605 ;
        POLYGON 253.085 42.725 253.355 42.725 253.085 42.600 ;
        POLYGON 254.880 42.725 254.880 42.715 254.865 42.715 ;
        RECT 254.880 42.715 256.265 42.725 ;
        POLYGON 254.860 42.715 254.860 42.705 254.850 42.705 ;
        RECT 254.860 42.705 256.265 42.715 ;
        POLYGON 254.850 42.705 254.850 42.650 254.775 42.650 ;
        RECT 254.850 42.670 256.265 42.705 ;
        POLYGON 256.265 42.910 256.515 42.910 256.265 42.670 ;
        POLYGON 258.275 42.910 258.275 42.875 258.245 42.875 ;
        RECT 258.275 42.875 259.820 42.910 ;
        POLYGON 258.245 42.875 258.245 42.740 258.140 42.740 ;
        RECT 258.245 42.740 259.820 42.875 ;
        POLYGON 258.140 42.740 258.140 42.725 258.130 42.725 ;
        RECT 258.140 42.725 259.820 42.740 ;
        POLYGON 258.130 42.725 258.130 42.670 258.080 42.670 ;
        RECT 258.130 42.670 259.820 42.725 ;
        RECT 254.850 42.660 256.255 42.670 ;
        POLYGON 256.255 42.670 256.265 42.670 256.255 42.660 ;
        POLYGON 258.080 42.670 258.080 42.660 258.070 42.660 ;
        RECT 258.080 42.660 259.820 42.670 ;
        RECT 254.850 42.650 256.200 42.660 ;
        POLYGON 254.775 42.650 254.775 42.600 254.705 42.600 ;
        RECT 254.775 42.610 256.200 42.650 ;
        POLYGON 256.200 42.660 256.255 42.660 256.200 42.610 ;
        POLYGON 258.070 42.660 258.070 42.610 258.025 42.610 ;
        RECT 258.070 42.610 259.820 42.660 ;
        RECT 254.775 42.600 256.005 42.610 ;
        POLYGON 246.655 42.600 246.675 42.600 246.675 42.590 ;
        RECT 246.675 42.595 249.225 42.600 ;
        POLYGON 249.225 42.600 249.265 42.595 249.225 42.595 ;
        POLYGON 250.215 42.600 250.215 42.595 250.175 42.595 ;
        RECT 250.215 42.595 252.980 42.600 ;
        RECT 246.675 42.590 249.300 42.595 ;
        POLYGON 249.300 42.595 249.385 42.590 249.300 42.590 ;
        POLYGON 250.170 42.595 250.170 42.590 250.110 42.590 ;
        RECT 250.170 42.590 252.980 42.595 ;
        RECT 243.075 42.515 244.700 42.590 ;
        RECT 238.730 42.485 241.090 42.515 ;
        RECT 231.245 42.355 235.595 42.485 ;
        RECT 209.390 42.155 224.120 42.355 ;
        POLYGON 224.120 42.355 224.200 42.155 224.120 42.155 ;
        POLYGON 231.245 42.355 231.280 42.355 231.280 42.290 ;
        RECT 231.280 42.290 235.595 42.355 ;
        POLYGON 231.280 42.290 231.345 42.290 231.345 42.160 ;
        RECT 231.345 42.220 235.595 42.290 ;
        POLYGON 235.595 42.485 235.765 42.220 235.595 42.220 ;
        POLYGON 238.730 42.485 238.935 42.485 238.935 42.220 ;
        RECT 238.935 42.320 241.090 42.485 ;
        POLYGON 241.090 42.515 241.270 42.320 241.090 42.320 ;
        POLYGON 243.075 42.515 243.100 42.515 243.100 42.495 ;
        RECT 243.100 42.495 244.700 42.515 ;
        POLYGON 243.100 42.495 243.245 42.495 243.245 42.365 ;
        RECT 243.245 42.485 244.700 42.495 ;
        POLYGON 244.700 42.590 244.840 42.485 244.700 42.485 ;
        POLYGON 246.675 42.590 246.775 42.590 246.775 42.550 ;
        RECT 246.775 42.585 249.385 42.590 ;
        POLYGON 249.385 42.590 249.485 42.585 249.385 42.585 ;
        POLYGON 250.110 42.590 250.110 42.585 250.045 42.585 ;
        RECT 250.110 42.585 252.980 42.590 ;
        RECT 246.775 42.580 249.525 42.585 ;
        POLYGON 249.525 42.585 249.610 42.580 249.525 42.580 ;
        POLYGON 249.895 42.585 249.895 42.580 249.785 42.580 ;
        RECT 249.895 42.580 252.980 42.585 ;
        RECT 246.775 42.550 252.980 42.580 ;
        POLYGON 252.980 42.600 253.085 42.600 252.980 42.550 ;
        POLYGON 254.705 42.600 254.705 42.550 254.635 42.550 ;
        RECT 254.705 42.550 256.005 42.600 ;
        POLYGON 246.775 42.550 246.930 42.550 246.930 42.485 ;
        RECT 246.930 42.515 252.895 42.550 ;
        POLYGON 252.895 42.550 252.975 42.550 252.895 42.515 ;
        POLYGON 254.635 42.550 254.635 42.535 254.615 42.535 ;
        RECT 254.635 42.535 256.005 42.550 ;
        POLYGON 254.615 42.535 254.615 42.515 254.585 42.515 ;
        RECT 254.615 42.515 256.005 42.535 ;
        RECT 246.930 42.485 252.810 42.515 ;
        RECT 243.245 42.465 244.845 42.485 ;
        POLYGON 244.845 42.485 244.870 42.465 244.845 42.465 ;
        POLYGON 246.930 42.485 246.970 42.485 246.970 42.470 ;
        RECT 246.970 42.480 252.810 42.485 ;
        POLYGON 252.810 42.515 252.895 42.515 252.810 42.480 ;
        POLYGON 254.585 42.515 254.585 42.490 254.550 42.490 ;
        RECT 254.585 42.490 256.005 42.515 ;
        POLYGON 254.550 42.490 254.550 42.480 254.540 42.480 ;
        RECT 254.550 42.480 256.005 42.490 ;
        RECT 246.970 42.470 252.760 42.480 ;
        POLYGON 246.970 42.470 246.980 42.470 246.980 42.465 ;
        RECT 246.980 42.465 252.760 42.470 ;
        RECT 243.245 42.365 244.870 42.465 ;
        POLYGON 243.245 42.365 243.300 42.365 243.300 42.320 ;
        RECT 243.300 42.330 244.870 42.365 ;
        POLYGON 244.870 42.465 245.065 42.330 244.870 42.330 ;
        POLYGON 246.980 42.465 247.005 42.465 247.005 42.455 ;
        RECT 247.005 42.460 252.760 42.465 ;
        POLYGON 252.760 42.480 252.810 42.480 252.760 42.460 ;
        POLYGON 254.540 42.480 254.540 42.460 254.510 42.460 ;
        RECT 254.540 42.460 256.005 42.480 ;
        RECT 247.005 42.455 252.545 42.460 ;
        POLYGON 247.010 42.455 247.075 42.455 247.075 42.430 ;
        RECT 247.075 42.430 252.545 42.455 ;
        POLYGON 247.075 42.430 247.195 42.430 247.195 42.390 ;
        RECT 247.195 42.390 252.545 42.430 ;
        POLYGON 247.195 42.390 247.245 42.390 247.245 42.375 ;
        RECT 247.245 42.380 252.545 42.390 ;
        POLYGON 252.545 42.460 252.760 42.460 252.545 42.380 ;
        POLYGON 254.510 42.460 254.510 42.435 254.475 42.435 ;
        RECT 254.510 42.435 256.005 42.460 ;
        POLYGON 256.005 42.610 256.200 42.610 256.005 42.435 ;
        POLYGON 258.025 42.610 258.025 42.595 258.010 42.595 ;
        RECT 258.025 42.595 259.820 42.610 ;
        POLYGON 258.010 42.595 258.010 42.550 257.975 42.550 ;
        RECT 258.010 42.550 259.820 42.595 ;
        POLYGON 257.975 42.550 257.975 42.510 257.935 42.510 ;
        RECT 257.975 42.510 259.820 42.550 ;
        POLYGON 257.935 42.510 257.935 42.435 257.865 42.435 ;
        RECT 257.935 42.490 259.820 42.510 ;
        POLYGON 259.820 42.950 260.130 42.950 259.820 42.490 ;
        POLYGON 262.650 42.945 262.650 42.820 262.590 42.820 ;
        RECT 262.650 42.935 265.705 42.950 ;
        POLYGON 265.705 43.365 265.850 43.365 265.705 42.935 ;
        POLYGON 270.460 43.365 270.460 43.290 270.445 43.290 ;
        RECT 270.460 43.290 277.650 43.375 ;
        POLYGON 270.445 43.290 270.445 43.055 270.390 43.055 ;
        RECT 270.445 43.055 277.650 43.290 ;
        POLYGON 270.390 43.055 270.390 42.990 270.375 42.990 ;
        RECT 270.390 42.990 277.650 43.055 ;
        POLYGON 270.375 42.990 270.375 42.935 270.360 42.935 ;
        RECT 270.375 42.935 277.650 42.990 ;
        RECT 262.650 42.820 265.490 42.935 ;
        POLYGON 262.590 42.820 262.590 42.490 262.430 42.490 ;
        RECT 262.590 42.490 265.490 42.820 ;
        RECT 257.935 42.435 259.655 42.490 ;
        POLYGON 254.475 42.435 254.475 42.380 254.390 42.380 ;
        RECT 254.475 42.380 255.815 42.435 ;
        RECT 247.245 42.375 252.525 42.380 ;
        POLYGON 247.245 42.375 247.365 42.375 247.365 42.330 ;
        RECT 247.365 42.370 252.525 42.375 ;
        POLYGON 252.525 42.380 252.545 42.380 252.525 42.370 ;
        POLYGON 254.390 42.380 254.390 42.370 254.370 42.370 ;
        RECT 254.390 42.370 255.815 42.380 ;
        RECT 247.365 42.335 252.415 42.370 ;
        POLYGON 252.415 42.370 252.525 42.370 252.415 42.335 ;
        POLYGON 254.370 42.370 254.370 42.335 254.315 42.335 ;
        RECT 254.370 42.335 255.815 42.370 ;
        RECT 247.365 42.330 252.325 42.335 ;
        RECT 243.300 42.320 245.065 42.330 ;
        RECT 238.935 42.230 241.270 42.320 ;
        POLYGON 241.270 42.320 241.355 42.230 241.270 42.230 ;
        POLYGON 243.300 42.320 243.375 42.320 243.375 42.260 ;
        RECT 243.375 42.300 245.065 42.320 ;
        POLYGON 245.065 42.330 245.110 42.300 245.065 42.300 ;
        POLYGON 247.365 42.330 247.455 42.330 247.455 42.300 ;
        RECT 247.455 42.305 252.325 42.330 ;
        POLYGON 252.325 42.335 252.415 42.335 252.325 42.305 ;
        POLYGON 254.315 42.335 254.315 42.305 254.270 42.305 ;
        RECT 254.315 42.305 255.815 42.335 ;
        RECT 247.455 42.300 252.100 42.305 ;
        RECT 243.375 42.260 245.110 42.300 ;
        POLYGON 243.375 42.260 243.410 42.260 243.410 42.230 ;
        RECT 243.410 42.245 245.110 42.260 ;
        POLYGON 245.110 42.300 245.190 42.245 245.110 42.245 ;
        POLYGON 247.455 42.300 247.485 42.300 247.485 42.290 ;
        RECT 247.485 42.290 252.100 42.300 ;
        POLYGON 247.485 42.290 247.510 42.290 247.510 42.285 ;
        RECT 247.510 42.285 252.100 42.290 ;
        POLYGON 247.510 42.285 247.650 42.285 247.650 42.245 ;
        RECT 247.650 42.245 252.100 42.285 ;
        RECT 243.410 42.230 245.190 42.245 ;
        RECT 238.935 42.220 241.355 42.230 ;
        RECT 231.345 42.155 235.765 42.220 ;
        RECT 209.390 41.940 224.200 42.155 ;
        POLYGON 224.200 42.155 224.295 41.940 224.200 41.940 ;
        POLYGON 231.345 42.155 231.350 42.155 231.350 42.150 ;
        RECT 231.350 42.150 235.765 42.155 ;
        POLYGON 231.350 42.150 231.460 42.150 231.460 41.940 ;
        RECT 231.460 41.940 235.765 42.150 ;
        RECT 209.390 41.770 224.295 41.940 ;
        POLYGON 224.295 41.940 224.375 41.770 224.295 41.770 ;
        POLYGON 231.460 41.940 231.550 41.940 231.550 41.770 ;
        RECT 231.550 41.895 235.765 41.940 ;
        POLYGON 235.765 42.220 235.975 41.895 235.765 41.895 ;
        POLYGON 238.935 42.220 238.965 42.220 238.965 42.185 ;
        RECT 238.965 42.185 241.355 42.220 ;
        POLYGON 238.965 42.185 239.125 42.185 239.125 41.985 ;
        RECT 239.125 42.125 241.355 42.185 ;
        POLYGON 241.355 42.230 241.465 42.125 241.355 42.125 ;
        POLYGON 243.410 42.230 243.545 42.230 243.545 42.125 ;
        RECT 243.545 42.200 245.190 42.230 ;
        POLYGON 245.190 42.245 245.265 42.200 245.190 42.200 ;
        POLYGON 247.650 42.245 247.740 42.245 247.740 42.220 ;
        RECT 247.740 42.235 252.100 42.245 ;
        POLYGON 252.100 42.305 252.325 42.305 252.100 42.235 ;
        POLYGON 254.270 42.305 254.270 42.280 254.230 42.280 ;
        RECT 254.270 42.280 255.815 42.305 ;
        POLYGON 255.815 42.435 256.005 42.435 255.815 42.280 ;
        POLYGON 257.865 42.435 257.865 42.355 257.795 42.355 ;
        RECT 257.865 42.355 259.655 42.435 ;
        POLYGON 257.795 42.350 257.795 42.280 257.725 42.280 ;
        RECT 257.795 42.280 259.655 42.355 ;
        POLYGON 254.230 42.280 254.230 42.275 254.220 42.275 ;
        RECT 254.230 42.275 255.735 42.280 ;
        POLYGON 254.220 42.275 254.220 42.240 254.165 42.240 ;
        RECT 254.220 42.240 255.735 42.275 ;
        POLYGON 254.165 42.240 254.165 42.235 254.160 42.235 ;
        RECT 254.165 42.235 255.735 42.240 ;
        RECT 247.740 42.225 252.065 42.235 ;
        POLYGON 252.065 42.235 252.095 42.235 252.065 42.225 ;
        POLYGON 254.160 42.235 254.160 42.225 254.145 42.225 ;
        RECT 254.160 42.225 255.735 42.235 ;
        RECT 247.740 42.220 251.925 42.225 ;
        POLYGON 247.740 42.220 247.805 42.220 247.805 42.200 ;
        RECT 247.805 42.200 251.925 42.220 ;
        RECT 243.545 42.125 245.265 42.200 ;
        POLYGON 245.265 42.200 245.380 42.125 245.265 42.125 ;
        POLYGON 247.805 42.200 247.895 42.200 247.895 42.175 ;
        RECT 247.895 42.185 251.925 42.200 ;
        POLYGON 251.925 42.225 252.065 42.225 251.925 42.185 ;
        POLYGON 254.145 42.225 254.145 42.220 254.135 42.220 ;
        RECT 254.145 42.220 255.735 42.225 ;
        POLYGON 254.130 42.220 254.130 42.185 254.075 42.185 ;
        RECT 254.130 42.210 255.735 42.220 ;
        POLYGON 255.735 42.280 255.815 42.280 255.735 42.210 ;
        POLYGON 257.725 42.280 257.725 42.210 257.660 42.210 ;
        RECT 257.725 42.260 259.655 42.280 ;
        POLYGON 259.655 42.490 259.820 42.490 259.655 42.260 ;
        POLYGON 262.430 42.490 262.430 42.450 262.405 42.450 ;
        RECT 262.430 42.450 265.490 42.490 ;
        POLYGON 262.405 42.450 262.405 42.335 262.345 42.335 ;
        RECT 262.405 42.370 265.490 42.450 ;
        POLYGON 265.490 42.935 265.705 42.935 265.490 42.370 ;
        POLYGON 270.360 42.930 270.360 42.735 270.310 42.735 ;
        RECT 270.360 42.840 277.650 42.935 ;
        POLYGON 277.650 44.075 277.780 44.075 277.650 42.840 ;
        POLYGON 287.780 44.095 287.780 42.840 287.715 42.840 ;
        RECT 287.780 42.840 303.120 44.110 ;
        RECT 270.360 42.735 277.455 42.840 ;
        POLYGON 270.310 42.735 270.310 42.690 270.295 42.690 ;
        RECT 270.310 42.690 277.455 42.735 ;
        POLYGON 270.295 42.690 270.295 42.370 270.195 42.370 ;
        RECT 270.295 42.370 277.455 42.690 ;
        RECT 262.405 42.335 265.455 42.370 ;
        POLYGON 262.345 42.335 262.345 42.260 262.300 42.260 ;
        RECT 262.345 42.295 265.455 42.335 ;
        POLYGON 265.455 42.370 265.490 42.370 265.455 42.295 ;
        POLYGON 270.195 42.365 270.195 42.300 270.175 42.300 ;
        RECT 270.195 42.300 277.455 42.370 ;
        RECT 262.345 42.260 265.255 42.295 ;
        RECT 257.725 42.210 259.495 42.260 ;
        RECT 254.130 42.185 255.455 42.210 ;
        RECT 247.895 42.175 251.860 42.185 ;
        POLYGON 247.895 42.175 247.945 42.175 247.945 42.160 ;
        RECT 247.945 42.170 251.860 42.175 ;
        POLYGON 251.860 42.185 251.920 42.185 251.860 42.170 ;
        POLYGON 254.075 42.185 254.075 42.170 254.050 42.170 ;
        RECT 254.075 42.170 255.455 42.185 ;
        RECT 247.945 42.160 251.615 42.170 ;
        POLYGON 247.945 42.160 248.005 42.160 248.005 42.150 ;
        RECT 248.005 42.150 251.615 42.160 ;
        POLYGON 248.010 42.150 248.115 42.150 248.115 42.125 ;
        RECT 248.115 42.125 251.615 42.150 ;
        RECT 239.125 42.030 241.465 42.125 ;
        POLYGON 241.465 42.125 241.560 42.030 241.465 42.030 ;
        POLYGON 243.545 42.125 243.630 42.125 243.630 42.060 ;
        RECT 243.630 42.060 245.380 42.125 ;
        POLYGON 243.630 42.060 243.645 42.060 243.645 42.050 ;
        RECT 243.645 42.050 245.380 42.060 ;
        POLYGON 243.645 42.050 243.665 42.050 243.665 42.030 ;
        RECT 243.665 42.045 245.380 42.050 ;
        POLYGON 245.380 42.125 245.510 42.045 245.380 42.045 ;
        POLYGON 248.115 42.125 248.295 42.125 248.295 42.085 ;
        RECT 248.295 42.110 251.615 42.125 ;
        POLYGON 251.615 42.170 251.860 42.170 251.615 42.110 ;
        POLYGON 254.050 42.170 254.050 42.110 253.945 42.110 ;
        RECT 254.050 42.110 255.455 42.170 ;
        RECT 248.295 42.105 251.605 42.110 ;
        POLYGON 251.605 42.110 251.615 42.110 251.605 42.105 ;
        POLYGON 253.945 42.110 253.945 42.105 253.935 42.105 ;
        RECT 253.945 42.105 255.455 42.110 ;
        RECT 248.295 42.085 251.425 42.105 ;
        POLYGON 248.295 42.085 248.315 42.085 248.315 42.080 ;
        RECT 248.315 42.080 251.425 42.085 ;
        POLYGON 248.315 42.080 248.380 42.080 248.380 42.065 ;
        RECT 248.380 42.070 251.425 42.080 ;
        POLYGON 251.425 42.105 251.605 42.105 251.425 42.070 ;
        POLYGON 253.935 42.105 253.935 42.085 253.900 42.085 ;
        RECT 253.935 42.085 255.455 42.105 ;
        POLYGON 253.900 42.085 253.900 42.075 253.880 42.075 ;
        RECT 253.900 42.075 255.455 42.085 ;
        POLYGON 253.880 42.075 253.880 42.070 253.875 42.070 ;
        RECT 253.880 42.070 255.455 42.075 ;
        RECT 248.380 42.065 251.350 42.070 ;
        POLYGON 248.390 42.065 248.510 42.065 248.510 42.045 ;
        RECT 248.510 42.055 251.350 42.065 ;
        POLYGON 251.350 42.070 251.425 42.070 251.350 42.055 ;
        POLYGON 253.875 42.070 253.875 42.055 253.850 42.055 ;
        RECT 253.875 42.055 255.455 42.070 ;
        RECT 248.510 42.045 251.145 42.055 ;
        RECT 243.665 42.030 245.510 42.045 ;
        RECT 239.125 41.985 241.560 42.030 ;
        POLYGON 239.125 41.985 239.130 41.985 239.130 41.980 ;
        RECT 239.130 41.980 241.560 41.985 ;
        POLYGON 239.130 41.980 239.200 41.980 239.200 41.900 ;
        RECT 239.200 41.925 241.560 41.980 ;
        POLYGON 241.560 42.030 241.670 41.925 241.560 41.925 ;
        POLYGON 243.665 42.030 243.810 42.030 243.810 41.925 ;
        RECT 243.810 41.960 245.510 42.030 ;
        POLYGON 245.510 42.045 245.660 41.960 245.510 41.960 ;
        POLYGON 248.510 42.045 248.845 42.045 248.845 41.990 ;
        RECT 248.845 42.015 251.145 42.045 ;
        POLYGON 251.145 42.055 251.345 42.055 251.145 42.015 ;
        POLYGON 253.850 42.055 253.850 42.050 253.845 42.050 ;
        RECT 253.850 42.050 255.455 42.055 ;
        POLYGON 253.845 42.050 253.845 42.030 253.800 42.030 ;
        RECT 253.845 42.030 255.455 42.050 ;
        POLYGON 253.800 42.030 253.800 42.015 253.770 42.015 ;
        RECT 253.800 42.015 255.455 42.030 ;
        RECT 248.845 42.005 251.065 42.015 ;
        POLYGON 251.065 42.015 251.145 42.015 251.065 42.005 ;
        POLYGON 253.770 42.015 253.770 42.005 253.755 42.005 ;
        RECT 253.770 42.005 255.455 42.015 ;
        RECT 248.845 41.990 250.915 42.005 ;
        POLYGON 248.845 41.990 248.870 41.990 248.870 41.985 ;
        RECT 248.870 41.985 250.915 41.990 ;
        POLYGON 250.915 42.005 251.065 42.005 250.915 41.985 ;
        POLYGON 253.755 42.005 253.755 41.985 253.715 41.985 ;
        RECT 253.755 41.990 255.455 42.005 ;
        POLYGON 255.455 42.210 255.735 42.210 255.455 41.990 ;
        POLYGON 257.660 42.210 257.660 42.160 257.610 42.160 ;
        RECT 257.660 42.160 259.495 42.210 ;
        POLYGON 257.610 42.160 257.610 42.150 257.595 42.150 ;
        RECT 257.610 42.150 259.495 42.160 ;
        POLYGON 257.595 42.150 257.595 41.990 257.440 41.990 ;
        RECT 257.595 42.040 259.495 42.150 ;
        POLYGON 259.495 42.260 259.655 42.260 259.495 42.040 ;
        POLYGON 262.300 42.255 262.300 42.150 262.240 42.150 ;
        RECT 262.300 42.150 265.255 42.260 ;
        POLYGON 262.240 42.150 262.240 42.040 262.170 42.040 ;
        RECT 262.240 42.040 265.255 42.150 ;
        RECT 257.595 41.990 259.210 42.040 ;
        RECT 253.755 41.985 255.280 41.990 ;
        POLYGON 248.875 41.985 248.940 41.985 248.940 41.980 ;
        RECT 248.940 41.980 250.680 41.985 ;
        POLYGON 248.940 41.980 248.955 41.980 248.955 41.975 ;
        RECT 248.955 41.975 250.680 41.980 ;
        POLYGON 248.965 41.975 249.105 41.975 249.105 41.960 ;
        RECT 249.105 41.960 250.680 41.975 ;
        RECT 243.810 41.955 245.660 41.960 ;
        POLYGON 245.660 41.960 245.665 41.955 245.660 41.955 ;
        POLYGON 249.105 41.960 249.155 41.960 249.155 41.955 ;
        RECT 249.155 41.955 250.680 41.960 ;
        POLYGON 250.680 41.985 250.910 41.985 250.680 41.955 ;
        POLYGON 253.715 41.985 253.715 41.955 253.660 41.955 ;
        RECT 253.715 41.955 255.280 41.985 ;
        RECT 243.810 41.925 245.665 41.955 ;
        RECT 239.200 41.895 241.670 41.925 ;
        RECT 231.550 41.875 235.975 41.895 ;
        POLYGON 235.975 41.895 235.985 41.875 235.975 41.875 ;
        POLYGON 239.200 41.895 239.220 41.895 239.220 41.875 ;
        RECT 239.220 41.875 241.670 41.895 ;
        RECT 231.550 41.845 235.985 41.875 ;
        POLYGON 235.985 41.875 236.005 41.845 235.985 41.845 ;
        POLYGON 239.220 41.875 239.245 41.875 239.245 41.845 ;
        RECT 239.245 41.855 241.670 41.875 ;
        POLYGON 241.670 41.925 241.740 41.855 241.670 41.855 ;
        POLYGON 243.810 41.925 243.905 41.925 243.905 41.855 ;
        RECT 243.905 41.880 245.665 41.925 ;
        POLYGON 245.665 41.955 245.815 41.880 245.665 41.880 ;
        POLYGON 249.155 41.955 249.300 41.955 249.300 41.940 ;
        RECT 249.300 41.940 250.435 41.955 ;
        POLYGON 250.435 41.955 250.680 41.955 250.435 41.940 ;
        POLYGON 253.660 41.955 253.660 41.940 253.630 41.940 ;
        RECT 253.660 41.940 255.280 41.955 ;
        POLYGON 249.300 41.940 249.380 41.940 249.380 41.935 ;
        RECT 249.380 41.935 250.405 41.940 ;
        POLYGON 250.405 41.940 250.430 41.940 250.405 41.935 ;
        POLYGON 253.630 41.940 253.630 41.935 253.620 41.935 ;
        RECT 253.630 41.935 255.280 41.940 ;
        POLYGON 249.380 41.935 249.695 41.935 249.695 41.920 ;
        RECT 249.695 41.925 250.220 41.935 ;
        POLYGON 250.220 41.935 250.400 41.935 250.220 41.925 ;
        POLYGON 253.620 41.935 253.620 41.925 253.605 41.925 ;
        RECT 253.620 41.925 255.280 41.935 ;
        RECT 249.695 41.920 249.890 41.925 ;
        POLYGON 249.890 41.925 250.220 41.925 249.890 41.920 ;
        POLYGON 253.605 41.925 253.605 41.920 253.595 41.920 ;
        RECT 253.605 41.920 255.280 41.925 ;
        POLYGON 253.595 41.920 253.595 41.910 253.580 41.910 ;
        RECT 253.595 41.910 255.280 41.920 ;
        POLYGON 253.580 41.910 253.580 41.880 253.515 41.880 ;
        RECT 253.580 41.880 255.280 41.910 ;
        RECT 243.905 41.875 245.815 41.880 ;
        POLYGON 245.815 41.880 245.820 41.875 245.815 41.875 ;
        POLYGON 253.515 41.880 253.515 41.875 253.505 41.875 ;
        RECT 253.515 41.875 255.280 41.880 ;
        RECT 243.905 41.865 245.820 41.875 ;
        POLYGON 245.820 41.875 245.840 41.865 245.820 41.865 ;
        POLYGON 253.505 41.875 253.505 41.865 253.485 41.865 ;
        RECT 253.505 41.865 255.280 41.875 ;
        POLYGON 255.280 41.990 255.455 41.990 255.280 41.865 ;
        POLYGON 257.440 41.990 257.440 41.960 257.410 41.960 ;
        RECT 257.440 41.960 259.210 41.990 ;
        POLYGON 257.410 41.960 257.410 41.865 257.305 41.865 ;
        RECT 257.410 41.865 259.210 41.960 ;
        RECT 243.905 41.855 245.840 41.865 ;
        RECT 239.245 41.845 241.740 41.855 ;
        RECT 231.550 41.790 236.005 41.845 ;
        POLYGON 236.005 41.845 236.040 41.790 236.005 41.790 ;
        POLYGON 239.245 41.845 239.295 41.845 239.295 41.790 ;
        RECT 239.295 41.790 241.740 41.845 ;
        RECT 231.550 41.785 236.040 41.790 ;
        POLYGON 236.040 41.790 236.045 41.785 236.040 41.785 ;
        POLYGON 239.295 41.790 239.300 41.790 239.300 41.785 ;
        RECT 239.300 41.785 241.740 41.790 ;
        RECT 231.550 41.770 236.045 41.785 ;
        RECT 209.390 41.645 224.375 41.770 ;
        POLYGON 209.390 41.645 209.825 41.645 209.825 40.540 ;
        RECT 209.825 41.320 224.375 41.645 ;
        POLYGON 224.375 41.770 224.575 41.320 224.375 41.320 ;
        POLYGON 231.550 41.770 231.580 41.770 231.580 41.715 ;
        RECT 231.580 41.740 236.045 41.770 ;
        POLYGON 236.045 41.785 236.075 41.740 236.045 41.740 ;
        POLYGON 239.300 41.785 239.340 41.785 239.340 41.740 ;
        RECT 239.340 41.745 241.740 41.785 ;
        POLYGON 241.740 41.855 241.865 41.745 241.740 41.745 ;
        POLYGON 243.905 41.855 243.955 41.855 243.955 41.820 ;
        RECT 243.955 41.820 245.840 41.855 ;
        POLYGON 243.955 41.820 244.020 41.820 244.020 41.770 ;
        RECT 244.020 41.815 245.840 41.820 ;
        POLYGON 245.840 41.865 245.945 41.815 245.840 41.815 ;
        POLYGON 253.485 41.865 253.485 41.835 253.420 41.835 ;
        RECT 253.485 41.835 255.165 41.865 ;
        POLYGON 253.420 41.835 253.420 41.815 253.375 41.815 ;
        RECT 253.420 41.815 255.165 41.835 ;
        RECT 244.020 41.800 245.945 41.815 ;
        POLYGON 245.945 41.815 245.970 41.800 245.945 41.800 ;
        POLYGON 253.375 41.815 253.375 41.805 253.355 41.805 ;
        RECT 253.375 41.805 255.165 41.815 ;
        RECT 244.020 41.770 245.970 41.800 ;
        POLYGON 244.020 41.770 244.055 41.770 244.055 41.745 ;
        RECT 244.055 41.745 245.970 41.770 ;
        RECT 239.340 41.740 241.865 41.745 ;
        RECT 231.580 41.715 236.075 41.740 ;
        POLYGON 231.580 41.715 231.685 41.715 231.685 41.515 ;
        RECT 231.685 41.640 236.075 41.715 ;
        POLYGON 236.075 41.740 236.145 41.640 236.075 41.640 ;
        POLYGON 239.340 41.740 239.425 41.740 239.425 41.645 ;
        RECT 239.425 41.730 241.865 41.740 ;
        POLYGON 241.865 41.745 241.880 41.730 241.865 41.730 ;
        POLYGON 244.055 41.745 244.080 41.745 244.080 41.730 ;
        RECT 244.080 41.735 245.970 41.745 ;
        POLYGON 245.970 41.800 246.120 41.735 245.970 41.735 ;
        POLYGON 253.355 41.800 253.355 41.735 253.215 41.735 ;
        RECT 253.355 41.780 255.165 41.805 ;
        POLYGON 255.165 41.865 255.280 41.865 255.165 41.780 ;
        POLYGON 257.305 41.865 257.305 41.835 257.275 41.835 ;
        RECT 257.305 41.835 259.210 41.865 ;
        POLYGON 257.275 41.835 257.275 41.780 257.215 41.780 ;
        RECT 257.275 41.780 259.210 41.835 ;
        RECT 253.355 41.735 254.865 41.780 ;
        RECT 244.080 41.730 246.120 41.735 ;
        RECT 239.425 41.640 241.880 41.730 ;
        RECT 231.685 41.575 236.145 41.640 ;
        POLYGON 236.145 41.640 236.195 41.575 236.145 41.575 ;
        POLYGON 239.425 41.640 239.485 41.640 239.485 41.575 ;
        RECT 239.485 41.575 241.880 41.640 ;
        RECT 231.685 41.515 236.195 41.575 ;
        POLYGON 231.685 41.515 231.800 41.515 231.800 41.325 ;
        RECT 231.800 41.435 236.195 41.515 ;
        POLYGON 236.195 41.575 236.295 41.435 236.195 41.435 ;
        POLYGON 239.485 41.575 239.610 41.575 239.610 41.435 ;
        RECT 239.610 41.535 241.880 41.575 ;
        POLYGON 241.880 41.730 242.105 41.535 241.880 41.535 ;
        POLYGON 244.080 41.730 244.260 41.730 244.260 41.615 ;
        RECT 244.260 41.690 246.120 41.730 ;
        POLYGON 246.120 41.735 246.235 41.690 246.120 41.690 ;
        POLYGON 253.215 41.735 253.215 41.690 253.110 41.690 ;
        RECT 253.215 41.690 254.865 41.735 ;
        RECT 244.260 41.660 246.240 41.690 ;
        POLYGON 246.240 41.690 246.310 41.660 246.240 41.660 ;
        POLYGON 253.110 41.690 253.110 41.680 253.085 41.680 ;
        RECT 253.110 41.680 254.865 41.690 ;
        POLYGON 253.085 41.680 253.085 41.660 253.040 41.660 ;
        RECT 253.085 41.660 254.865 41.680 ;
        RECT 244.260 41.615 246.310 41.660 ;
        POLYGON 244.260 41.615 244.380 41.615 244.380 41.535 ;
        RECT 244.380 41.570 246.310 41.615 ;
        POLYGON 246.310 41.660 246.535 41.570 246.310 41.570 ;
        POLYGON 253.040 41.660 253.040 41.635 252.980 41.635 ;
        RECT 253.040 41.635 254.865 41.660 ;
        POLYGON 252.975 41.635 252.975 41.600 252.895 41.600 ;
        RECT 252.975 41.600 254.865 41.635 ;
        POLYGON 252.895 41.600 252.895 41.575 252.840 41.575 ;
        RECT 252.895 41.575 254.865 41.600 ;
        POLYGON 254.865 41.780 255.165 41.780 254.865 41.575 ;
        POLYGON 257.215 41.780 257.215 41.765 257.200 41.765 ;
        RECT 257.215 41.765 259.210 41.780 ;
        POLYGON 257.200 41.765 257.200 41.735 257.165 41.735 ;
        RECT 257.200 41.735 259.210 41.765 ;
        POLYGON 257.165 41.735 257.165 41.645 257.070 41.645 ;
        RECT 257.165 41.685 259.210 41.735 ;
        POLYGON 259.210 42.040 259.495 42.040 259.210 41.685 ;
        POLYGON 262.170 42.035 262.170 41.890 262.080 41.890 ;
        RECT 262.170 41.890 265.255 42.040 ;
        POLYGON 262.080 41.890 262.080 41.785 262.015 41.785 ;
        RECT 262.080 41.815 265.255 41.890 ;
        POLYGON 265.255 42.295 265.455 42.295 265.255 41.815 ;
        POLYGON 270.175 42.295 270.175 42.070 270.105 42.070 ;
        RECT 270.175 42.070 277.455 42.300 ;
        POLYGON 270.105 42.070 270.105 42.055 270.100 42.055 ;
        RECT 270.105 42.055 277.455 42.070 ;
        POLYGON 270.100 42.055 270.100 41.815 270.015 41.815 ;
        RECT 270.100 41.815 277.455 42.055 ;
        RECT 262.080 41.785 264.995 41.815 ;
        POLYGON 262.015 41.785 262.015 41.705 261.960 41.705 ;
        RECT 262.015 41.705 264.995 41.785 ;
        POLYGON 261.960 41.705 261.960 41.690 261.945 41.690 ;
        RECT 261.960 41.690 264.995 41.705 ;
        RECT 257.165 41.645 259.150 41.685 ;
        POLYGON 257.070 41.645 257.070 41.575 256.990 41.575 ;
        RECT 257.070 41.610 259.150 41.645 ;
        POLYGON 259.150 41.685 259.210 41.685 259.150 41.610 ;
        POLYGON 261.945 41.685 261.945 41.665 261.930 41.665 ;
        RECT 261.945 41.665 264.995 41.690 ;
        POLYGON 261.930 41.665 261.930 41.635 261.910 41.635 ;
        RECT 261.930 41.635 264.995 41.665 ;
        POLYGON 261.910 41.635 261.910 41.615 261.895 41.615 ;
        RECT 261.910 41.615 264.995 41.635 ;
        RECT 257.070 41.575 258.905 41.610 ;
        POLYGON 252.840 41.575 252.840 41.570 252.825 41.570 ;
        RECT 252.840 41.570 254.770 41.575 ;
        RECT 244.380 41.565 246.545 41.570 ;
        POLYGON 246.545 41.570 246.550 41.565 246.545 41.565 ;
        POLYGON 252.825 41.570 252.825 41.565 252.810 41.565 ;
        RECT 252.825 41.565 254.770 41.570 ;
        RECT 244.380 41.535 246.550 41.565 ;
        RECT 239.610 41.495 242.105 41.535 ;
        POLYGON 242.105 41.535 242.145 41.495 242.105 41.495 ;
        POLYGON 244.380 41.535 244.425 41.535 244.425 41.505 ;
        RECT 244.425 41.530 246.550 41.535 ;
        POLYGON 246.550 41.565 246.650 41.530 246.550 41.530 ;
        POLYGON 252.805 41.565 252.805 41.545 252.760 41.545 ;
        RECT 252.805 41.545 254.770 41.565 ;
        POLYGON 252.760 41.545 252.760 41.530 252.720 41.530 ;
        RECT 252.760 41.530 254.770 41.545 ;
        RECT 244.425 41.505 246.655 41.530 ;
        POLYGON 244.425 41.505 244.435 41.505 244.435 41.500 ;
        RECT 244.435 41.500 246.655 41.505 ;
        POLYGON 246.655 41.530 246.750 41.500 246.655 41.500 ;
        POLYGON 252.720 41.530 252.720 41.500 252.640 41.500 ;
        RECT 252.720 41.515 254.770 41.530 ;
        POLYGON 254.770 41.575 254.865 41.575 254.770 41.515 ;
        POLYGON 256.990 41.575 256.990 41.570 256.985 41.570 ;
        RECT 256.990 41.570 258.905 41.575 ;
        POLYGON 256.985 41.570 256.985 41.525 256.930 41.525 ;
        RECT 256.985 41.525 258.905 41.570 ;
        POLYGON 256.930 41.525 256.930 41.515 256.920 41.515 ;
        RECT 256.930 41.515 258.905 41.525 ;
        RECT 252.720 41.510 254.755 41.515 ;
        POLYGON 254.755 41.515 254.770 41.515 254.755 41.510 ;
        POLYGON 256.920 41.515 256.920 41.510 256.915 41.510 ;
        RECT 256.920 41.510 258.905 41.515 ;
        RECT 252.720 41.500 254.550 41.510 ;
        POLYGON 244.440 41.500 244.445 41.500 244.445 41.495 ;
        RECT 244.445 41.495 246.750 41.500 ;
        RECT 239.610 41.485 242.145 41.495 ;
        POLYGON 242.145 41.495 242.160 41.485 242.145 41.485 ;
        POLYGON 244.445 41.495 244.465 41.495 244.465 41.485 ;
        RECT 244.465 41.490 246.750 41.495 ;
        POLYGON 246.750 41.500 246.775 41.490 246.750 41.490 ;
        POLYGON 252.640 41.500 252.640 41.490 252.610 41.490 ;
        RECT 252.640 41.490 254.550 41.500 ;
        RECT 244.465 41.485 246.775 41.490 ;
        RECT 239.610 41.465 242.160 41.485 ;
        POLYGON 242.160 41.485 242.185 41.465 242.160 41.465 ;
        POLYGON 244.465 41.485 244.495 41.485 244.495 41.465 ;
        RECT 244.495 41.465 246.775 41.485 ;
        RECT 239.610 41.435 242.185 41.465 ;
        RECT 231.800 41.350 236.295 41.435 ;
        POLYGON 236.295 41.435 236.355 41.350 236.295 41.350 ;
        POLYGON 239.610 41.435 239.615 41.435 239.615 41.430 ;
        RECT 239.615 41.430 242.185 41.435 ;
        POLYGON 239.615 41.430 239.655 41.430 239.655 41.380 ;
        RECT 239.655 41.380 242.185 41.430 ;
        POLYGON 239.655 41.380 239.685 41.380 239.685 41.350 ;
        RECT 239.685 41.350 242.185 41.380 ;
        RECT 231.800 41.320 236.355 41.350 ;
        RECT 209.825 40.885 224.575 41.320 ;
        POLYGON 224.575 41.320 224.785 40.885 224.575 40.885 ;
        POLYGON 231.800 41.320 231.900 41.320 231.900 41.160 ;
        RECT 231.900 41.300 236.355 41.320 ;
        POLYGON 236.355 41.350 236.390 41.300 236.355 41.300 ;
        POLYGON 239.685 41.350 239.735 41.350 239.735 41.300 ;
        RECT 239.735 41.340 242.185 41.350 ;
        POLYGON 242.185 41.465 242.340 41.340 242.185 41.340 ;
        POLYGON 244.495 41.465 244.705 41.465 244.705 41.340 ;
        RECT 244.705 41.425 246.775 41.465 ;
        POLYGON 246.775 41.490 246.970 41.425 246.775 41.425 ;
        POLYGON 252.610 41.490 252.610 41.465 252.545 41.465 ;
        RECT 252.610 41.465 254.550 41.490 ;
        POLYGON 252.545 41.465 252.545 41.460 252.525 41.460 ;
        RECT 252.545 41.460 254.550 41.465 ;
        POLYGON 252.525 41.460 252.525 41.445 252.490 41.445 ;
        RECT 252.525 41.445 254.550 41.460 ;
        POLYGON 252.490 41.445 252.490 41.425 252.430 41.425 ;
        RECT 252.490 41.425 254.550 41.445 ;
        RECT 244.705 41.420 246.970 41.425 ;
        POLYGON 246.970 41.425 246.975 41.420 246.970 41.420 ;
        POLYGON 252.430 41.425 252.430 41.420 252.415 41.420 ;
        RECT 252.430 41.420 254.550 41.425 ;
        RECT 244.705 41.410 246.975 41.420 ;
        POLYGON 246.975 41.420 247.010 41.410 246.975 41.410 ;
        POLYGON 252.415 41.420 252.415 41.410 252.385 41.410 ;
        RECT 252.415 41.410 254.550 41.420 ;
        RECT 244.705 41.390 247.010 41.410 ;
        POLYGON 247.010 41.410 247.075 41.390 247.010 41.390 ;
        POLYGON 252.385 41.410 252.385 41.390 252.325 41.390 ;
        RECT 252.385 41.390 254.550 41.410 ;
        RECT 244.705 41.355 247.075 41.390 ;
        POLYGON 247.075 41.390 247.195 41.355 247.075 41.355 ;
        POLYGON 252.325 41.390 252.325 41.355 252.210 41.355 ;
        RECT 252.325 41.380 254.550 41.390 ;
        POLYGON 254.550 41.510 254.755 41.510 254.550 41.380 ;
        POLYGON 256.915 41.510 256.915 41.380 256.760 41.380 ;
        RECT 256.915 41.380 258.905 41.510 ;
        RECT 252.325 41.355 254.230 41.380 ;
        RECT 244.705 41.345 247.195 41.355 ;
        POLYGON 247.195 41.355 247.240 41.345 247.195 41.345 ;
        POLYGON 252.210 41.355 252.210 41.345 252.180 41.345 ;
        RECT 252.210 41.345 254.230 41.355 ;
        RECT 244.705 41.340 247.245 41.345 ;
        RECT 239.735 41.300 242.340 41.340 ;
        RECT 231.900 41.165 236.390 41.300 ;
        POLYGON 236.390 41.300 236.485 41.165 236.390 41.165 ;
        POLYGON 239.735 41.300 239.870 41.300 239.870 41.165 ;
        RECT 239.870 41.185 242.340 41.300 ;
        POLYGON 242.340 41.340 242.525 41.185 242.340 41.185 ;
        POLYGON 244.705 41.340 244.840 41.340 244.840 41.260 ;
        RECT 244.840 41.295 247.245 41.340 ;
        POLYGON 247.245 41.345 247.395 41.295 247.245 41.295 ;
        POLYGON 252.180 41.345 252.180 41.330 252.130 41.330 ;
        RECT 252.180 41.330 254.230 41.345 ;
        POLYGON 252.130 41.330 252.130 41.320 252.100 41.320 ;
        RECT 252.130 41.320 254.230 41.330 ;
        POLYGON 252.095 41.320 252.095 41.310 252.065 41.310 ;
        RECT 252.095 41.310 254.230 41.320 ;
        POLYGON 252.065 41.310 252.065 41.295 252.005 41.295 ;
        RECT 252.065 41.295 254.230 41.310 ;
        RECT 244.840 41.290 247.395 41.295 ;
        POLYGON 247.395 41.295 247.425 41.290 247.395 41.290 ;
        POLYGON 252.005 41.295 252.005 41.290 251.985 41.290 ;
        RECT 252.005 41.290 254.230 41.295 ;
        RECT 244.840 41.270 247.425 41.290 ;
        POLYGON 247.425 41.290 247.505 41.270 247.425 41.270 ;
        POLYGON 251.985 41.290 251.985 41.275 251.925 41.275 ;
        RECT 251.985 41.275 254.230 41.290 ;
        POLYGON 251.920 41.275 251.920 41.270 251.905 41.270 ;
        RECT 251.920 41.270 254.230 41.275 ;
        RECT 244.840 41.260 247.510 41.270 ;
        POLYGON 244.840 41.260 244.900 41.260 244.900 41.230 ;
        RECT 244.900 41.230 247.510 41.260 ;
        POLYGON 244.900 41.230 244.985 41.230 244.985 41.185 ;
        RECT 244.985 41.215 247.510 41.230 ;
        POLYGON 247.510 41.270 247.735 41.215 247.510 41.215 ;
        POLYGON 251.905 41.270 251.905 41.255 251.860 41.255 ;
        RECT 251.905 41.255 254.230 41.270 ;
        POLYGON 251.860 41.255 251.860 41.230 251.765 41.230 ;
        RECT 251.860 41.230 254.230 41.255 ;
        POLYGON 251.765 41.230 251.765 41.215 251.700 41.215 ;
        RECT 251.765 41.215 254.230 41.230 ;
        RECT 244.985 41.195 247.740 41.215 ;
        POLYGON 247.740 41.215 247.815 41.195 247.740 41.195 ;
        POLYGON 251.700 41.215 251.700 41.195 251.615 41.195 ;
        RECT 251.700 41.195 254.230 41.215 ;
        RECT 244.985 41.185 247.815 41.195 ;
        RECT 239.870 41.165 242.525 41.185 ;
        RECT 231.900 41.160 236.485 41.165 ;
        POLYGON 231.900 41.160 232.065 41.160 232.065 40.885 ;
        RECT 232.065 41.125 236.485 41.160 ;
        POLYGON 236.485 41.165 236.510 41.125 236.485 41.125 ;
        POLYGON 239.870 41.165 239.910 41.165 239.910 41.125 ;
        RECT 239.910 41.150 242.525 41.165 ;
        POLYGON 242.525 41.185 242.570 41.150 242.525 41.150 ;
        POLYGON 244.985 41.185 245.050 41.185 245.050 41.150 ;
        RECT 245.050 41.180 247.815 41.185 ;
        POLYGON 247.815 41.195 247.895 41.180 247.815 41.180 ;
        POLYGON 251.605 41.195 251.605 41.180 251.545 41.180 ;
        RECT 251.605 41.190 254.230 41.195 ;
        POLYGON 254.230 41.380 254.550 41.380 254.230 41.190 ;
        POLYGON 256.760 41.380 256.760 41.375 256.755 41.375 ;
        RECT 256.760 41.375 258.905 41.380 ;
        POLYGON 256.755 41.375 256.755 41.345 256.720 41.345 ;
        RECT 256.755 41.345 258.905 41.375 ;
        POLYGON 256.720 41.345 256.720 41.315 256.680 41.315 ;
        RECT 256.720 41.330 258.905 41.345 ;
        POLYGON 258.905 41.610 259.150 41.610 258.905 41.330 ;
        POLYGON 261.895 41.610 261.895 41.590 261.880 41.590 ;
        RECT 261.895 41.590 264.995 41.615 ;
        POLYGON 261.880 41.590 261.880 41.535 261.840 41.535 ;
        RECT 261.880 41.535 264.995 41.590 ;
        POLYGON 261.840 41.535 261.840 41.465 261.790 41.465 ;
        RECT 261.840 41.465 264.995 41.535 ;
        POLYGON 261.790 41.465 261.790 41.405 261.750 41.405 ;
        RECT 261.790 41.405 264.995 41.465 ;
        POLYGON 261.750 41.405 261.750 41.380 261.735 41.380 ;
        RECT 261.750 41.380 264.995 41.405 ;
        POLYGON 261.735 41.380 261.735 41.335 261.700 41.335 ;
        RECT 261.735 41.335 264.995 41.380 ;
        RECT 256.720 41.315 258.790 41.330 ;
        POLYGON 256.680 41.315 256.680 41.230 256.570 41.230 ;
        RECT 256.680 41.230 258.790 41.315 ;
        POLYGON 256.570 41.230 256.570 41.190 256.520 41.190 ;
        RECT 256.570 41.195 258.790 41.230 ;
        POLYGON 258.790 41.330 258.905 41.330 258.790 41.195 ;
        POLYGON 261.700 41.330 261.700 41.195 261.595 41.195 ;
        RECT 261.700 41.270 264.995 41.335 ;
        POLYGON 264.995 41.815 265.255 41.815 264.995 41.270 ;
        POLYGON 270.015 41.815 270.015 41.445 269.885 41.445 ;
        RECT 270.015 41.495 277.455 41.815 ;
        POLYGON 277.455 42.840 277.650 42.840 277.455 41.495 ;
        POLYGON 287.715 42.835 287.715 41.495 287.645 41.495 ;
        RECT 287.715 41.495 303.120 42.840 ;
        RECT 270.015 41.445 277.205 41.495 ;
        POLYGON 269.885 41.445 269.885 41.335 269.845 41.335 ;
        RECT 269.885 41.335 277.205 41.445 ;
        POLYGON 269.845 41.335 269.845 41.315 269.840 41.315 ;
        RECT 269.845 41.315 277.205 41.335 ;
        POLYGON 269.840 41.315 269.840 41.270 269.820 41.270 ;
        RECT 269.840 41.270 277.205 41.315 ;
        RECT 261.700 41.195 264.850 41.270 ;
        RECT 256.570 41.190 258.750 41.195 ;
        RECT 251.605 41.180 254.185 41.190 ;
        RECT 245.050 41.170 247.895 41.180 ;
        POLYGON 247.895 41.180 247.945 41.170 247.895 41.170 ;
        POLYGON 251.545 41.180 251.545 41.170 251.505 41.170 ;
        RECT 251.545 41.170 254.185 41.180 ;
        RECT 245.050 41.155 247.945 41.170 ;
        POLYGON 247.945 41.170 248.005 41.155 247.945 41.155 ;
        POLYGON 251.505 41.170 251.505 41.155 251.445 41.155 ;
        RECT 251.505 41.165 254.185 41.170 ;
        POLYGON 254.185 41.190 254.230 41.190 254.185 41.165 ;
        POLYGON 256.520 41.190 256.520 41.185 256.515 41.185 ;
        RECT 256.520 41.185 258.750 41.190 ;
        POLYGON 256.515 41.185 256.515 41.165 256.490 41.165 ;
        RECT 256.515 41.165 258.750 41.185 ;
        RECT 251.505 41.155 254.090 41.165 ;
        RECT 245.050 41.150 248.010 41.155 ;
        RECT 239.910 41.140 242.570 41.150 ;
        POLYGON 242.570 41.150 242.585 41.140 242.570 41.140 ;
        POLYGON 245.050 41.150 245.070 41.150 245.070 41.140 ;
        RECT 245.070 41.140 248.010 41.150 ;
        RECT 239.910 41.125 242.585 41.140 ;
        RECT 232.065 41.070 236.510 41.125 ;
        POLYGON 236.510 41.125 236.555 41.070 236.510 41.070 ;
        POLYGON 239.910 41.125 239.965 41.125 239.965 41.070 ;
        RECT 239.965 41.070 242.585 41.125 ;
        RECT 232.065 40.885 236.555 41.070 ;
        RECT 209.825 40.540 224.785 40.885 ;
        POLYGON 209.825 40.540 210.035 40.540 210.035 40.075 ;
        RECT 210.035 40.510 224.785 40.540 ;
        POLYGON 224.785 40.885 224.970 40.510 224.785 40.510 ;
        POLYGON 232.065 40.885 232.075 40.885 232.075 40.870 ;
        RECT 232.075 40.870 236.555 40.885 ;
        POLYGON 232.075 40.870 232.240 40.870 232.240 40.625 ;
        RECT 232.240 40.855 236.555 40.870 ;
        POLYGON 236.555 41.070 236.725 40.855 236.555 40.855 ;
        POLYGON 239.965 41.070 240.180 41.070 240.180 40.855 ;
        RECT 240.180 40.955 242.585 41.070 ;
        POLYGON 242.585 41.140 242.840 40.955 242.585 40.955 ;
        POLYGON 245.070 41.140 245.090 41.140 245.090 41.130 ;
        RECT 245.090 41.130 248.010 41.140 ;
        POLYGON 245.095 41.130 245.265 41.130 245.265 41.040 ;
        RECT 245.265 41.110 248.010 41.130 ;
        POLYGON 248.010 41.155 248.230 41.110 248.010 41.110 ;
        POLYGON 251.445 41.155 251.445 41.150 251.425 41.150 ;
        RECT 251.445 41.150 254.090 41.155 ;
        POLYGON 251.420 41.150 251.420 41.145 251.395 41.145 ;
        RECT 251.420 41.145 254.090 41.150 ;
        POLYGON 251.395 41.145 251.395 41.140 251.350 41.140 ;
        RECT 251.395 41.140 254.090 41.145 ;
        POLYGON 251.350 41.140 251.350 41.135 251.345 41.135 ;
        RECT 251.350 41.135 254.090 41.140 ;
        POLYGON 251.345 41.135 251.345 41.110 251.200 41.110 ;
        RECT 251.345 41.115 254.090 41.135 ;
        POLYGON 254.090 41.165 254.185 41.165 254.090 41.115 ;
        POLYGON 256.490 41.165 256.490 41.115 256.420 41.115 ;
        RECT 256.490 41.155 258.750 41.165 ;
        POLYGON 258.750 41.195 258.790 41.195 258.750 41.155 ;
        POLYGON 261.595 41.195 261.595 41.155 261.565 41.155 ;
        RECT 261.595 41.155 264.850 41.195 ;
        RECT 256.490 41.115 258.410 41.155 ;
        RECT 251.345 41.110 253.925 41.115 ;
        RECT 245.265 41.105 248.230 41.110 ;
        POLYGON 248.230 41.110 248.290 41.105 248.230 41.105 ;
        POLYGON 251.200 41.110 251.200 41.105 251.175 41.105 ;
        RECT 251.200 41.105 253.925 41.110 ;
        RECT 245.265 41.100 248.295 41.105 ;
        POLYGON 248.295 41.105 248.315 41.100 248.295 41.100 ;
        POLYGON 251.175 41.105 251.175 41.100 251.145 41.100 ;
        RECT 251.175 41.100 253.925 41.105 ;
        RECT 245.265 41.090 248.315 41.100 ;
        POLYGON 248.315 41.100 248.380 41.090 248.315 41.090 ;
        POLYGON 251.140 41.100 251.140 41.090 251.070 41.090 ;
        RECT 251.140 41.090 253.925 41.100 ;
        RECT 245.265 41.050 248.390 41.090 ;
        POLYGON 248.390 41.090 248.645 41.050 248.390 41.050 ;
        POLYGON 251.065 41.090 251.065 41.080 251.020 41.080 ;
        RECT 251.065 41.080 253.925 41.090 ;
        POLYGON 251.020 41.080 251.020 41.065 250.910 41.065 ;
        RECT 251.020 41.065 253.925 41.080 ;
        POLYGON 250.910 41.065 250.910 41.050 250.795 41.050 ;
        RECT 250.910 41.050 253.925 41.065 ;
        RECT 245.265 41.040 248.645 41.050 ;
        POLYGON 245.265 41.040 245.435 41.040 245.435 40.955 ;
        RECT 245.435 41.030 248.645 41.040 ;
        POLYGON 248.645 41.050 248.840 41.030 248.645 41.030 ;
        POLYGON 250.795 41.050 250.795 41.035 250.680 41.035 ;
        RECT 250.795 41.035 253.925 41.050 ;
        POLYGON 250.680 41.035 250.680 41.030 250.635 41.030 ;
        RECT 250.680 41.030 253.925 41.035 ;
        RECT 245.435 41.025 248.845 41.030 ;
        POLYGON 248.845 41.030 248.875 41.025 248.845 41.025 ;
        POLYGON 250.635 41.030 250.635 41.025 250.570 41.025 ;
        RECT 250.635 41.025 253.925 41.030 ;
        POLYGON 253.925 41.115 254.090 41.115 253.925 41.025 ;
        POLYGON 256.420 41.115 256.420 41.025 256.305 41.025 ;
        RECT 256.420 41.025 258.410 41.115 ;
        RECT 245.435 41.020 248.875 41.025 ;
        POLYGON 248.875 41.025 248.935 41.020 248.875 41.020 ;
        POLYGON 250.570 41.025 250.570 41.020 250.505 41.020 ;
        RECT 250.570 41.020 253.900 41.025 ;
        RECT 245.435 41.010 248.965 41.020 ;
        POLYGON 248.965 41.020 249.050 41.010 248.965 41.010 ;
        POLYGON 250.505 41.020 250.505 41.015 250.440 41.015 ;
        RECT 250.505 41.015 253.900 41.020 ;
        POLYGON 250.435 41.015 250.435 41.010 250.430 41.010 ;
        RECT 250.435 41.010 253.900 41.015 ;
        POLYGON 253.900 41.025 253.925 41.025 253.900 41.010 ;
        POLYGON 256.305 41.025 256.305 41.010 256.285 41.010 ;
        RECT 256.305 41.010 258.410 41.025 ;
        RECT 245.435 40.995 249.050 41.010 ;
        POLYGON 249.050 41.010 249.295 40.995 249.050 40.995 ;
        POLYGON 250.400 41.010 250.400 40.995 250.245 40.995 ;
        RECT 250.400 40.995 253.670 41.010 ;
        RECT 245.435 40.990 249.300 40.995 ;
        POLYGON 249.300 40.995 249.365 40.990 249.300 40.990 ;
        POLYGON 250.220 40.995 250.220 40.990 250.100 40.990 ;
        RECT 250.220 40.990 253.670 40.995 ;
        RECT 245.435 40.985 249.380 40.990 ;
        POLYGON 249.380 40.990 249.455 40.985 249.380 40.985 ;
        POLYGON 250.100 40.990 250.100 40.985 249.975 40.985 ;
        RECT 250.100 40.985 253.670 40.990 ;
        RECT 245.435 40.980 249.850 40.985 ;
        POLYGON 249.850 40.985 249.855 40.980 249.850 40.980 ;
        POLYGON 249.975 40.985 249.975 40.980 249.855 40.980 ;
        RECT 249.975 40.980 253.670 40.985 ;
        RECT 245.435 40.955 253.670 40.980 ;
        RECT 240.180 40.925 242.840 40.955 ;
        POLYGON 242.840 40.955 242.880 40.925 242.840 40.925 ;
        POLYGON 245.435 40.955 245.500 40.955 245.500 40.925 ;
        RECT 245.500 40.925 253.670 40.955 ;
        RECT 240.180 40.920 242.880 40.925 ;
        POLYGON 242.880 40.925 242.885 40.920 242.880 40.920 ;
        POLYGON 245.500 40.925 245.515 40.925 245.515 40.920 ;
        RECT 245.515 40.920 253.670 40.925 ;
        RECT 240.180 40.855 242.885 40.920 ;
        RECT 232.240 40.760 236.725 40.855 ;
        POLYGON 236.725 40.855 236.800 40.760 236.725 40.760 ;
        POLYGON 240.180 40.855 240.225 40.855 240.225 40.810 ;
        RECT 240.225 40.825 242.885 40.855 ;
        POLYGON 242.885 40.920 243.010 40.825 242.885 40.825 ;
        POLYGON 245.515 40.920 245.580 40.920 245.580 40.890 ;
        RECT 245.580 40.895 253.670 40.920 ;
        POLYGON 253.670 41.010 253.900 41.010 253.670 40.895 ;
        POLYGON 256.285 41.010 256.285 41.000 256.270 41.000 ;
        RECT 256.285 41.000 258.410 41.010 ;
        POLYGON 256.270 41.000 256.270 40.995 256.265 40.995 ;
        RECT 256.270 40.995 258.410 41.000 ;
        POLYGON 256.265 40.995 256.265 40.990 256.255 40.990 ;
        RECT 256.265 40.990 258.410 40.995 ;
        POLYGON 256.255 40.990 256.255 40.950 256.200 40.950 ;
        RECT 256.255 40.950 258.410 40.990 ;
        POLYGON 256.200 40.950 256.200 40.895 256.120 40.895 ;
        RECT 256.200 40.895 258.410 40.950 ;
        RECT 245.580 40.890 253.505 40.895 ;
        POLYGON 245.580 40.890 245.665 40.890 245.665 40.850 ;
        RECT 245.665 40.850 253.505 40.890 ;
        POLYGON 245.665 40.850 245.715 40.850 245.715 40.825 ;
        RECT 245.715 40.825 253.505 40.850 ;
        RECT 240.225 40.810 243.010 40.825 ;
        POLYGON 240.225 40.810 240.255 40.810 240.255 40.785 ;
        RECT 240.255 40.785 243.010 40.810 ;
        POLYGON 240.255 40.785 240.280 40.785 240.280 40.760 ;
        RECT 240.280 40.765 243.010 40.785 ;
        POLYGON 243.010 40.825 243.100 40.765 243.010 40.765 ;
        POLYGON 245.715 40.825 245.815 40.825 245.815 40.780 ;
        RECT 245.815 40.815 253.505 40.825 ;
        POLYGON 253.505 40.895 253.670 40.895 253.505 40.815 ;
        POLYGON 256.120 40.895 256.120 40.815 256.005 40.815 ;
        RECT 256.120 40.815 258.410 40.895 ;
        RECT 245.815 40.780 253.420 40.815 ;
        POLYGON 245.815 40.780 245.845 40.780 245.845 40.765 ;
        RECT 245.845 40.775 253.420 40.780 ;
        POLYGON 253.420 40.815 253.505 40.815 253.420 40.775 ;
        POLYGON 256.005 40.815 256.005 40.775 255.950 40.775 ;
        RECT 256.005 40.795 258.410 40.815 ;
        POLYGON 258.410 41.155 258.750 41.155 258.410 40.795 ;
        POLYGON 261.565 41.155 261.565 41.050 261.485 41.050 ;
        RECT 261.565 41.050 264.850 41.155 ;
        POLYGON 261.485 41.050 261.485 41.010 261.455 41.010 ;
        RECT 261.485 41.010 264.850 41.050 ;
        POLYGON 261.455 41.010 261.455 40.795 261.280 40.795 ;
        RECT 261.455 40.980 264.850 41.010 ;
        POLYGON 264.850 41.270 264.995 41.270 264.850 40.980 ;
        POLYGON 269.820 41.265 269.820 40.985 269.710 40.985 ;
        RECT 269.820 40.985 277.205 41.270 ;
        RECT 261.455 40.795 264.720 40.980 ;
        RECT 256.005 40.775 258.295 40.795 ;
        RECT 245.845 40.770 253.415 40.775 ;
        POLYGON 253.415 40.775 253.420 40.775 253.415 40.770 ;
        POLYGON 255.950 40.775 255.950 40.770 255.940 40.770 ;
        RECT 255.950 40.770 258.295 40.775 ;
        RECT 245.845 40.765 253.235 40.770 ;
        RECT 240.280 40.760 243.100 40.765 ;
        RECT 232.240 40.625 236.800 40.760 ;
        POLYGON 232.240 40.625 232.310 40.625 232.310 40.515 ;
        RECT 232.310 40.510 236.800 40.625 ;
        RECT 210.035 40.075 224.970 40.510 ;
        POLYGON 210.035 40.075 210.290 40.075 210.290 39.500 ;
        RECT 210.290 40.020 224.970 40.075 ;
        POLYGON 224.970 40.510 225.225 40.020 224.970 40.020 ;
        POLYGON 232.310 40.510 232.500 40.510 232.500 40.225 ;
        RECT 232.500 40.495 236.800 40.510 ;
        POLYGON 236.800 40.760 237.005 40.495 236.800 40.495 ;
        POLYGON 240.280 40.760 240.335 40.760 240.335 40.710 ;
        RECT 240.335 40.710 243.100 40.760 ;
        POLYGON 240.335 40.710 240.575 40.710 240.575 40.495 ;
        RECT 240.575 40.665 243.100 40.710 ;
        POLYGON 243.100 40.765 243.245 40.665 243.100 40.665 ;
        POLYGON 245.845 40.765 245.940 40.765 245.940 40.725 ;
        RECT 245.940 40.725 253.235 40.765 ;
        POLYGON 245.940 40.725 246.080 40.725 246.080 40.665 ;
        RECT 246.080 40.695 253.235 40.725 ;
        POLYGON 253.235 40.770 253.415 40.770 253.235 40.695 ;
        POLYGON 255.940 40.770 255.940 40.700 255.840 40.700 ;
        RECT 255.940 40.700 258.295 40.770 ;
        POLYGON 255.840 40.700 255.840 40.695 255.835 40.695 ;
        RECT 255.840 40.695 258.295 40.700 ;
        RECT 246.080 40.665 253.165 40.695 ;
        POLYGON 253.165 40.695 253.235 40.695 253.165 40.665 ;
        POLYGON 255.835 40.695 255.835 40.680 255.815 40.680 ;
        RECT 255.835 40.685 258.295 40.695 ;
        POLYGON 258.295 40.795 258.410 40.795 258.295 40.685 ;
        POLYGON 261.280 40.790 261.280 40.685 261.190 40.685 ;
        RECT 261.280 40.730 264.720 40.795 ;
        POLYGON 264.720 40.980 264.850 40.980 264.720 40.730 ;
        POLYGON 269.710 40.980 269.710 40.730 269.610 40.730 ;
        RECT 269.710 40.730 277.205 40.985 ;
        RECT 261.280 40.685 264.420 40.730 ;
        RECT 255.835 40.680 258.135 40.685 ;
        POLYGON 255.815 40.680 255.815 40.665 255.790 40.665 ;
        RECT 255.815 40.665 258.135 40.680 ;
        RECT 240.575 40.580 243.245 40.665 ;
        POLYGON 243.245 40.665 243.375 40.580 243.245 40.580 ;
        POLYGON 246.080 40.665 246.215 40.665 246.215 40.610 ;
        RECT 246.215 40.610 252.980 40.665 ;
        POLYGON 246.220 40.610 246.245 40.610 246.245 40.600 ;
        RECT 246.245 40.600 252.980 40.610 ;
        POLYGON 246.245 40.600 246.285 40.600 246.285 40.580 ;
        RECT 246.285 40.585 252.980 40.600 ;
        POLYGON 252.980 40.665 253.165 40.665 252.980 40.585 ;
        POLYGON 255.790 40.665 255.790 40.655 255.775 40.655 ;
        RECT 255.790 40.655 258.135 40.665 ;
        POLYGON 255.775 40.655 255.775 40.630 255.735 40.630 ;
        RECT 255.775 40.630 258.135 40.655 ;
        POLYGON 255.735 40.630 255.735 40.585 255.665 40.585 ;
        RECT 255.735 40.585 258.135 40.630 ;
        RECT 246.285 40.580 252.970 40.585 ;
        POLYGON 252.970 40.585 252.980 40.585 252.970 40.580 ;
        POLYGON 255.665 40.585 255.665 40.580 255.655 40.580 ;
        RECT 255.665 40.580 258.135 40.585 ;
        RECT 240.575 40.515 243.375 40.580 ;
        POLYGON 243.375 40.580 243.470 40.515 243.375 40.515 ;
        POLYGON 246.285 40.580 246.310 40.580 246.310 40.570 ;
        RECT 246.310 40.570 252.905 40.580 ;
        POLYGON 246.310 40.570 246.460 40.570 246.460 40.515 ;
        RECT 246.460 40.555 252.905 40.570 ;
        POLYGON 252.905 40.580 252.970 40.580 252.905 40.555 ;
        POLYGON 255.655 40.580 255.655 40.555 255.615 40.555 ;
        RECT 255.655 40.555 258.135 40.580 ;
        RECT 246.460 40.515 252.760 40.555 ;
        RECT 240.575 40.495 243.470 40.515 ;
        RECT 232.500 40.475 237.005 40.495 ;
        POLYGON 237.005 40.495 237.025 40.475 237.005 40.475 ;
        POLYGON 240.575 40.495 240.595 40.495 240.595 40.475 ;
        RECT 240.595 40.475 243.470 40.495 ;
        RECT 232.500 40.405 237.025 40.475 ;
        POLYGON 237.025 40.475 237.085 40.405 237.025 40.405 ;
        POLYGON 240.595 40.475 240.675 40.475 240.675 40.405 ;
        RECT 240.675 40.420 243.470 40.475 ;
        POLYGON 243.470 40.515 243.625 40.420 243.470 40.420 ;
        POLYGON 246.460 40.515 246.505 40.515 246.505 40.500 ;
        RECT 246.505 40.505 252.760 40.515 ;
        POLYGON 252.760 40.555 252.905 40.555 252.760 40.505 ;
        POLYGON 255.615 40.555 255.615 40.505 255.535 40.505 ;
        RECT 255.615 40.535 258.135 40.555 ;
        POLYGON 258.135 40.685 258.295 40.685 258.135 40.535 ;
        POLYGON 261.190 40.680 261.190 40.555 261.085 40.555 ;
        RECT 261.190 40.555 264.420 40.685 ;
        POLYGON 261.085 40.555 261.085 40.535 261.070 40.535 ;
        RECT 261.085 40.535 264.420 40.555 ;
        RECT 255.615 40.505 258.010 40.535 ;
        RECT 246.505 40.500 252.705 40.505 ;
        POLYGON 246.505 40.500 246.545 40.500 246.545 40.485 ;
        RECT 246.545 40.485 252.705 40.500 ;
        POLYGON 252.705 40.505 252.760 40.505 252.705 40.485 ;
        POLYGON 255.535 40.505 255.535 40.485 255.505 40.485 ;
        RECT 255.535 40.485 258.010 40.505 ;
        POLYGON 246.545 40.485 246.755 40.485 246.755 40.420 ;
        RECT 246.755 40.465 252.635 40.485 ;
        POLYGON 252.635 40.485 252.705 40.485 252.635 40.465 ;
        POLYGON 255.505 40.485 255.505 40.465 255.470 40.465 ;
        RECT 255.505 40.465 258.010 40.485 ;
        RECT 246.755 40.435 252.545 40.465 ;
        POLYGON 252.545 40.465 252.635 40.465 252.545 40.435 ;
        POLYGON 255.470 40.465 255.470 40.435 255.425 40.435 ;
        RECT 255.470 40.435 258.010 40.465 ;
        RECT 246.755 40.420 252.435 40.435 ;
        RECT 240.675 40.405 243.630 40.420 ;
        RECT 232.500 40.225 237.085 40.405 ;
        POLYGON 232.500 40.225 232.650 40.225 232.650 40.020 ;
        RECT 232.650 40.115 237.085 40.225 ;
        POLYGON 237.085 40.405 237.335 40.115 237.085 40.115 ;
        POLYGON 240.675 40.405 240.830 40.405 240.830 40.270 ;
        RECT 240.830 40.400 243.630 40.405 ;
        POLYGON 243.630 40.420 243.660 40.400 243.630 40.400 ;
        POLYGON 246.755 40.420 246.775 40.420 246.775 40.415 ;
        RECT 246.775 40.415 252.435 40.420 ;
        POLYGON 246.775 40.415 246.820 40.415 246.820 40.400 ;
        RECT 246.820 40.405 252.435 40.415 ;
        POLYGON 252.435 40.435 252.545 40.435 252.435 40.405 ;
        POLYGON 255.425 40.435 255.425 40.430 255.420 40.430 ;
        RECT 255.425 40.430 258.010 40.435 ;
        POLYGON 255.420 40.430 255.420 40.415 255.395 40.415 ;
        RECT 255.420 40.415 258.010 40.430 ;
        POLYGON 258.010 40.535 258.135 40.535 258.010 40.415 ;
        POLYGON 261.070 40.535 261.070 40.415 260.970 40.415 ;
        RECT 261.070 40.415 264.420 40.535 ;
        POLYGON 255.395 40.415 255.395 40.405 255.375 40.405 ;
        RECT 255.395 40.405 257.850 40.415 ;
        RECT 246.820 40.400 252.350 40.405 ;
        RECT 240.830 40.270 243.660 40.400 ;
        POLYGON 240.830 40.270 241.010 40.270 241.010 40.130 ;
        RECT 241.010 40.225 243.660 40.270 ;
        POLYGON 243.660 40.400 243.950 40.225 243.660 40.225 ;
        POLYGON 246.820 40.400 247.010 40.400 247.010 40.350 ;
        RECT 247.010 40.380 252.350 40.400 ;
        POLYGON 252.350 40.405 252.435 40.405 252.350 40.380 ;
        POLYGON 255.375 40.405 255.375 40.380 255.335 40.380 ;
        RECT 255.375 40.380 257.850 40.405 ;
        RECT 247.010 40.375 252.325 40.380 ;
        POLYGON 252.325 40.380 252.350 40.380 252.325 40.375 ;
        POLYGON 255.335 40.380 255.335 40.375 255.325 40.375 ;
        RECT 255.335 40.375 257.850 40.380 ;
        RECT 247.010 40.350 252.155 40.375 ;
        POLYGON 247.010 40.350 247.080 40.350 247.080 40.335 ;
        RECT 247.080 40.335 252.155 40.350 ;
        POLYGON 252.155 40.375 252.325 40.375 252.155 40.335 ;
        POLYGON 255.325 40.375 255.325 40.350 255.280 40.350 ;
        RECT 255.325 40.350 257.850 40.375 ;
        POLYGON 255.280 40.350 255.280 40.335 255.255 40.335 ;
        RECT 255.280 40.335 257.850 40.350 ;
        POLYGON 247.085 40.335 247.130 40.335 247.130 40.325 ;
        RECT 247.130 40.325 252.045 40.335 ;
        POLYGON 247.130 40.325 247.245 40.325 247.245 40.300 ;
        RECT 247.245 40.315 252.045 40.325 ;
        POLYGON 252.045 40.335 252.155 40.335 252.045 40.315 ;
        POLYGON 255.255 40.335 255.255 40.315 255.225 40.315 ;
        RECT 255.255 40.315 257.850 40.335 ;
        RECT 247.245 40.300 251.860 40.315 ;
        POLYGON 247.245 40.300 247.340 40.300 247.340 40.280 ;
        RECT 247.340 40.280 251.860 40.300 ;
        POLYGON 251.860 40.315 252.040 40.315 251.860 40.280 ;
        POLYGON 255.225 40.315 255.225 40.280 255.165 40.280 ;
        RECT 255.225 40.280 257.850 40.315 ;
        POLYGON 247.340 40.280 247.480 40.280 247.480 40.255 ;
        RECT 247.480 40.255 251.615 40.280 ;
        POLYGON 247.485 40.255 247.585 40.255 247.585 40.240 ;
        RECT 247.585 40.245 251.615 40.255 ;
        POLYGON 251.615 40.280 251.855 40.280 251.615 40.245 ;
        POLYGON 255.165 40.280 255.165 40.245 255.105 40.245 ;
        RECT 255.165 40.275 257.850 40.280 ;
        POLYGON 257.850 40.415 258.010 40.415 257.850 40.275 ;
        POLYGON 260.970 40.415 260.970 40.385 260.945 40.385 ;
        RECT 260.970 40.385 264.420 40.415 ;
        POLYGON 260.945 40.385 260.945 40.275 260.855 40.275 ;
        RECT 260.945 40.275 264.420 40.385 ;
        RECT 255.165 40.245 257.595 40.275 ;
        RECT 247.585 40.240 251.530 40.245 ;
        POLYGON 247.590 40.240 247.700 40.240 247.700 40.225 ;
        RECT 247.700 40.235 251.530 40.240 ;
        POLYGON 251.530 40.245 251.615 40.245 251.530 40.235 ;
        POLYGON 255.105 40.245 255.105 40.235 255.085 40.235 ;
        RECT 255.105 40.235 257.595 40.245 ;
        RECT 247.700 40.225 251.350 40.235 ;
        RECT 241.010 40.220 243.950 40.225 ;
        POLYGON 243.950 40.225 243.955 40.220 243.950 40.220 ;
        POLYGON 247.700 40.225 247.740 40.225 247.740 40.220 ;
        RECT 247.740 40.220 251.350 40.225 ;
        RECT 241.010 40.185 243.955 40.220 ;
        POLYGON 243.955 40.220 244.020 40.185 243.955 40.185 ;
        POLYGON 247.740 40.220 247.835 40.220 247.835 40.210 ;
        RECT 247.835 40.215 251.350 40.220 ;
        POLYGON 251.350 40.235 251.530 40.235 251.350 40.215 ;
        POLYGON 255.085 40.235 255.085 40.215 255.050 40.215 ;
        RECT 255.085 40.215 257.595 40.235 ;
        RECT 247.835 40.210 251.180 40.215 ;
        POLYGON 247.840 40.210 248.010 40.210 248.010 40.190 ;
        RECT 248.010 40.200 251.180 40.210 ;
        POLYGON 251.180 40.215 251.345 40.215 251.180 40.200 ;
        POLYGON 255.050 40.215 255.050 40.200 255.025 40.200 ;
        RECT 255.050 40.200 257.595 40.215 ;
        RECT 248.010 40.190 251.065 40.200 ;
        POLYGON 251.065 40.200 251.175 40.200 251.065 40.190 ;
        POLYGON 255.025 40.200 255.025 40.190 255.005 40.190 ;
        RECT 255.025 40.190 257.595 40.200 ;
        POLYGON 248.010 40.190 248.095 40.190 248.095 40.185 ;
        RECT 248.095 40.185 250.435 40.190 ;
        RECT 241.010 40.130 244.020 40.185 ;
        POLYGON 241.010 40.130 241.025 40.130 241.025 40.115 ;
        RECT 241.025 40.115 244.020 40.130 ;
        RECT 232.650 40.030 237.335 40.115 ;
        POLYGON 237.335 40.115 237.410 40.030 237.335 40.030 ;
        POLYGON 241.025 40.115 241.130 40.115 241.130 40.030 ;
        RECT 241.130 40.050 244.020 40.115 ;
        POLYGON 244.020 40.185 244.260 40.050 244.020 40.050 ;
        POLYGON 248.100 40.185 248.295 40.185 248.295 40.170 ;
        RECT 248.295 40.170 250.435 40.185 ;
        POLYGON 248.370 40.170 248.645 40.170 248.645 40.160 ;
        RECT 248.645 40.160 250.435 40.170 ;
        POLYGON 250.435 40.190 251.065 40.190 250.435 40.160 ;
        POLYGON 255.005 40.190 255.005 40.160 254.955 40.160 ;
        RECT 255.005 40.160 257.595 40.190 ;
        POLYGON 248.660 40.160 248.940 40.160 248.940 40.150 ;
        RECT 248.940 40.150 249.695 40.160 ;
        POLYGON 249.695 40.160 250.365 40.160 249.695 40.150 ;
        POLYGON 254.955 40.160 254.955 40.150 254.935 40.150 ;
        RECT 254.955 40.150 257.595 40.160 ;
        POLYGON 254.935 40.150 254.935 40.110 254.865 40.110 ;
        RECT 254.935 40.110 257.595 40.150 ;
        POLYGON 254.865 40.110 254.865 40.065 254.770 40.065 ;
        RECT 254.865 40.065 257.595 40.110 ;
        POLYGON 254.770 40.065 254.770 40.055 254.755 40.055 ;
        RECT 254.770 40.055 257.595 40.065 ;
        POLYGON 254.755 40.055 254.755 40.050 254.745 40.050 ;
        RECT 254.755 40.050 257.595 40.055 ;
        POLYGON 257.595 40.275 257.850 40.275 257.595 40.050 ;
        POLYGON 260.855 40.275 260.855 40.200 260.795 40.200 ;
        RECT 260.855 40.200 264.420 40.275 ;
        POLYGON 264.420 40.730 264.720 40.730 264.420 40.200 ;
        POLYGON 269.610 40.730 269.610 40.250 269.420 40.250 ;
        RECT 269.610 40.250 277.205 40.730 ;
        POLYGON 269.420 40.250 269.420 40.200 269.395 40.200 ;
        RECT 269.420 40.200 277.205 40.250 ;
        POLYGON 260.795 40.200 260.795 40.090 260.695 40.090 ;
        RECT 260.795 40.095 264.355 40.200 ;
        POLYGON 264.355 40.200 264.420 40.200 264.355 40.095 ;
        POLYGON 269.395 40.195 269.395 40.140 269.370 40.140 ;
        RECT 269.395 40.185 277.205 40.200 ;
        POLYGON 277.205 41.495 277.455 41.495 277.205 40.185 ;
        POLYGON 287.645 41.480 287.645 40.220 287.580 40.220 ;
        RECT 287.645 40.220 303.120 41.495 ;
        RECT 269.395 40.140 277.040 40.185 ;
        POLYGON 269.370 40.140 269.370 40.095 269.350 40.095 ;
        RECT 269.370 40.095 277.040 40.140 ;
        RECT 260.795 40.090 264.105 40.095 ;
        POLYGON 260.695 40.090 260.695 40.050 260.660 40.050 ;
        RECT 260.695 40.050 264.105 40.090 ;
        RECT 241.130 40.030 244.260 40.050 ;
        RECT 232.650 40.020 237.410 40.030 ;
        RECT 210.290 40.015 225.225 40.020 ;
        POLYGON 225.225 40.020 225.230 40.015 225.225 40.015 ;
        POLYGON 232.650 40.020 232.655 40.020 232.655 40.015 ;
        RECT 232.655 40.015 237.410 40.020 ;
        RECT 210.290 39.710 225.230 40.015 ;
        POLYGON 225.230 40.015 225.390 39.710 225.230 39.710 ;
        POLYGON 232.655 40.015 232.880 40.015 232.880 39.710 ;
        RECT 232.880 39.870 237.410 40.015 ;
        POLYGON 237.410 40.030 237.555 39.870 237.410 39.870 ;
        POLYGON 241.130 40.030 241.315 40.030 241.315 39.885 ;
        RECT 241.315 39.960 244.260 40.030 ;
        POLYGON 244.260 40.050 244.425 39.960 244.260 39.960 ;
        POLYGON 254.745 40.050 254.745 39.960 254.570 39.960 ;
        RECT 254.745 39.960 257.415 40.050 ;
        RECT 241.315 39.955 244.425 39.960 ;
        POLYGON 244.425 39.960 244.435 39.955 244.425 39.955 ;
        POLYGON 254.570 39.960 254.570 39.955 254.560 39.955 ;
        RECT 254.570 39.955 257.415 39.960 ;
        RECT 241.315 39.885 244.440 39.955 ;
        POLYGON 254.560 39.955 254.560 39.950 254.550 39.950 ;
        RECT 254.560 39.950 257.415 39.955 ;
        POLYGON 241.315 39.885 241.330 39.885 241.330 39.870 ;
        RECT 241.330 39.870 244.440 39.885 ;
        RECT 232.880 39.750 237.555 39.870 ;
        POLYGON 237.555 39.870 237.670 39.750 237.555 39.750 ;
        POLYGON 241.330 39.870 241.480 39.870 241.480 39.760 ;
        RECT 241.480 39.760 244.440 39.870 ;
        POLYGON 241.480 39.760 241.490 39.760 241.490 39.750 ;
        RECT 241.490 39.755 244.440 39.760 ;
        POLYGON 244.440 39.950 244.840 39.755 244.440 39.755 ;
        POLYGON 254.550 39.950 254.550 39.900 254.455 39.900 ;
        RECT 254.550 39.910 257.415 39.950 ;
        POLYGON 257.415 40.050 257.595 40.050 257.415 39.910 ;
        POLYGON 260.660 40.050 260.660 39.910 260.530 39.910 ;
        RECT 260.660 39.910 264.105 40.050 ;
        RECT 254.550 39.900 257.345 39.910 ;
        POLYGON 254.455 39.900 254.455 39.795 254.230 39.795 ;
        RECT 254.455 39.850 257.345 39.900 ;
        POLYGON 257.345 39.910 257.415 39.910 257.345 39.850 ;
        POLYGON 260.530 39.910 260.530 39.850 260.475 39.850 ;
        RECT 260.530 39.850 264.105 39.910 ;
        RECT 254.455 39.795 257.165 39.850 ;
        POLYGON 254.230 39.795 254.230 39.770 254.185 39.770 ;
        RECT 254.230 39.770 257.165 39.795 ;
        POLYGON 254.185 39.770 254.185 39.755 254.155 39.755 ;
        RECT 254.185 39.755 257.165 39.770 ;
        RECT 241.490 39.750 244.840 39.755 ;
        RECT 232.880 39.710 237.670 39.750 ;
        RECT 210.290 39.495 225.390 39.710 ;
        POLYGON 225.390 39.710 225.510 39.495 225.390 39.495 ;
        POLYGON 232.880 39.710 232.910 39.710 232.910 39.670 ;
        RECT 232.910 39.705 237.670 39.710 ;
        POLYGON 237.670 39.750 237.715 39.705 237.670 39.705 ;
        POLYGON 241.490 39.750 241.555 39.750 241.555 39.705 ;
        RECT 241.555 39.725 244.840 39.750 ;
        POLYGON 244.840 39.755 244.900 39.725 244.840 39.725 ;
        POLYGON 254.155 39.755 254.155 39.725 254.090 39.725 ;
        RECT 254.155 39.725 257.165 39.755 ;
        RECT 241.555 39.705 244.900 39.725 ;
        RECT 232.910 39.670 237.715 39.705 ;
        POLYGON 232.910 39.670 232.970 39.670 232.970 39.580 ;
        RECT 232.970 39.580 237.715 39.670 ;
        POLYGON 232.970 39.580 233.035 39.580 233.035 39.495 ;
        RECT 233.035 39.495 237.715 39.580 ;
        POLYGON 237.715 39.705 237.910 39.495 237.715 39.495 ;
        POLYGON 241.555 39.705 241.710 39.705 241.710 39.595 ;
        RECT 241.710 39.695 244.900 39.705 ;
        POLYGON 244.900 39.725 244.955 39.695 244.900 39.695 ;
        POLYGON 254.090 39.725 254.090 39.695 254.030 39.695 ;
        RECT 254.090 39.705 257.165 39.725 ;
        POLYGON 257.165 39.850 257.345 39.850 257.165 39.705 ;
        POLYGON 260.475 39.850 260.475 39.790 260.420 39.790 ;
        RECT 260.475 39.790 264.105 39.850 ;
        POLYGON 260.420 39.790 260.420 39.745 260.385 39.745 ;
        RECT 260.420 39.745 264.105 39.790 ;
        POLYGON 260.385 39.745 260.385 39.705 260.350 39.705 ;
        RECT 260.385 39.705 264.105 39.745 ;
        RECT 254.090 39.695 256.880 39.705 ;
        RECT 241.710 39.635 244.955 39.695 ;
        POLYGON 244.955 39.695 245.090 39.635 244.955 39.635 ;
        POLYGON 254.030 39.695 254.030 39.645 253.925 39.645 ;
        RECT 254.030 39.645 256.880 39.695 ;
        POLYGON 253.925 39.645 253.925 39.635 253.900 39.635 ;
        RECT 253.925 39.635 256.880 39.645 ;
        RECT 241.710 39.595 245.095 39.635 ;
        POLYGON 241.710 39.595 241.850 39.595 241.850 39.495 ;
        RECT 241.850 39.560 245.095 39.595 ;
        POLYGON 245.095 39.635 245.265 39.560 245.095 39.560 ;
        POLYGON 253.900 39.635 253.900 39.580 253.790 39.580 ;
        RECT 253.900 39.580 256.880 39.635 ;
        POLYGON 253.790 39.580 253.790 39.560 253.740 39.560 ;
        RECT 253.790 39.560 256.880 39.580 ;
        RECT 241.850 39.495 245.265 39.560 ;
        POLYGON 245.265 39.560 245.395 39.495 245.265 39.495 ;
        POLYGON 253.740 39.560 253.740 39.530 253.670 39.530 ;
        RECT 253.740 39.530 256.880 39.560 ;
        POLYGON 253.670 39.530 253.670 39.495 253.590 39.495 ;
        RECT 253.670 39.495 256.880 39.530 ;
        POLYGON 256.880 39.705 257.165 39.705 256.880 39.495 ;
        POLYGON 260.350 39.705 260.350 39.495 260.155 39.495 ;
        RECT 260.350 39.685 264.105 39.705 ;
        POLYGON 264.105 40.095 264.355 40.095 264.105 39.685 ;
        POLYGON 269.350 40.095 269.350 39.690 269.170 39.690 ;
        RECT 269.350 39.690 277.040 40.095 ;
        RECT 260.350 39.495 263.975 39.685 ;
        POLYGON 263.975 39.685 264.105 39.685 263.975 39.495 ;
        POLYGON 269.170 39.685 269.170 39.500 269.085 39.500 ;
        RECT 269.170 39.500 277.040 39.690 ;
        POLYGON 277.040 40.185 277.205 40.185 277.040 39.505 ;
        POLYGON 287.580 40.185 287.580 39.540 287.545 39.540 ;
        RECT 287.580 39.540 303.120 40.220 ;
        RECT 269.085 39.495 277.040 39.500 ;
        RECT 182.060 39.335 197.810 39.495 ;
        RECT 161.675 39.320 164.520 39.335 ;
        RECT 117.510 39.305 158.170 39.320 ;
        POLYGON 158.170 39.320 158.210 39.320 158.170 39.305 ;
        POLYGON 161.645 39.320 161.645 39.305 161.625 39.305 ;
        RECT 161.645 39.305 164.520 39.320 ;
        RECT 117.510 39.265 158.025 39.305 ;
        POLYGON 117.510 39.265 117.515 39.265 117.515 39.260 ;
        RECT 117.515 39.260 158.025 39.265 ;
        RECT 58.745 38.160 115.350 39.260 ;
        POLYGON 115.350 39.260 115.885 38.160 115.350 38.160 ;
        POLYGON 117.515 39.260 117.520 39.260 117.520 39.190 ;
        RECT 117.520 39.250 158.025 39.260 ;
        POLYGON 158.025 39.305 158.170 39.305 158.025 39.250 ;
        POLYGON 161.625 39.305 161.625 39.280 161.585 39.280 ;
        RECT 161.625 39.280 164.520 39.305 ;
        POLYGON 161.585 39.280 161.585 39.250 161.540 39.250 ;
        RECT 161.585 39.250 164.520 39.280 ;
        RECT 117.520 39.220 157.950 39.250 ;
        POLYGON 157.950 39.250 158.025 39.250 157.950 39.220 ;
        POLYGON 161.540 39.250 161.540 39.220 161.500 39.220 ;
        RECT 161.540 39.220 164.520 39.250 ;
        RECT 117.520 39.155 157.695 39.220 ;
        POLYGON 117.520 39.155 117.525 39.155 117.525 39.120 ;
        RECT 117.525 39.135 157.695 39.155 ;
        POLYGON 157.695 39.220 157.950 39.220 157.695 39.135 ;
        POLYGON 161.500 39.220 161.500 39.210 161.485 39.210 ;
        RECT 161.500 39.210 164.520 39.220 ;
        POLYGON 161.485 39.210 161.485 39.135 161.370 39.135 ;
        RECT 161.485 39.135 164.520 39.210 ;
        RECT 117.525 39.120 157.640 39.135 ;
        POLYGON 157.640 39.135 157.695 39.135 157.640 39.120 ;
        POLYGON 161.370 39.135 161.370 39.120 161.350 39.120 ;
        RECT 161.370 39.120 164.520 39.135 ;
        RECT 117.525 39.080 157.440 39.120 ;
        POLYGON 117.525 39.080 117.535 39.080 117.535 38.980 ;
        RECT 117.535 39.060 157.440 39.080 ;
        POLYGON 157.440 39.120 157.640 39.120 157.440 39.060 ;
        POLYGON 161.350 39.120 161.350 39.065 161.265 39.065 ;
        RECT 161.350 39.065 164.520 39.120 ;
        POLYGON 161.265 39.065 161.265 39.060 161.260 39.060 ;
        RECT 161.265 39.060 164.520 39.065 ;
        RECT 117.535 39.020 157.270 39.060 ;
        POLYGON 157.270 39.060 157.440 39.060 157.270 39.020 ;
        POLYGON 161.260 39.060 161.260 39.055 161.250 39.055 ;
        RECT 161.260 39.055 164.520 39.060 ;
        POLYGON 161.250 39.055 161.250 39.020 161.195 39.020 ;
        RECT 161.250 39.020 164.520 39.055 ;
        RECT 117.535 39.000 157.190 39.020 ;
        POLYGON 157.190 39.020 157.270 39.020 157.190 39.000 ;
        POLYGON 161.195 39.020 161.195 39.000 161.160 39.000 ;
        RECT 161.195 39.000 164.520 39.020 ;
        RECT 117.535 38.980 157.105 39.000 ;
        POLYGON 157.105 39.000 157.190 39.000 157.105 38.980 ;
        POLYGON 161.160 39.000 161.160 38.980 161.130 38.980 ;
        RECT 161.160 38.980 164.520 39.000 ;
        RECT 117.535 38.950 156.930 38.980 ;
        POLYGON 156.930 38.980 157.100 38.980 156.930 38.950 ;
        POLYGON 161.130 38.980 161.130 38.950 161.080 38.950 ;
        RECT 161.130 38.950 164.520 38.980 ;
        RECT 117.535 38.920 156.660 38.950 ;
        POLYGON 117.535 38.920 117.580 38.920 117.580 38.345 ;
        RECT 117.580 38.910 156.660 38.920 ;
        POLYGON 156.660 38.950 156.930 38.950 156.660 38.910 ;
        POLYGON 161.080 38.950 161.080 38.910 161.015 38.910 ;
        RECT 161.080 38.910 164.520 38.950 ;
        RECT 117.580 38.900 156.560 38.910 ;
        POLYGON 156.560 38.910 156.660 38.910 156.560 38.900 ;
        POLYGON 161.015 38.910 161.015 38.900 161.000 38.900 ;
        RECT 161.015 38.900 164.520 38.910 ;
        RECT 117.580 38.890 156.490 38.900 ;
        POLYGON 156.490 38.900 156.555 38.900 156.490 38.890 ;
        POLYGON 161.000 38.900 161.000 38.890 160.985 38.890 ;
        RECT 161.000 38.890 164.520 38.900 ;
        RECT 117.580 38.880 156.375 38.890 ;
        POLYGON 156.375 38.890 156.485 38.890 156.375 38.880 ;
        POLYGON 160.985 38.890 160.985 38.880 160.965 38.880 ;
        RECT 160.985 38.880 164.520 38.890 ;
        RECT 117.580 38.855 156.065 38.880 ;
        POLYGON 156.065 38.880 156.375 38.880 156.065 38.855 ;
        POLYGON 160.965 38.880 160.965 38.855 160.925 38.855 ;
        RECT 160.965 38.855 164.520 38.880 ;
        RECT 117.580 38.845 155.690 38.855 ;
        RECT 117.580 38.830 153.400 38.845 ;
        POLYGON 153.400 38.845 153.420 38.845 153.420 38.840 ;
        RECT 153.420 38.840 155.690 38.845 ;
        POLYGON 155.690 38.855 155.985 38.855 155.690 38.840 ;
        POLYGON 160.925 38.855 160.925 38.840 160.900 38.840 ;
        RECT 160.925 38.840 164.520 38.855 ;
        POLYGON 153.400 38.840 153.410 38.830 153.400 38.830 ;
        POLYGON 153.425 38.840 153.735 38.840 153.735 38.830 ;
        RECT 153.735 38.830 155.370 38.840 ;
        POLYGON 155.370 38.840 155.685 38.840 155.370 38.830 ;
        POLYGON 160.900 38.840 160.900 38.830 160.885 38.830 ;
        RECT 160.900 38.830 164.520 38.840 ;
        RECT 117.580 38.800 153.410 38.830 ;
        POLYGON 154.000 38.830 154.305 38.830 154.305 38.825 ;
        RECT 154.305 38.825 154.915 38.830 ;
        POLYGON 154.915 38.830 155.370 38.830 154.915 38.825 ;
        POLYGON 160.885 38.830 160.885 38.825 160.875 38.825 ;
        RECT 160.885 38.825 164.520 38.830 ;
        POLYGON 153.410 38.825 153.425 38.800 153.410 38.800 ;
        POLYGON 160.875 38.825 160.875 38.800 160.835 38.800 ;
        RECT 160.875 38.805 164.520 38.825 ;
        POLYGON 164.520 39.335 165.045 39.335 164.520 38.805 ;
        POLYGON 168.885 39.335 168.885 39.275 168.840 39.275 ;
        RECT 168.885 39.275 173.920 39.335 ;
        POLYGON 168.840 39.275 168.840 39.210 168.795 39.210 ;
        RECT 168.840 39.210 173.920 39.275 ;
        POLYGON 168.795 39.210 168.795 39.110 168.730 39.110 ;
        RECT 168.795 39.110 173.920 39.210 ;
        POLYGON 168.730 39.110 168.730 39.045 168.685 39.045 ;
        RECT 168.730 39.090 173.920 39.110 ;
        POLYGON 173.920 39.335 174.025 39.335 173.920 39.090 ;
        POLYGON 182.015 39.335 182.015 39.090 181.955 39.090 ;
        RECT 182.015 39.090 197.810 39.335 ;
        RECT 168.730 39.045 173.390 39.090 ;
        POLYGON 168.685 39.045 168.685 38.865 168.555 38.865 ;
        RECT 168.685 38.865 173.390 39.045 ;
        POLYGON 168.555 38.865 168.555 38.805 168.510 38.805 ;
        RECT 168.555 38.805 173.390 38.865 ;
        RECT 160.875 38.800 164.000 38.805 ;
        RECT 117.580 38.765 153.425 38.800 ;
        POLYGON 153.425 38.800 153.445 38.765 153.425 38.765 ;
        RECT 117.580 38.755 153.445 38.765 ;
        POLYGON 160.830 38.800 160.830 38.760 160.770 38.760 ;
        RECT 160.830 38.760 164.000 38.800 ;
        POLYGON 153.445 38.760 153.450 38.755 153.445 38.755 ;
        POLYGON 160.770 38.760 160.770 38.755 160.760 38.755 ;
        RECT 160.770 38.755 164.000 38.760 ;
        RECT 117.580 38.700 153.450 38.755 ;
        POLYGON 160.760 38.755 160.760 38.750 160.755 38.750 ;
        RECT 160.760 38.750 164.000 38.755 ;
        POLYGON 153.450 38.750 153.480 38.700 153.450 38.700 ;
        POLYGON 160.755 38.750 160.755 38.700 160.665 38.700 ;
        RECT 160.755 38.700 164.000 38.750 ;
        RECT 117.580 38.555 153.480 38.700 ;
        POLYGON 153.480 38.700 153.560 38.555 153.480 38.555 ;
        RECT 117.580 38.485 153.560 38.555 ;
        POLYGON 160.660 38.700 160.660 38.550 160.390 38.550 ;
        RECT 160.660 38.550 164.000 38.700 ;
        POLYGON 153.560 38.550 153.600 38.485 153.560 38.485 ;
        POLYGON 160.390 38.550 160.390 38.485 160.275 38.485 ;
        RECT 160.390 38.485 164.000 38.550 ;
        RECT 117.580 38.440 153.600 38.485 ;
        POLYGON 153.600 38.485 153.625 38.440 153.600 38.440 ;
        POLYGON 160.275 38.485 160.275 38.440 160.185 38.440 ;
        RECT 160.275 38.440 164.000 38.485 ;
        RECT 117.580 38.430 153.625 38.440 ;
        POLYGON 153.625 38.440 153.630 38.430 153.625 38.430 ;
        POLYGON 160.185 38.440 160.185 38.430 160.160 38.430 ;
        RECT 160.185 38.430 164.000 38.440 ;
        RECT 117.580 38.320 153.630 38.430 ;
        POLYGON 153.630 38.430 153.690 38.320 153.630 38.320 ;
        POLYGON 117.580 38.320 117.590 38.320 117.590 38.205 ;
        RECT 117.590 38.275 153.690 38.320 ;
        POLYGON 160.160 38.430 160.160 38.315 159.930 38.315 ;
        RECT 160.160 38.325 164.000 38.430 ;
        POLYGON 164.000 38.805 164.520 38.805 164.000 38.325 ;
        POLYGON 168.510 38.805 168.510 38.665 168.405 38.665 ;
        RECT 168.510 38.665 173.390 38.805 ;
        POLYGON 168.405 38.665 168.405 38.570 168.335 38.570 ;
        RECT 168.405 38.570 173.390 38.665 ;
        POLYGON 168.335 38.570 168.335 38.465 168.255 38.465 ;
        RECT 168.335 38.465 173.390 38.570 ;
        POLYGON 168.255 38.465 168.255 38.445 168.240 38.445 ;
        RECT 168.255 38.445 173.390 38.465 ;
        POLYGON 168.240 38.445 168.240 38.330 168.145 38.330 ;
        RECT 168.240 38.330 173.390 38.445 ;
        RECT 160.160 38.315 163.940 38.325 ;
        POLYGON 153.690 38.315 153.715 38.275 153.690 38.275 ;
        POLYGON 159.925 38.315 159.925 38.275 159.850 38.275 ;
        RECT 159.925 38.275 163.940 38.315 ;
        POLYGON 163.940 38.325 164.000 38.325 163.940 38.275 ;
        POLYGON 168.145 38.325 168.145 38.280 168.105 38.280 ;
        RECT 168.145 38.280 173.390 38.330 ;
        RECT 117.590 38.230 153.715 38.275 ;
        POLYGON 153.715 38.275 153.740 38.230 153.715 38.230 ;
        POLYGON 159.850 38.275 159.850 38.230 159.765 38.230 ;
        RECT 159.850 38.230 163.350 38.275 ;
        RECT 117.590 38.205 153.740 38.230 ;
        POLYGON 159.765 38.230 159.765 38.225 159.755 38.225 ;
        RECT 159.765 38.225 163.350 38.230 ;
        POLYGON 153.740 38.225 153.755 38.205 153.740 38.205 ;
        RECT 58.745 38.055 115.885 38.160 ;
        POLYGON 58.745 38.055 59.505 38.055 59.505 36.635 ;
        RECT 59.505 38.010 115.885 38.055 ;
        POLYGON 115.885 38.160 115.955 38.010 115.885 38.010 ;
        RECT 117.590 38.155 153.755 38.205 ;
        POLYGON 159.755 38.225 159.755 38.200 159.700 38.200 ;
        RECT 159.755 38.200 163.350 38.225 ;
        POLYGON 117.590 38.155 117.600 38.155 117.600 38.065 ;
        RECT 117.600 38.140 153.755 38.155 ;
        POLYGON 153.755 38.200 153.790 38.140 153.755 38.140 ;
        RECT 117.600 38.095 153.790 38.140 ;
        POLYGON 159.695 38.200 159.695 38.135 159.555 38.135 ;
        RECT 159.695 38.135 163.350 38.200 ;
        POLYGON 153.790 38.135 153.815 38.095 153.790 38.095 ;
        POLYGON 159.555 38.135 159.555 38.095 159.470 38.095 ;
        RECT 159.555 38.095 163.350 38.135 ;
        RECT 117.600 38.085 153.815 38.095 ;
        POLYGON 153.815 38.095 153.820 38.085 153.815 38.085 ;
        POLYGON 159.470 38.095 159.470 38.085 159.445 38.085 ;
        RECT 159.470 38.085 163.350 38.095 ;
        RECT 117.600 38.040 153.820 38.085 ;
        POLYGON 153.820 38.085 153.845 38.040 153.820 38.040 ;
        RECT 117.600 38.010 153.845 38.040 ;
        POLYGON 159.445 38.085 159.445 38.035 159.340 38.035 ;
        RECT 159.445 38.035 163.350 38.085 ;
        RECT 59.505 37.750 115.955 38.010 ;
        POLYGON 115.955 38.010 116.095 37.750 115.955 37.750 ;
        POLYGON 117.600 38.010 117.620 38.010 117.620 37.780 ;
        RECT 117.620 37.975 153.845 38.010 ;
        POLYGON 153.845 38.035 153.880 37.975 153.845 37.975 ;
        POLYGON 159.340 38.035 159.340 37.975 159.210 37.975 ;
        RECT 159.340 37.975 163.350 38.035 ;
        RECT 117.620 37.940 153.880 37.975 ;
        POLYGON 159.210 37.975 159.210 37.970 159.200 37.970 ;
        RECT 159.210 37.970 163.350 37.975 ;
        POLYGON 153.880 37.970 153.900 37.940 153.880 37.940 ;
        RECT 117.620 37.915 153.900 37.940 ;
        POLYGON 159.200 37.970 159.200 37.935 159.125 37.935 ;
        RECT 159.200 37.935 163.350 37.970 ;
        POLYGON 153.900 37.935 153.915 37.915 153.900 37.915 ;
        POLYGON 159.125 37.935 159.125 37.915 159.085 37.915 ;
        RECT 159.125 37.915 163.350 37.935 ;
        RECT 117.620 37.805 153.915 37.915 ;
        POLYGON 153.915 37.915 153.975 37.805 153.915 37.805 ;
        POLYGON 159.085 37.915 159.085 37.805 158.820 37.805 ;
        RECT 159.085 37.805 163.350 37.915 ;
        RECT 117.620 37.795 153.975 37.805 ;
        POLYGON 153.975 37.805 153.980 37.795 153.975 37.795 ;
        RECT 117.620 37.785 153.980 37.795 ;
        POLYGON 158.820 37.805 158.820 37.790 158.785 37.790 ;
        RECT 158.820 37.790 163.350 37.805 ;
        POLYGON 153.980 37.790 153.985 37.785 153.980 37.785 ;
        RECT 117.620 37.760 153.985 37.785 ;
        POLYGON 158.780 37.790 158.780 37.780 158.755 37.780 ;
        RECT 158.780 37.780 163.350 37.790 ;
        POLYGON 163.350 38.275 163.940 38.275 163.350 37.780 ;
        POLYGON 168.105 38.275 168.105 38.210 168.050 38.210 ;
        RECT 168.105 38.210 173.390 38.280 ;
        POLYGON 168.050 38.210 168.050 38.080 167.950 38.080 ;
        RECT 168.050 38.080 173.390 38.210 ;
        POLYGON 167.950 38.080 167.950 38.040 167.920 38.040 ;
        RECT 167.950 38.040 173.390 38.080 ;
        POLYGON 167.920 38.040 167.920 37.955 167.845 37.955 ;
        RECT 167.920 38.000 173.390 38.040 ;
        POLYGON 173.390 39.090 173.920 39.090 173.390 38.000 ;
        POLYGON 181.955 39.085 181.955 38.895 181.910 38.895 ;
        RECT 181.955 38.895 197.810 39.090 ;
        POLYGON 181.910 38.895 181.910 38.085 181.675 38.085 ;
        RECT 181.910 38.085 197.810 38.895 ;
        POLYGON 181.675 38.085 181.675 38.000 181.650 38.000 ;
        RECT 181.675 38.000 197.810 38.085 ;
        RECT 167.920 37.955 173.185 38.000 ;
        POLYGON 167.845 37.955 167.845 37.780 167.695 37.780 ;
        RECT 167.845 37.780 173.185 37.955 ;
        POLYGON 153.985 37.780 154.000 37.760 153.985 37.760 ;
        RECT 117.620 37.750 154.000 37.760 ;
        POLYGON 158.755 37.780 158.755 37.755 158.690 37.755 ;
        RECT 158.755 37.755 163.105 37.780 ;
        RECT 59.505 36.785 116.095 37.750 ;
        POLYGON 116.095 37.750 116.600 36.785 116.095 36.785 ;
        POLYGON 117.620 37.750 117.640 37.750 117.640 37.500 ;
        RECT 117.640 37.740 154.000 37.750 ;
        POLYGON 154.000 37.755 154.010 37.740 154.000 37.740 ;
        POLYGON 158.690 37.755 158.690 37.740 158.655 37.740 ;
        RECT 158.690 37.740 163.105 37.755 ;
        RECT 117.640 37.680 154.010 37.740 ;
        POLYGON 158.655 37.740 158.655 37.735 158.645 37.735 ;
        RECT 158.655 37.735 163.105 37.740 ;
        POLYGON 154.010 37.735 154.045 37.680 154.010 37.680 ;
        RECT 117.640 37.625 154.045 37.680 ;
        POLYGON 158.645 37.735 158.645 37.675 158.500 37.675 ;
        RECT 158.645 37.675 163.105 37.735 ;
        POLYGON 154.045 37.675 154.075 37.625 154.045 37.625 ;
        POLYGON 158.500 37.675 158.500 37.625 158.365 37.625 ;
        RECT 158.500 37.625 163.105 37.675 ;
        RECT 117.640 37.585 154.075 37.625 ;
        POLYGON 154.075 37.625 154.095 37.585 154.075 37.585 ;
        POLYGON 158.365 37.625 158.365 37.585 158.255 37.585 ;
        RECT 158.365 37.595 163.105 37.625 ;
        POLYGON 163.105 37.780 163.350 37.780 163.105 37.595 ;
        POLYGON 167.695 37.780 167.695 37.690 167.620 37.690 ;
        RECT 167.695 37.690 173.185 37.780 ;
        POLYGON 167.620 37.690 167.620 37.595 167.535 37.595 ;
        RECT 167.620 37.625 173.185 37.690 ;
        POLYGON 173.185 38.000 173.390 38.000 173.185 37.625 ;
        POLYGON 181.650 37.995 181.650 37.855 181.610 37.855 ;
        RECT 181.650 37.855 197.810 38.000 ;
        POLYGON 181.610 37.855 181.610 37.645 181.545 37.645 ;
        RECT 181.610 37.645 197.810 37.855 ;
        POLYGON 181.545 37.645 181.545 37.630 181.540 37.630 ;
        RECT 181.545 37.630 197.810 37.645 ;
        RECT 167.620 37.595 172.905 37.625 ;
        RECT 158.365 37.585 162.920 37.595 ;
        RECT 117.640 37.580 154.095 37.585 ;
        POLYGON 154.095 37.585 154.100 37.580 154.095 37.580 ;
        RECT 117.640 37.570 154.100 37.580 ;
        POLYGON 158.255 37.585 158.255 37.575 158.230 37.575 ;
        RECT 158.255 37.575 162.920 37.585 ;
        POLYGON 154.100 37.575 154.105 37.570 154.100 37.570 ;
        POLYGON 158.230 37.575 158.230 37.570 158.210 37.570 ;
        RECT 158.230 37.570 162.920 37.575 ;
        RECT 117.640 37.560 154.105 37.570 ;
        POLYGON 158.210 37.570 158.210 37.565 158.195 37.565 ;
        RECT 158.210 37.565 162.920 37.570 ;
        POLYGON 154.105 37.565 154.110 37.560 154.105 37.560 ;
        RECT 117.640 37.535 154.110 37.560 ;
        POLYGON 158.195 37.565 158.195 37.555 158.170 37.555 ;
        RECT 158.195 37.555 162.920 37.565 ;
        POLYGON 154.110 37.555 154.125 37.535 154.110 37.535 ;
        RECT 117.640 37.525 154.125 37.535 ;
        POLYGON 158.170 37.555 158.170 37.530 158.090 37.530 ;
        RECT 158.170 37.530 162.920 37.555 ;
        POLYGON 154.125 37.530 154.130 37.525 154.125 37.525 ;
        POLYGON 158.090 37.530 158.090 37.525 158.075 37.525 ;
        RECT 158.090 37.525 162.920 37.530 ;
        RECT 117.640 37.515 154.130 37.525 ;
        POLYGON 154.130 37.525 154.135 37.515 154.130 37.515 ;
        RECT 117.640 37.495 154.135 37.515 ;
        POLYGON 158.075 37.525 158.075 37.510 158.025 37.510 ;
        RECT 158.075 37.510 162.920 37.525 ;
        POLYGON 117.640 37.495 117.645 37.495 117.645 37.430 ;
        RECT 117.645 37.490 154.135 37.495 ;
        POLYGON 154.135 37.510 154.150 37.490 154.135 37.490 ;
        POLYGON 158.025 37.510 158.025 37.490 157.965 37.490 ;
        RECT 158.025 37.490 162.920 37.510 ;
        RECT 117.645 37.450 154.150 37.490 ;
        POLYGON 154.150 37.490 154.170 37.450 154.150 37.450 ;
        RECT 117.645 37.435 154.170 37.450 ;
        POLYGON 157.950 37.490 157.950 37.445 157.790 37.445 ;
        RECT 157.950 37.455 162.920 37.490 ;
        POLYGON 162.920 37.595 163.105 37.595 162.920 37.455 ;
        POLYGON 167.535 37.590 167.535 37.535 167.485 37.535 ;
        RECT 167.535 37.535 172.905 37.595 ;
        POLYGON 167.485 37.535 167.485 37.455 167.410 37.455 ;
        RECT 167.485 37.455 172.905 37.535 ;
        RECT 157.950 37.445 162.740 37.455 ;
        POLYGON 154.170 37.445 154.180 37.435 154.170 37.435 ;
        RECT 117.645 37.425 154.180 37.435 ;
        POLYGON 157.790 37.445 157.790 37.430 157.735 37.430 ;
        RECT 157.790 37.430 162.740 37.445 ;
        POLYGON 154.180 37.430 154.185 37.425 154.180 37.425 ;
        POLYGON 157.735 37.430 157.735 37.425 157.720 37.425 ;
        RECT 157.735 37.425 162.740 37.430 ;
        RECT 117.645 37.415 154.185 37.425 ;
        POLYGON 157.720 37.425 157.720 37.420 157.700 37.420 ;
        RECT 157.720 37.420 162.740 37.425 ;
        POLYGON 154.185 37.420 154.190 37.415 154.185 37.415 ;
        POLYGON 117.645 37.415 117.690 37.415 117.690 36.795 ;
        RECT 117.690 37.380 154.190 37.415 ;
        POLYGON 157.695 37.420 157.695 37.410 157.640 37.410 ;
        RECT 157.695 37.410 162.740 37.420 ;
        POLYGON 154.190 37.410 154.210 37.380 154.190 37.380 ;
        POLYGON 157.640 37.410 157.640 37.380 157.505 37.380 ;
        RECT 157.640 37.380 162.740 37.410 ;
        RECT 117.690 37.370 154.210 37.380 ;
        POLYGON 157.505 37.380 157.505 37.375 157.485 37.375 ;
        RECT 157.505 37.375 162.740 37.380 ;
        POLYGON 154.210 37.375 154.215 37.370 154.210 37.370 ;
        RECT 117.690 37.335 154.215 37.370 ;
        POLYGON 157.485 37.375 157.485 37.365 157.440 37.365 ;
        RECT 157.485 37.365 162.740 37.375 ;
        POLYGON 154.215 37.365 154.235 37.335 154.215 37.335 ;
        POLYGON 157.430 37.365 157.430 37.335 157.270 37.335 ;
        RECT 157.430 37.335 162.740 37.365 ;
        RECT 117.690 37.325 154.235 37.335 ;
        POLYGON 157.265 37.335 157.265 37.330 157.230 37.330 ;
        RECT 157.265 37.330 162.740 37.335 ;
        POLYGON 154.235 37.330 154.240 37.325 154.235 37.325 ;
        POLYGON 157.230 37.330 157.230 37.325 157.190 37.325 ;
        RECT 157.230 37.325 162.740 37.330 ;
        POLYGON 162.740 37.455 162.920 37.455 162.740 37.325 ;
        POLYGON 167.410 37.455 167.410 37.415 167.375 37.415 ;
        RECT 167.410 37.415 172.905 37.455 ;
        POLYGON 167.375 37.415 167.375 37.325 167.290 37.325 ;
        RECT 167.375 37.325 172.905 37.415 ;
        RECT 117.690 37.315 154.240 37.325 ;
        POLYGON 154.240 37.325 154.245 37.315 154.240 37.315 ;
        POLYGON 157.190 37.325 157.190 37.315 157.145 37.315 ;
        RECT 157.190 37.315 162.120 37.325 ;
        RECT 117.690 37.295 154.245 37.315 ;
        POLYGON 157.145 37.315 157.145 37.310 157.100 37.310 ;
        RECT 157.145 37.310 162.120 37.315 ;
        POLYGON 154.245 37.310 154.255 37.295 154.245 37.295 ;
        POLYGON 157.095 37.310 157.095 37.295 156.970 37.295 ;
        RECT 157.095 37.295 162.120 37.310 ;
        RECT 117.690 37.290 154.255 37.295 ;
        POLYGON 154.255 37.295 154.260 37.290 154.255 37.290 ;
        POLYGON 156.970 37.295 156.970 37.290 156.930 37.290 ;
        RECT 156.970 37.290 162.120 37.295 ;
        RECT 117.690 37.270 154.260 37.290 ;
        POLYGON 154.260 37.290 154.270 37.270 154.260 37.270 ;
        POLYGON 156.925 37.290 156.925 37.280 156.845 37.280 ;
        RECT 156.925 37.280 162.120 37.290 ;
        POLYGON 156.845 37.280 156.845 37.270 156.720 37.270 ;
        RECT 156.845 37.270 162.120 37.280 ;
        RECT 117.690 37.260 154.270 37.270 ;
        POLYGON 156.720 37.270 156.720 37.265 156.660 37.265 ;
        RECT 156.720 37.265 162.120 37.270 ;
        POLYGON 154.270 37.265 154.275 37.260 154.270 37.260 ;
        RECT 117.690 37.245 154.275 37.260 ;
        POLYGON 156.660 37.265 156.660 37.255 156.560 37.255 ;
        RECT 156.660 37.255 162.120 37.265 ;
        POLYGON 154.275 37.255 154.285 37.245 154.275 37.245 ;
        POLYGON 156.555 37.255 156.555 37.250 156.525 37.250 ;
        RECT 156.555 37.250 162.120 37.255 ;
        POLYGON 156.485 37.250 156.485 37.245 156.375 37.245 ;
        RECT 156.485 37.245 162.120 37.250 ;
        RECT 117.690 37.235 154.285 37.245 ;
        POLYGON 156.370 37.245 156.370 37.240 156.305 37.240 ;
        RECT 156.370 37.240 162.120 37.245 ;
        POLYGON 154.285 37.240 154.290 37.235 154.285 37.235 ;
        POLYGON 156.305 37.240 156.305 37.235 156.235 37.235 ;
        RECT 156.305 37.235 162.120 37.240 ;
        RECT 117.690 37.225 154.290 37.235 ;
        POLYGON 156.235 37.235 156.235 37.230 156.170 37.230 ;
        RECT 156.235 37.230 162.120 37.235 ;
        POLYGON 154.290 37.230 154.295 37.225 154.290 37.225 ;
        POLYGON 156.060 37.230 156.060 37.225 155.985 37.225 ;
        RECT 156.060 37.225 162.120 37.230 ;
        RECT 117.690 37.215 154.295 37.225 ;
        POLYGON 155.985 37.225 155.985 37.220 155.690 37.220 ;
        RECT 155.985 37.220 162.120 37.225 ;
        POLYGON 154.295 37.220 154.300 37.215 154.295 37.215 ;
        POLYGON 155.685 37.220 155.685 37.215 155.530 37.215 ;
        RECT 155.685 37.215 162.120 37.220 ;
        RECT 117.690 37.205 154.300 37.215 ;
        POLYGON 155.530 37.215 155.530 37.210 155.370 37.210 ;
        RECT 155.530 37.210 162.120 37.215 ;
        POLYGON 154.300 37.210 154.305 37.205 154.300 37.205 ;
        POLYGON 155.355 37.210 155.355 37.205 154.855 37.205 ;
        RECT 155.355 37.205 162.120 37.210 ;
        RECT 117.690 36.905 162.120 37.205 ;
        POLYGON 162.120 37.325 162.740 37.325 162.120 36.905 ;
        POLYGON 167.290 37.325 167.290 37.155 167.135 37.155 ;
        RECT 167.290 37.155 172.905 37.325 ;
        POLYGON 167.135 37.155 167.135 37.125 167.110 37.125 ;
        RECT 167.135 37.125 172.905 37.155 ;
        POLYGON 167.110 37.125 167.110 37.040 167.030 37.040 ;
        RECT 167.110 37.105 172.905 37.125 ;
        POLYGON 172.905 37.625 173.185 37.625 172.905 37.105 ;
        POLYGON 181.540 37.625 181.540 37.105 181.360 37.105 ;
        RECT 181.540 37.215 197.810 37.630 ;
        POLYGON 197.810 39.495 198.000 39.495 197.810 37.215 ;
        POLYGON 210.290 39.495 210.395 39.495 210.395 39.270 ;
        RECT 210.395 39.270 225.510 39.495 ;
        POLYGON 210.395 39.270 210.730 39.270 210.730 38.585 ;
        RECT 210.730 39.165 225.510 39.270 ;
        POLYGON 225.510 39.495 225.700 39.165 225.510 39.165 ;
        POLYGON 233.035 39.495 233.300 39.495 233.300 39.165 ;
        RECT 233.300 39.280 237.910 39.495 ;
        POLYGON 237.910 39.495 238.120 39.280 237.910 39.280 ;
        POLYGON 241.850 39.495 242.160 39.495 242.160 39.280 ;
        RECT 242.160 39.455 245.395 39.495 ;
        POLYGON 245.395 39.495 245.495 39.455 245.395 39.455 ;
        POLYGON 253.590 39.495 253.590 39.460 253.505 39.460 ;
        RECT 253.590 39.460 256.720 39.495 ;
        POLYGON 253.505 39.460 253.505 39.455 253.495 39.455 ;
        RECT 253.505 39.455 256.720 39.460 ;
        RECT 242.160 39.385 245.495 39.455 ;
        POLYGON 245.495 39.455 245.665 39.385 245.495 39.385 ;
        POLYGON 253.495 39.455 253.495 39.420 253.420 39.420 ;
        RECT 253.495 39.420 256.720 39.455 ;
        POLYGON 253.415 39.420 253.415 39.385 253.335 39.385 ;
        RECT 253.415 39.385 256.720 39.420 ;
        RECT 242.160 39.330 245.665 39.385 ;
        POLYGON 245.665 39.385 245.815 39.330 245.665 39.330 ;
        POLYGON 253.335 39.385 253.335 39.340 253.235 39.340 ;
        RECT 253.335 39.375 256.720 39.385 ;
        POLYGON 256.720 39.495 256.880 39.495 256.720 39.375 ;
        POLYGON 260.155 39.495 260.155 39.470 260.130 39.470 ;
        RECT 260.155 39.470 263.820 39.495 ;
        POLYGON 260.130 39.470 260.130 39.385 260.055 39.385 ;
        RECT 260.130 39.385 263.820 39.470 ;
        POLYGON 260.055 39.385 260.055 39.375 260.045 39.375 ;
        RECT 260.055 39.375 263.820 39.385 ;
        RECT 253.335 39.340 256.255 39.375 ;
        POLYGON 253.235 39.340 253.235 39.330 253.205 39.330 ;
        RECT 253.235 39.330 256.255 39.340 ;
        RECT 242.160 39.280 245.815 39.330 ;
        POLYGON 245.815 39.330 245.940 39.280 245.815 39.280 ;
        POLYGON 253.205 39.330 253.205 39.315 253.165 39.315 ;
        RECT 253.205 39.315 256.255 39.330 ;
        POLYGON 253.165 39.315 253.165 39.280 253.080 39.280 ;
        RECT 253.165 39.280 256.255 39.315 ;
        RECT 233.300 39.265 238.120 39.280 ;
        POLYGON 238.120 39.280 238.135 39.265 238.120 39.265 ;
        POLYGON 242.160 39.280 242.185 39.280 242.185 39.265 ;
        RECT 242.185 39.265 245.940 39.280 ;
        RECT 233.300 39.215 238.135 39.265 ;
        POLYGON 238.135 39.265 238.190 39.215 238.135 39.215 ;
        POLYGON 242.185 39.265 242.270 39.265 242.270 39.215 ;
        RECT 242.270 39.260 245.940 39.265 ;
        POLYGON 245.940 39.280 245.995 39.260 245.940 39.260 ;
        POLYGON 253.080 39.280 253.080 39.260 253.030 39.260 ;
        RECT 253.080 39.260 256.255 39.280 ;
        RECT 242.270 39.215 245.995 39.260 ;
        RECT 233.300 39.165 238.190 39.215 ;
        RECT 210.730 38.930 225.700 39.165 ;
        POLYGON 225.700 39.165 225.835 38.930 225.700 38.930 ;
        POLYGON 233.300 39.165 233.475 39.165 233.475 38.945 ;
        RECT 233.475 39.095 238.190 39.165 ;
        POLYGON 238.190 39.215 238.320 39.095 238.190 39.095 ;
        POLYGON 242.270 39.215 242.380 39.215 242.380 39.150 ;
        RECT 242.380 39.180 245.995 39.215 ;
        POLYGON 245.995 39.260 246.235 39.180 245.995 39.180 ;
        POLYGON 253.030 39.260 253.030 39.240 252.980 39.240 ;
        RECT 253.030 39.240 256.255 39.260 ;
        POLYGON 252.970 39.240 252.970 39.230 252.955 39.230 ;
        RECT 252.970 39.230 256.255 39.240 ;
        POLYGON 252.955 39.230 252.955 39.215 252.905 39.215 ;
        RECT 252.955 39.215 256.255 39.230 ;
        POLYGON 252.905 39.215 252.905 39.180 252.805 39.180 ;
        RECT 252.905 39.180 256.255 39.215 ;
        RECT 242.380 39.175 246.235 39.180 ;
        POLYGON 246.235 39.180 246.245 39.175 246.235 39.175 ;
        POLYGON 252.805 39.180 252.805 39.175 252.795 39.175 ;
        RECT 252.805 39.175 256.255 39.180 ;
        RECT 242.380 39.155 246.245 39.175 ;
        POLYGON 246.245 39.175 246.310 39.155 246.245 39.155 ;
        POLYGON 252.795 39.175 252.795 39.165 252.765 39.165 ;
        RECT 252.795 39.165 256.255 39.175 ;
        POLYGON 252.760 39.165 252.760 39.155 252.725 39.155 ;
        RECT 252.760 39.155 256.255 39.165 ;
        RECT 242.380 39.150 246.310 39.155 ;
        POLYGON 242.385 39.150 242.440 39.150 242.440 39.115 ;
        RECT 242.440 39.115 246.310 39.150 ;
        POLYGON 242.440 39.115 242.470 39.115 242.470 39.095 ;
        RECT 242.470 39.110 246.310 39.115 ;
        POLYGON 246.310 39.155 246.470 39.110 246.310 39.110 ;
        POLYGON 252.725 39.155 252.725 39.150 252.705 39.150 ;
        RECT 252.725 39.150 256.255 39.155 ;
        POLYGON 252.705 39.150 252.705 39.145 252.700 39.145 ;
        RECT 252.705 39.145 256.255 39.150 ;
        POLYGON 252.700 39.145 252.700 39.125 252.635 39.125 ;
        RECT 252.700 39.125 256.255 39.145 ;
        POLYGON 252.635 39.125 252.635 39.110 252.580 39.110 ;
        RECT 252.635 39.110 256.255 39.125 ;
        RECT 242.470 39.100 246.470 39.110 ;
        POLYGON 246.470 39.110 246.505 39.100 246.470 39.100 ;
        POLYGON 252.580 39.110 252.580 39.100 252.545 39.100 ;
        RECT 252.580 39.100 256.255 39.110 ;
        RECT 242.470 39.095 246.505 39.100 ;
        RECT 233.475 38.945 238.320 39.095 ;
        POLYGON 233.475 38.945 233.485 38.945 233.485 38.930 ;
        RECT 233.485 38.930 238.320 38.945 ;
        RECT 210.730 38.585 225.835 38.930 ;
        POLYGON 210.730 38.585 211.000 38.585 211.000 38.020 ;
        RECT 211.000 38.335 225.835 38.585 ;
        POLYGON 225.835 38.930 226.200 38.335 225.835 38.335 ;
        POLYGON 233.485 38.930 233.620 38.930 233.620 38.770 ;
        RECT 233.620 38.825 238.320 38.930 ;
        POLYGON 238.320 39.095 238.605 38.825 238.320 38.825 ;
        POLYGON 242.470 39.095 242.885 39.095 242.885 38.840 ;
        RECT 242.885 39.090 246.505 39.095 ;
        POLYGON 246.505 39.100 246.545 39.090 246.505 39.090 ;
        POLYGON 252.545 39.100 252.545 39.090 252.505 39.090 ;
        RECT 252.545 39.090 256.255 39.100 ;
        RECT 242.885 39.045 246.545 39.090 ;
        POLYGON 246.545 39.090 246.710 39.045 246.545 39.045 ;
        POLYGON 252.505 39.090 252.505 39.075 252.450 39.075 ;
        RECT 252.505 39.075 256.255 39.090 ;
        POLYGON 252.450 39.075 252.450 39.070 252.435 39.070 ;
        RECT 252.450 39.070 256.255 39.075 ;
        POLYGON 252.430 39.070 252.430 39.050 252.350 39.050 ;
        RECT 252.430 39.065 256.255 39.070 ;
        POLYGON 256.255 39.375 256.720 39.375 256.255 39.065 ;
        POLYGON 260.045 39.375 260.045 39.065 259.735 39.065 ;
        RECT 260.045 39.260 263.820 39.375 ;
        POLYGON 263.820 39.495 263.975 39.495 263.820 39.265 ;
        POLYGON 269.085 39.495 269.085 39.265 268.980 39.265 ;
        RECT 269.085 39.265 276.895 39.495 ;
        RECT 260.045 39.065 263.495 39.260 ;
        RECT 252.430 39.050 255.775 39.065 ;
        POLYGON 252.350 39.050 252.350 39.045 252.325 39.045 ;
        RECT 252.350 39.045 255.775 39.050 ;
        RECT 242.885 39.035 246.710 39.045 ;
        POLYGON 246.710 39.045 246.775 39.035 246.710 39.035 ;
        POLYGON 252.325 39.045 252.325 39.035 252.290 39.035 ;
        RECT 252.325 39.035 255.775 39.045 ;
        RECT 242.885 39.030 246.775 39.035 ;
        POLYGON 246.775 39.035 246.805 39.030 246.775 39.030 ;
        POLYGON 252.290 39.035 252.290 39.030 252.270 39.030 ;
        RECT 252.290 39.030 255.775 39.035 ;
        RECT 242.885 39.025 246.805 39.030 ;
        POLYGON 246.805 39.030 246.820 39.025 246.805 39.025 ;
        POLYGON 252.270 39.030 252.270 39.025 252.250 39.025 ;
        RECT 252.270 39.025 255.775 39.030 ;
        RECT 242.885 38.995 246.820 39.025 ;
        POLYGON 246.820 39.025 246.960 38.995 246.820 38.995 ;
        POLYGON 252.250 39.025 252.250 39.010 252.195 39.010 ;
        RECT 252.250 39.010 255.775 39.025 ;
        POLYGON 252.195 39.010 252.195 39.005 252.155 39.005 ;
        RECT 252.195 39.005 255.775 39.010 ;
        POLYGON 252.155 39.005 252.155 38.995 252.100 38.995 ;
        RECT 252.155 38.995 255.775 39.005 ;
        RECT 242.885 38.990 246.960 38.995 ;
        POLYGON 246.960 38.995 247.005 38.990 246.960 38.990 ;
        POLYGON 252.100 38.995 252.100 38.990 252.080 38.990 ;
        RECT 252.100 38.990 255.775 38.995 ;
        RECT 242.885 38.975 247.010 38.990 ;
        POLYGON 247.010 38.990 247.085 38.975 247.010 38.975 ;
        POLYGON 252.080 38.990 252.080 38.980 252.040 38.980 ;
        RECT 252.080 38.980 255.775 38.990 ;
        POLYGON 252.040 38.980 252.040 38.975 252.015 38.975 ;
        RECT 252.040 38.975 255.775 38.980 ;
        RECT 242.885 38.970 247.085 38.975 ;
        POLYGON 247.085 38.975 247.125 38.970 247.085 38.970 ;
        POLYGON 252.015 38.975 252.015 38.970 251.990 38.970 ;
        RECT 252.015 38.970 255.775 38.975 ;
        RECT 242.885 38.955 247.130 38.970 ;
        POLYGON 247.130 38.970 247.215 38.955 247.130 38.955 ;
        POLYGON 251.990 38.970 251.990 38.960 251.940 38.960 ;
        RECT 251.990 38.960 255.775 38.970 ;
        POLYGON 251.940 38.960 251.940 38.955 251.905 38.955 ;
        RECT 251.940 38.955 255.775 38.960 ;
        RECT 242.885 38.935 247.215 38.955 ;
        POLYGON 247.215 38.955 247.335 38.935 247.215 38.935 ;
        POLYGON 251.905 38.955 251.905 38.950 251.865 38.950 ;
        RECT 251.905 38.950 255.775 38.955 ;
        POLYGON 251.855 38.950 251.855 38.935 251.765 38.935 ;
        RECT 251.855 38.935 255.775 38.950 ;
        RECT 242.885 38.920 247.340 38.935 ;
        POLYGON 247.340 38.935 247.480 38.920 247.340 38.920 ;
        POLYGON 251.765 38.935 251.765 38.920 251.670 38.920 ;
        RECT 251.765 38.920 255.775 38.935 ;
        RECT 242.885 38.910 247.485 38.920 ;
        POLYGON 247.485 38.920 247.585 38.910 247.485 38.910 ;
        POLYGON 251.670 38.920 251.670 38.915 251.615 38.915 ;
        RECT 251.670 38.915 255.775 38.920 ;
        POLYGON 251.615 38.915 251.615 38.910 251.575 38.910 ;
        RECT 251.615 38.910 255.775 38.915 ;
        RECT 242.885 38.895 247.590 38.910 ;
        POLYGON 247.590 38.910 247.735 38.895 247.590 38.895 ;
        POLYGON 251.575 38.910 251.575 38.905 251.530 38.905 ;
        RECT 251.575 38.905 255.775 38.910 ;
        POLYGON 251.530 38.905 251.530 38.895 251.430 38.895 ;
        RECT 251.530 38.895 255.775 38.905 ;
        RECT 242.885 38.890 247.740 38.895 ;
        POLYGON 247.740 38.895 247.765 38.890 247.740 38.890 ;
        POLYGON 251.430 38.895 251.430 38.890 251.380 38.890 ;
        RECT 251.430 38.890 255.775 38.895 ;
        RECT 242.885 38.885 247.765 38.890 ;
        POLYGON 247.765 38.890 247.835 38.885 247.765 38.885 ;
        POLYGON 251.340 38.890 251.340 38.885 251.285 38.885 ;
        RECT 251.340 38.885 255.775 38.890 ;
        RECT 242.885 38.875 247.840 38.885 ;
        POLYGON 247.840 38.885 248.000 38.875 247.840 38.875 ;
        POLYGON 251.285 38.885 251.285 38.875 251.180 38.875 ;
        RECT 251.285 38.875 255.775 38.885 ;
        RECT 242.885 38.870 248.010 38.875 ;
        POLYGON 248.010 38.875 248.065 38.870 248.010 38.870 ;
        POLYGON 251.175 38.875 251.175 38.870 251.075 38.870 ;
        RECT 251.175 38.870 255.775 38.875 ;
        RECT 242.885 38.860 248.100 38.870 ;
        POLYGON 248.100 38.870 248.285 38.860 248.100 38.860 ;
        POLYGON 251.065 38.870 251.065 38.860 250.815 38.860 ;
        RECT 251.065 38.860 255.775 38.870 ;
        RECT 242.885 38.850 248.370 38.860 ;
        POLYGON 248.370 38.860 248.635 38.850 248.370 38.850 ;
        POLYGON 250.815 38.860 250.815 38.850 250.560 38.850 ;
        RECT 250.815 38.850 255.775 38.860 ;
        RECT 242.885 38.845 248.660 38.850 ;
        POLYGON 248.660 38.850 248.745 38.845 248.660 38.845 ;
        POLYGON 250.560 38.850 250.560 38.845 250.435 38.845 ;
        RECT 250.560 38.845 255.775 38.850 ;
        RECT 242.885 38.840 248.940 38.845 ;
        POLYGON 248.940 38.845 248.945 38.840 248.940 38.840 ;
        POLYGON 250.365 38.845 250.365 38.840 250.015 38.840 ;
        RECT 250.365 38.840 255.775 38.845 ;
        POLYGON 242.885 38.840 242.910 38.840 242.910 38.825 ;
        RECT 242.910 38.835 249.355 38.840 ;
        POLYGON 249.355 38.840 249.540 38.835 249.355 38.835 ;
        POLYGON 250.015 38.840 250.015 38.835 249.665 38.835 ;
        RECT 250.015 38.835 255.775 38.840 ;
        RECT 242.910 38.825 255.775 38.835 ;
        RECT 233.620 38.795 238.605 38.825 ;
        POLYGON 238.605 38.825 238.640 38.795 238.605 38.795 ;
        POLYGON 242.910 38.825 242.970 38.825 242.970 38.795 ;
        RECT 242.970 38.795 255.775 38.825 ;
        RECT 233.620 38.770 238.640 38.795 ;
        POLYGON 233.620 38.770 233.880 38.770 233.880 38.465 ;
        RECT 233.880 38.725 238.640 38.770 ;
        POLYGON 238.640 38.795 238.710 38.725 238.640 38.725 ;
        POLYGON 242.970 38.795 243.100 38.795 243.100 38.725 ;
        RECT 243.100 38.775 255.775 38.795 ;
        POLYGON 255.775 39.065 256.255 39.065 255.775 38.775 ;
        POLYGON 259.735 39.065 259.735 38.985 259.655 38.985 ;
        RECT 259.735 38.985 263.495 39.065 ;
        POLYGON 259.655 38.985 259.655 38.820 259.495 38.820 ;
        RECT 259.655 38.825 263.495 38.985 ;
        POLYGON 263.495 39.260 263.820 39.260 263.495 38.825 ;
        POLYGON 268.980 39.265 268.980 39.105 268.910 39.105 ;
        RECT 268.980 39.105 276.895 39.265 ;
        POLYGON 268.910 39.105 268.910 38.965 268.845 38.965 ;
        RECT 268.910 38.965 276.895 39.105 ;
        POLYGON 268.845 38.965 268.845 38.830 268.780 38.830 ;
        RECT 268.845 38.905 276.895 38.965 ;
        POLYGON 276.895 39.495 277.040 39.495 276.895 38.905 ;
        POLYGON 287.545 39.495 287.545 38.925 287.515 38.925 ;
        RECT 287.545 38.925 303.120 39.540 ;
        RECT 268.845 38.830 276.535 38.905 ;
        RECT 259.655 38.820 263.240 38.825 ;
        POLYGON 259.495 38.820 259.495 38.775 259.450 38.775 ;
        RECT 259.495 38.775 263.240 38.820 ;
        RECT 243.100 38.740 255.720 38.775 ;
        POLYGON 255.720 38.775 255.775 38.775 255.720 38.740 ;
        POLYGON 259.450 38.775 259.450 38.740 259.415 38.740 ;
        RECT 259.450 38.740 263.240 38.775 ;
        RECT 243.100 38.725 255.295 38.740 ;
        RECT 233.880 38.510 238.710 38.725 ;
        POLYGON 238.710 38.725 238.965 38.510 238.710 38.510 ;
        POLYGON 243.100 38.725 243.190 38.725 243.190 38.680 ;
        RECT 243.190 38.680 255.295 38.725 ;
        POLYGON 243.190 38.680 243.455 38.680 243.455 38.540 ;
        RECT 243.455 38.540 255.295 38.680 ;
        POLYGON 243.455 38.540 243.505 38.540 243.505 38.510 ;
        RECT 243.505 38.510 255.295 38.540 ;
        RECT 233.880 38.465 238.965 38.510 ;
        POLYGON 233.880 38.465 233.990 38.465 233.990 38.335 ;
        RECT 233.990 38.375 238.965 38.465 ;
        POLYGON 238.965 38.510 239.125 38.375 238.965 38.375 ;
        POLYGON 243.505 38.510 243.645 38.510 243.645 38.435 ;
        RECT 243.645 38.505 255.295 38.510 ;
        POLYGON 255.295 38.740 255.720 38.740 255.295 38.505 ;
        POLYGON 259.415 38.740 259.415 38.605 259.280 38.605 ;
        RECT 259.415 38.605 263.240 38.740 ;
        POLYGON 259.280 38.605 259.280 38.545 259.210 38.545 ;
        RECT 259.280 38.545 263.240 38.605 ;
        POLYGON 259.210 38.545 259.210 38.505 259.165 38.505 ;
        RECT 259.210 38.505 263.240 38.545 ;
        POLYGON 263.240 38.825 263.495 38.825 263.240 38.505 ;
        POLYGON 268.780 38.825 268.780 38.725 268.730 38.725 ;
        RECT 268.780 38.725 276.535 38.830 ;
        POLYGON 268.730 38.725 268.730 38.680 268.705 38.680 ;
        RECT 268.730 38.680 276.535 38.725 ;
        POLYGON 268.705 38.680 268.705 38.505 268.620 38.505 ;
        RECT 268.705 38.505 276.535 38.680 ;
        RECT 243.645 38.500 255.280 38.505 ;
        POLYGON 255.280 38.505 255.295 38.505 255.280 38.500 ;
        POLYGON 259.165 38.505 259.165 38.500 259.160 38.500 ;
        RECT 259.165 38.500 263.145 38.505 ;
        RECT 243.645 38.435 254.885 38.500 ;
        POLYGON 243.645 38.435 243.770 38.435 243.770 38.375 ;
        RECT 243.770 38.375 254.885 38.435 ;
        RECT 233.990 38.370 239.125 38.375 ;
        POLYGON 239.125 38.375 239.130 38.370 239.125 38.370 ;
        POLYGON 243.770 38.375 243.780 38.375 243.780 38.370 ;
        RECT 243.780 38.370 254.885 38.375 ;
        RECT 233.990 38.335 239.130 38.370 ;
        RECT 211.000 38.170 226.200 38.335 ;
        POLYGON 226.200 38.335 226.300 38.170 226.200 38.170 ;
        POLYGON 233.990 38.335 234.010 38.335 234.010 38.315 ;
        RECT 234.010 38.315 239.130 38.335 ;
        POLYGON 234.010 38.315 234.140 38.315 234.140 38.170 ;
        RECT 234.140 38.200 239.130 38.315 ;
        POLYGON 239.130 38.370 239.330 38.200 239.130 38.200 ;
        POLYGON 243.780 38.370 243.960 38.370 243.960 38.285 ;
        RECT 243.960 38.300 254.885 38.370 ;
        POLYGON 254.885 38.500 255.280 38.500 254.885 38.300 ;
        POLYGON 259.160 38.500 259.160 38.490 259.150 38.490 ;
        RECT 259.160 38.490 263.145 38.500 ;
        POLYGON 259.150 38.490 259.150 38.300 258.940 38.300 ;
        RECT 259.150 38.385 263.145 38.490 ;
        POLYGON 263.145 38.505 263.240 38.505 263.145 38.385 ;
        POLYGON 268.620 38.505 268.620 38.390 268.565 38.390 ;
        RECT 268.620 38.390 276.535 38.505 ;
        RECT 259.150 38.300 262.770 38.385 ;
        RECT 243.960 38.285 254.770 38.300 ;
        POLYGON 243.960 38.285 244.130 38.285 244.130 38.200 ;
        RECT 244.130 38.245 254.770 38.285 ;
        POLYGON 254.770 38.300 254.885 38.300 254.770 38.245 ;
        POLYGON 258.940 38.300 258.940 38.270 258.905 38.270 ;
        RECT 258.940 38.270 262.770 38.300 ;
        POLYGON 258.905 38.270 258.905 38.245 258.880 38.245 ;
        RECT 258.905 38.245 262.770 38.270 ;
        RECT 244.130 38.200 254.225 38.245 ;
        RECT 234.140 38.170 239.330 38.200 ;
        RECT 211.000 38.075 226.300 38.170 ;
        POLYGON 226.300 38.170 226.360 38.075 226.300 38.075 ;
        POLYGON 234.140 38.170 234.225 38.170 234.225 38.075 ;
        RECT 234.225 38.075 239.330 38.170 ;
        RECT 211.000 38.020 226.360 38.075 ;
        POLYGON 211.000 38.020 211.420 38.020 211.420 37.220 ;
        RECT 211.420 37.510 226.360 38.020 ;
        POLYGON 226.360 38.075 226.730 37.510 226.360 37.510 ;
        POLYGON 234.225 38.075 234.380 38.075 234.380 37.910 ;
        RECT 234.380 37.980 239.330 38.075 ;
        POLYGON 239.330 38.200 239.615 37.980 239.330 37.980 ;
        POLYGON 244.130 38.200 244.440 38.200 244.440 38.050 ;
        RECT 244.440 38.050 254.225 38.200 ;
        POLYGON 244.440 38.050 244.525 38.050 244.525 38.010 ;
        RECT 244.525 38.010 254.225 38.050 ;
        POLYGON 244.530 38.010 244.595 38.010 244.595 37.980 ;
        RECT 244.595 37.995 254.225 38.010 ;
        POLYGON 254.225 38.245 254.770 38.245 254.225 37.995 ;
        POLYGON 258.880 38.245 258.880 38.160 258.790 38.160 ;
        RECT 258.880 38.160 262.770 38.245 ;
        POLYGON 258.790 38.160 258.790 38.125 258.750 38.125 ;
        RECT 258.790 38.125 262.770 38.160 ;
        POLYGON 258.750 38.125 258.750 37.995 258.605 37.995 ;
        RECT 258.750 37.995 262.770 38.125 ;
        RECT 244.595 37.980 254.090 37.995 ;
        RECT 234.380 37.950 239.615 37.980 ;
        POLYGON 239.615 37.980 239.655 37.950 239.615 37.950 ;
        POLYGON 244.595 37.980 244.660 37.980 244.660 37.950 ;
        RECT 244.660 37.950 254.090 37.980 ;
        RECT 234.380 37.925 239.655 37.950 ;
        POLYGON 239.655 37.950 239.690 37.925 239.655 37.925 ;
        POLYGON 244.660 37.950 244.715 37.950 244.715 37.925 ;
        RECT 244.715 37.930 254.090 37.950 ;
        POLYGON 254.090 37.995 254.225 37.995 254.090 37.930 ;
        POLYGON 258.605 37.995 258.605 37.930 258.530 37.930 ;
        RECT 258.605 37.940 262.770 37.995 ;
        POLYGON 262.770 38.385 263.145 38.385 262.770 37.945 ;
        POLYGON 268.565 38.385 268.565 38.015 268.385 38.015 ;
        RECT 268.565 38.015 276.535 38.390 ;
        POLYGON 268.385 38.015 268.385 37.950 268.350 37.950 ;
        RECT 268.385 37.950 276.535 38.015 ;
        RECT 258.605 37.930 262.115 37.940 ;
        RECT 244.715 37.925 254.045 37.930 ;
        RECT 234.380 37.910 239.690 37.925 ;
        POLYGON 234.380 37.910 234.570 37.910 234.570 37.695 ;
        RECT 234.570 37.705 239.690 37.910 ;
        POLYGON 239.690 37.925 239.975 37.705 239.690 37.705 ;
        POLYGON 244.715 37.925 244.750 37.925 244.750 37.910 ;
        RECT 244.750 37.910 254.045 37.925 ;
        POLYGON 254.045 37.930 254.090 37.930 254.045 37.910 ;
        POLYGON 258.530 37.930 258.530 37.910 258.505 37.910 ;
        RECT 258.530 37.910 262.115 37.930 ;
        POLYGON 244.750 37.910 245.095 37.910 245.095 37.755 ;
        RECT 245.095 37.755 253.505 37.910 ;
        POLYGON 245.095 37.755 245.220 37.755 245.220 37.705 ;
        RECT 245.220 37.705 253.505 37.755 ;
        RECT 234.570 37.695 239.975 37.705 ;
        POLYGON 234.570 37.695 234.750 37.695 234.750 37.510 ;
        RECT 234.750 37.530 239.975 37.695 ;
        POLYGON 239.975 37.705 240.225 37.530 239.975 37.530 ;
        POLYGON 245.220 37.705 245.385 37.705 245.385 37.640 ;
        RECT 245.385 37.690 253.505 37.705 ;
        POLYGON 253.505 37.910 254.045 37.910 253.505 37.690 ;
        POLYGON 258.505 37.910 258.505 37.900 258.495 37.900 ;
        RECT 258.505 37.900 262.115 37.910 ;
        POLYGON 258.495 37.900 258.495 37.825 258.410 37.825 ;
        RECT 258.495 37.825 262.115 37.900 ;
        POLYGON 258.410 37.825 258.410 37.730 258.295 37.730 ;
        RECT 258.410 37.730 262.115 37.825 ;
        POLYGON 258.295 37.730 258.295 37.690 258.245 37.690 ;
        RECT 258.295 37.690 262.115 37.730 ;
        RECT 245.385 37.640 253.235 37.690 ;
        POLYGON 245.385 37.640 245.555 37.640 245.555 37.580 ;
        RECT 245.555 37.590 253.235 37.640 ;
        POLYGON 253.235 37.690 253.505 37.690 253.235 37.590 ;
        POLYGON 258.245 37.690 258.245 37.600 258.135 37.600 ;
        RECT 258.245 37.600 262.115 37.690 ;
        POLYGON 258.135 37.600 258.135 37.590 258.125 37.590 ;
        RECT 258.135 37.590 262.115 37.600 ;
        RECT 245.555 37.580 253.195 37.590 ;
        POLYGON 245.560 37.580 245.600 37.580 245.600 37.560 ;
        RECT 245.600 37.575 253.195 37.580 ;
        POLYGON 253.195 37.590 253.235 37.590 253.195 37.575 ;
        POLYGON 258.125 37.590 258.125 37.575 258.110 37.575 ;
        RECT 258.125 37.575 262.115 37.590 ;
        RECT 245.600 37.565 253.155 37.575 ;
        POLYGON 253.155 37.575 253.195 37.575 253.155 37.565 ;
        POLYGON 258.110 37.575 258.110 37.565 258.095 37.565 ;
        RECT 258.110 37.565 262.115 37.575 ;
        RECT 245.600 37.560 252.970 37.565 ;
        POLYGON 245.605 37.560 245.695 37.560 245.695 37.530 ;
        RECT 245.695 37.530 252.970 37.560 ;
        RECT 234.750 37.510 240.225 37.530 ;
        POLYGON 240.225 37.530 240.255 37.510 240.225 37.510 ;
        POLYGON 245.695 37.530 245.760 37.530 245.760 37.510 ;
        RECT 245.760 37.510 252.970 37.530 ;
        RECT 211.420 37.430 226.730 37.510 ;
        POLYGON 226.730 37.510 226.785 37.430 226.730 37.430 ;
        POLYGON 234.750 37.510 234.830 37.510 234.830 37.430 ;
        RECT 234.830 37.455 240.255 37.510 ;
        POLYGON 240.255 37.510 240.335 37.455 240.255 37.455 ;
        POLYGON 245.760 37.510 245.940 37.510 245.940 37.455 ;
        RECT 245.940 37.505 252.970 37.510 ;
        POLYGON 252.970 37.565 253.155 37.565 252.970 37.505 ;
        POLYGON 258.095 37.565 258.095 37.505 258.015 37.505 ;
        RECT 258.095 37.505 262.115 37.565 ;
        RECT 245.940 37.455 252.705 37.505 ;
        RECT 234.830 37.430 240.335 37.455 ;
        RECT 211.420 37.215 226.785 37.430 ;
        RECT 181.540 37.105 197.580 37.215 ;
        RECT 167.110 37.040 172.665 37.105 ;
        POLYGON 167.030 37.040 167.030 36.905 166.895 36.905 ;
        RECT 167.030 36.905 172.665 37.040 ;
        RECT 117.690 36.865 162.055 36.905 ;
        POLYGON 162.055 36.905 162.120 36.905 162.055 36.865 ;
        POLYGON 166.895 36.905 166.895 36.865 166.855 36.865 ;
        RECT 166.895 36.865 172.665 36.905 ;
        RECT 117.690 36.785 161.805 36.865 ;
        RECT 59.505 36.635 116.600 36.785 ;
        POLYGON 59.505 36.635 60.145 36.635 60.145 35.585 ;
        RECT 60.145 35.585 116.600 36.635 ;
        POLYGON 116.600 36.785 117.280 35.585 116.600 35.585 ;
        POLYGON 117.690 36.785 117.695 36.785 117.695 36.725 ;
        RECT 117.695 36.720 161.805 36.785 ;
        POLYGON 161.805 36.865 162.055 36.865 161.805 36.720 ;
        POLYGON 166.855 36.865 166.855 36.720 166.710 36.720 ;
        RECT 166.855 36.725 172.665 36.865 ;
        POLYGON 172.665 37.105 172.905 37.105 172.665 36.725 ;
        POLYGON 181.360 37.105 181.360 36.730 181.230 36.730 ;
        RECT 181.360 36.730 197.580 37.105 ;
        RECT 166.855 36.720 172.615 36.725 ;
        RECT 117.695 36.690 161.485 36.720 ;
        POLYGON 117.695 36.690 117.745 36.690 117.745 36.020 ;
        RECT 117.745 36.530 161.485 36.690 ;
        POLYGON 161.485 36.720 161.805 36.720 161.485 36.530 ;
        POLYGON 166.710 36.720 166.710 36.605 166.595 36.605 ;
        RECT 166.710 36.645 172.615 36.720 ;
        POLYGON 172.615 36.725 172.665 36.725 172.615 36.645 ;
        POLYGON 181.230 36.725 181.230 36.645 181.200 36.645 ;
        RECT 181.230 36.645 197.580 36.730 ;
        RECT 166.710 36.605 172.270 36.645 ;
        POLYGON 166.595 36.605 166.595 36.570 166.555 36.570 ;
        RECT 166.595 36.570 172.270 36.605 ;
        POLYGON 166.555 36.570 166.555 36.530 166.515 36.530 ;
        RECT 166.555 36.530 172.270 36.570 ;
        RECT 117.745 36.370 161.175 36.530 ;
        POLYGON 161.175 36.530 161.485 36.530 161.175 36.370 ;
        POLYGON 166.515 36.530 166.515 36.370 166.345 36.370 ;
        RECT 166.515 36.370 172.270 36.530 ;
        RECT 117.745 36.260 160.970 36.370 ;
        POLYGON 160.970 36.370 161.175 36.370 160.970 36.260 ;
        POLYGON 166.345 36.370 166.345 36.260 166.225 36.260 ;
        RECT 166.345 36.260 172.270 36.370 ;
        RECT 117.745 36.190 160.830 36.260 ;
        POLYGON 160.830 36.260 160.970 36.260 160.830 36.190 ;
        POLYGON 166.225 36.260 166.225 36.225 166.190 36.225 ;
        RECT 166.225 36.225 172.270 36.260 ;
        POLYGON 166.190 36.225 166.190 36.190 166.150 36.190 ;
        RECT 166.190 36.190 172.270 36.225 ;
        RECT 117.745 36.050 160.520 36.190 ;
        POLYGON 160.520 36.190 160.830 36.190 160.520 36.050 ;
        POLYGON 166.150 36.190 166.150 36.115 166.070 36.115 ;
        RECT 166.150 36.150 172.270 36.190 ;
        POLYGON 172.270 36.645 172.615 36.645 172.270 36.150 ;
        POLYGON 181.200 36.640 181.200 36.420 181.125 36.420 ;
        RECT 181.200 36.420 197.580 36.645 ;
        POLYGON 181.125 36.420 181.125 36.155 181.020 36.155 ;
        RECT 181.125 36.155 197.580 36.420 ;
        RECT 166.150 36.115 171.875 36.150 ;
        POLYGON 166.070 36.115 166.070 36.100 166.050 36.100 ;
        RECT 166.070 36.100 171.875 36.115 ;
        POLYGON 166.050 36.100 166.050 36.050 165.995 36.050 ;
        RECT 166.050 36.050 171.875 36.100 ;
        RECT 117.745 35.985 160.160 36.050 ;
        POLYGON 117.745 35.985 117.750 35.985 117.750 35.950 ;
        RECT 117.750 35.905 160.160 35.985 ;
        POLYGON 117.750 35.905 117.775 35.905 117.775 35.600 ;
        RECT 117.775 35.885 160.160 35.905 ;
        POLYGON 160.160 36.050 160.520 36.050 160.160 35.885 ;
        POLYGON 165.995 36.050 165.995 35.920 165.845 35.920 ;
        RECT 165.995 35.920 171.875 36.050 ;
        POLYGON 165.845 35.920 165.845 35.885 165.805 35.885 ;
        RECT 165.845 35.885 171.875 35.920 ;
        RECT 117.775 35.775 159.865 35.885 ;
        POLYGON 159.865 35.885 160.160 35.885 159.865 35.775 ;
        POLYGON 165.805 35.885 165.805 35.775 165.675 35.775 ;
        RECT 165.805 35.775 171.875 35.885 ;
        RECT 117.775 35.765 159.845 35.775 ;
        POLYGON 159.845 35.775 159.865 35.775 159.845 35.765 ;
        POLYGON 165.675 35.775 165.675 35.765 165.665 35.765 ;
        RECT 165.675 35.765 171.875 35.775 ;
        RECT 117.775 35.625 159.470 35.765 ;
        POLYGON 159.470 35.765 159.845 35.765 159.470 35.625 ;
        POLYGON 165.665 35.765 165.665 35.690 165.575 35.690 ;
        RECT 165.665 35.690 171.875 35.765 ;
        POLYGON 165.575 35.690 165.575 35.675 165.560 35.675 ;
        RECT 165.575 35.675 171.875 35.690 ;
        POLYGON 165.560 35.675 165.560 35.625 165.495 35.625 ;
        RECT 165.560 35.630 171.875 35.675 ;
        POLYGON 171.875 36.150 172.270 36.150 171.875 35.630 ;
        POLYGON 181.020 36.150 181.020 35.915 180.925 35.915 ;
        RECT 181.020 35.915 197.580 36.155 ;
        POLYGON 180.925 35.915 180.925 35.630 180.810 35.630 ;
        RECT 180.925 35.630 197.580 35.915 ;
        RECT 165.560 35.625 171.435 35.630 ;
        RECT 117.775 35.585 159.145 35.625 ;
        RECT 14.030 34.580 22.645 35.585 ;
        POLYGON 14.030 34.580 14.625 34.580 14.625 29.755 ;
        RECT 14.625 29.755 22.645 34.580 ;
        POLYGON 14.625 29.755 16.145 29.755 16.145 21.130 ;
        RECT 16.145 29.560 22.645 29.755 ;
        POLYGON 22.645 35.585 23.480 29.560 22.645 29.560 ;
        POLYGON 60.145 35.585 60.990 35.585 60.990 34.200 ;
        RECT 60.990 35.180 117.280 35.585 ;
        POLYGON 117.280 35.585 117.530 35.180 117.280 35.180 ;
        POLYGON 117.775 35.585 117.780 35.585 117.780 35.560 ;
        RECT 117.780 35.535 159.145 35.585 ;
        POLYGON 117.780 35.535 117.815 35.535 117.815 35.310 ;
        RECT 117.815 35.520 159.145 35.535 ;
        POLYGON 159.145 35.625 159.470 35.625 159.145 35.520 ;
        POLYGON 165.495 35.625 165.495 35.610 165.475 35.610 ;
        RECT 165.495 35.610 171.435 35.625 ;
        POLYGON 165.475 35.610 165.475 35.520 165.365 35.520 ;
        RECT 165.475 35.520 171.435 35.610 ;
        RECT 117.815 35.395 158.755 35.520 ;
        POLYGON 158.755 35.520 159.145 35.520 158.755 35.395 ;
        POLYGON 165.365 35.520 165.365 35.395 165.210 35.395 ;
        RECT 165.365 35.395 171.435 35.520 ;
        RECT 117.815 35.390 158.740 35.395 ;
        POLYGON 158.740 35.395 158.755 35.395 158.740 35.390 ;
        POLYGON 165.210 35.395 165.210 35.390 165.200 35.390 ;
        RECT 165.210 35.390 171.435 35.395 ;
        RECT 117.815 35.310 158.435 35.390 ;
        POLYGON 158.435 35.390 158.740 35.390 158.435 35.310 ;
        POLYGON 165.200 35.390 165.200 35.320 165.115 35.320 ;
        RECT 165.200 35.320 171.435 35.390 ;
        POLYGON 165.115 35.320 165.115 35.310 165.105 35.310 ;
        RECT 165.115 35.310 171.435 35.320 ;
        RECT 117.815 35.300 158.025 35.310 ;
        POLYGON 117.815 35.300 117.830 35.300 117.830 35.200 ;
        RECT 117.830 35.205 158.025 35.300 ;
        POLYGON 158.025 35.310 158.430 35.310 158.025 35.205 ;
        POLYGON 165.105 35.310 165.105 35.300 165.090 35.300 ;
        RECT 165.105 35.300 171.435 35.310 ;
        POLYGON 165.090 35.300 165.090 35.260 165.045 35.260 ;
        RECT 165.090 35.260 171.435 35.300 ;
        POLYGON 165.040 35.260 165.040 35.205 164.965 35.205 ;
        RECT 165.040 35.205 171.435 35.260 ;
        RECT 117.830 35.180 157.710 35.205 ;
        RECT 60.990 34.780 117.530 35.180 ;
        POLYGON 117.530 35.180 117.775 34.780 117.530 34.780 ;
        POLYGON 117.830 35.180 117.835 35.180 117.835 35.165 ;
        RECT 117.835 35.140 157.710 35.180 ;
        POLYGON 157.710 35.205 158.025 35.205 157.710 35.140 ;
        POLYGON 164.965 35.205 164.965 35.140 164.880 35.140 ;
        RECT 164.965 35.140 171.435 35.205 ;
        RECT 117.835 35.135 157.600 35.140 ;
        POLYGON 117.835 35.135 117.885 35.135 117.885 34.805 ;
        RECT 117.885 35.115 157.600 35.135 ;
        POLYGON 157.600 35.140 157.710 35.140 157.600 35.115 ;
        POLYGON 164.880 35.140 164.880 35.115 164.845 35.115 ;
        RECT 164.880 35.115 171.435 35.140 ;
        RECT 117.885 35.045 157.270 35.115 ;
        POLYGON 157.270 35.115 157.600 35.115 157.270 35.045 ;
        POLYGON 164.845 35.115 164.845 35.045 164.750 35.045 ;
        RECT 164.845 35.090 171.435 35.115 ;
        POLYGON 171.435 35.630 171.875 35.630 171.435 35.090 ;
        POLYGON 180.810 35.630 180.810 35.320 180.685 35.320 ;
        RECT 180.810 35.485 197.580 35.630 ;
        POLYGON 197.580 37.215 197.810 37.215 197.580 35.485 ;
        POLYGON 211.420 37.215 211.430 37.215 211.430 37.205 ;
        RECT 211.430 37.210 226.785 37.215 ;
        POLYGON 226.785 37.430 226.940 37.210 226.785 37.210 ;
        RECT 211.430 37.205 226.940 37.210 ;
        POLYGON 234.830 37.430 235.050 37.430 235.050 37.205 ;
        RECT 235.050 37.240 240.335 37.430 ;
        POLYGON 240.335 37.455 240.645 37.240 240.335 37.240 ;
        POLYGON 245.940 37.455 246.220 37.455 246.220 37.390 ;
        RECT 246.220 37.435 252.705 37.455 ;
        POLYGON 252.705 37.505 252.970 37.505 252.705 37.435 ;
        POLYGON 258.015 37.505 258.015 37.500 258.010 37.500 ;
        RECT 258.015 37.500 262.115 37.505 ;
        POLYGON 258.010 37.500 258.010 37.435 257.925 37.435 ;
        RECT 258.010 37.435 262.115 37.500 ;
        RECT 246.220 37.390 252.435 37.435 ;
        POLYGON 246.220 37.390 246.375 37.390 246.375 37.360 ;
        RECT 246.375 37.380 252.435 37.390 ;
        POLYGON 252.435 37.435 252.705 37.435 252.435 37.380 ;
        POLYGON 257.925 37.435 257.925 37.380 257.855 37.380 ;
        RECT 257.925 37.380 262.115 37.435 ;
        RECT 246.375 37.365 252.340 37.380 ;
        POLYGON 252.340 37.380 252.435 37.380 252.340 37.365 ;
        POLYGON 257.855 37.380 257.855 37.375 257.850 37.375 ;
        RECT 257.855 37.375 262.115 37.380 ;
        POLYGON 257.850 37.375 257.850 37.365 257.835 37.365 ;
        RECT 257.850 37.365 262.115 37.375 ;
        RECT 246.375 37.360 252.155 37.365 ;
        POLYGON 246.380 37.360 246.505 37.360 246.505 37.340 ;
        RECT 246.505 37.340 252.155 37.360 ;
        POLYGON 246.505 37.340 246.680 37.340 246.680 37.315 ;
        RECT 246.680 37.330 252.155 37.340 ;
        POLYGON 252.155 37.365 252.340 37.365 252.155 37.330 ;
        POLYGON 257.835 37.365 257.835 37.330 257.790 37.330 ;
        RECT 257.835 37.330 262.115 37.365 ;
        RECT 246.680 37.325 252.080 37.330 ;
        POLYGON 252.080 37.330 252.155 37.330 252.080 37.325 ;
        POLYGON 257.790 37.330 257.790 37.325 257.780 37.325 ;
        RECT 257.790 37.325 262.115 37.330 ;
        RECT 246.680 37.315 251.855 37.325 ;
        POLYGON 246.685 37.315 246.805 37.315 246.805 37.295 ;
        RECT 246.805 37.295 251.855 37.315 ;
        POLYGON 251.855 37.325 252.080 37.325 251.855 37.295 ;
        POLYGON 257.780 37.325 257.780 37.295 257.740 37.295 ;
        RECT 257.780 37.295 262.115 37.325 ;
        POLYGON 246.805 37.295 247.130 37.295 247.130 37.265 ;
        RECT 247.130 37.265 251.530 37.295 ;
        POLYGON 251.530 37.295 251.855 37.295 251.530 37.265 ;
        POLYGON 257.740 37.295 257.740 37.265 257.700 37.265 ;
        RECT 257.740 37.265 262.115 37.295 ;
        POLYGON 247.130 37.265 247.195 37.265 247.195 37.260 ;
        RECT 247.195 37.260 251.180 37.265 ;
        POLYGON 247.210 37.260 247.485 37.260 247.485 37.245 ;
        RECT 247.485 37.245 251.180 37.260 ;
        POLYGON 251.180 37.265 251.480 37.265 251.180 37.245 ;
        POLYGON 257.700 37.265 257.700 37.245 257.670 37.245 ;
        RECT 257.700 37.245 262.115 37.265 ;
        POLYGON 247.485 37.245 247.750 37.245 247.750 37.240 ;
        RECT 247.750 37.240 251.000 37.245 ;
        POLYGON 251.000 37.245 251.180 37.245 251.000 37.240 ;
        POLYGON 257.670 37.245 257.670 37.240 257.665 37.240 ;
        RECT 257.670 37.240 262.115 37.245 ;
        RECT 235.050 37.205 240.645 37.240 ;
        POLYGON 240.645 37.240 240.700 37.205 240.645 37.205 ;
        POLYGON 247.760 37.240 248.050 37.240 248.050 37.230 ;
        RECT 248.050 37.230 250.625 37.240 ;
        POLYGON 250.625 37.240 250.995 37.240 250.625 37.230 ;
        POLYGON 257.665 37.240 257.665 37.230 257.650 37.230 ;
        RECT 257.665 37.235 262.115 37.240 ;
        POLYGON 262.115 37.940 262.770 37.940 262.115 37.235 ;
        POLYGON 268.350 37.945 268.350 37.800 268.270 37.800 ;
        RECT 268.350 37.800 276.535 37.950 ;
        POLYGON 268.270 37.800 268.270 37.240 267.965 37.240 ;
        RECT 268.270 37.655 276.535 37.800 ;
        POLYGON 276.535 38.905 276.895 38.905 276.535 37.655 ;
        POLYGON 287.515 38.905 287.515 37.690 287.450 37.690 ;
        RECT 287.515 37.690 303.120 38.925 ;
        RECT 268.270 37.240 276.380 37.655 ;
        RECT 257.665 37.230 262.085 37.235 ;
        POLYGON 248.055 37.230 248.315 37.230 248.315 37.225 ;
        RECT 248.315 37.225 250.365 37.230 ;
        POLYGON 250.365 37.230 250.620 37.230 250.365 37.225 ;
        POLYGON 257.650 37.230 257.650 37.225 257.645 37.225 ;
        RECT 257.650 37.225 262.085 37.230 ;
        POLYGON 248.315 37.225 248.730 37.225 248.730 37.220 ;
        RECT 248.730 37.220 249.920 37.225 ;
        POLYGON 249.920 37.225 250.365 37.225 249.920 37.220 ;
        POLYGON 257.645 37.225 257.645 37.220 257.635 37.220 ;
        RECT 257.645 37.220 262.085 37.225 ;
        POLYGON 257.635 37.220 257.635 37.205 257.615 37.205 ;
        RECT 257.635 37.205 262.085 37.220 ;
        POLYGON 262.085 37.235 262.115 37.235 262.085 37.205 ;
        POLYGON 267.965 37.235 267.965 37.205 267.945 37.205 ;
        RECT 267.965 37.205 276.380 37.240 ;
        POLYGON 276.380 37.655 276.535 37.655 276.380 37.205 ;
        POLYGON 287.450 37.655 287.450 37.215 287.425 37.215 ;
        RECT 287.450 37.215 303.120 37.690 ;
        POLYGON 211.430 37.205 211.475 37.205 211.475 37.120 ;
        RECT 211.475 37.120 226.940 37.205 ;
        POLYGON 211.475 37.120 211.645 37.120 211.645 36.800 ;
        RECT 211.645 37.020 226.940 37.120 ;
        POLYGON 226.940 37.205 227.075 37.020 226.940 37.020 ;
        POLYGON 235.050 37.205 235.235 37.205 235.235 37.020 ;
        RECT 235.235 37.125 240.700 37.205 ;
        POLYGON 240.700 37.205 240.830 37.125 240.700 37.125 ;
        POLYGON 257.615 37.205 257.615 37.190 257.595 37.190 ;
        RECT 257.615 37.190 261.950 37.205 ;
        POLYGON 257.595 37.190 257.595 37.125 257.500 37.125 ;
        RECT 257.595 37.125 261.950 37.190 ;
        RECT 235.235 37.020 240.830 37.125 ;
        RECT 211.645 36.800 227.075 37.020 ;
        POLYGON 211.645 36.800 212.275 36.800 212.275 35.690 ;
        RECT 212.275 36.710 227.075 36.800 ;
        POLYGON 227.075 37.020 227.295 36.710 227.075 36.710 ;
        POLYGON 235.235 37.020 235.275 37.020 235.275 36.985 ;
        RECT 235.275 37.015 240.830 37.020 ;
        POLYGON 240.830 37.125 241.010 37.015 240.830 37.015 ;
        POLYGON 257.500 37.125 257.500 37.065 257.415 37.065 ;
        RECT 257.500 37.065 261.950 37.125 ;
        POLYGON 261.950 37.205 262.085 37.205 261.950 37.065 ;
        POLYGON 267.945 37.205 267.945 37.120 267.900 37.120 ;
        RECT 267.945 37.120 276.115 37.205 ;
        POLYGON 267.900 37.120 267.900 37.065 267.865 37.065 ;
        RECT 267.900 37.065 276.115 37.120 ;
        POLYGON 257.415 37.065 257.415 37.015 257.345 37.015 ;
        RECT 257.415 37.015 261.690 37.065 ;
        RECT 235.275 36.985 241.010 37.015 ;
        POLYGON 235.275 36.985 235.560 36.985 235.560 36.710 ;
        RECT 235.560 36.825 241.010 36.985 ;
        POLYGON 241.010 37.015 241.315 36.825 241.010 36.825 ;
        POLYGON 257.345 37.015 257.345 36.905 257.165 36.905 ;
        RECT 257.345 36.905 261.690 37.015 ;
        POLYGON 257.165 36.905 257.165 36.825 257.040 36.825 ;
        RECT 257.165 36.825 261.690 36.905 ;
        RECT 235.560 36.810 241.315 36.825 ;
        POLYGON 241.315 36.825 241.335 36.810 241.315 36.810 ;
        POLYGON 257.040 36.825 257.040 36.810 257.015 36.810 ;
        RECT 257.040 36.810 261.690 36.825 ;
        POLYGON 261.690 37.065 261.950 37.065 261.690 36.810 ;
        POLYGON 267.865 37.065 267.865 36.930 267.780 36.930 ;
        RECT 267.865 36.930 276.115 37.065 ;
        POLYGON 267.780 36.930 267.780 36.810 267.705 36.810 ;
        RECT 267.780 36.810 276.115 36.930 ;
        RECT 235.560 36.735 241.335 36.810 ;
        POLYGON 241.335 36.810 241.475 36.735 241.335 36.735 ;
        POLYGON 257.015 36.810 257.015 36.735 256.875 36.735 ;
        RECT 257.015 36.735 261.070 36.810 ;
        RECT 235.560 36.710 241.480 36.735 ;
        RECT 212.275 36.705 227.295 36.710 ;
        POLYGON 227.295 36.710 227.300 36.705 227.295 36.705 ;
        POLYGON 235.560 36.710 235.565 36.710 235.565 36.705 ;
        RECT 235.565 36.705 241.480 36.710 ;
        RECT 212.275 36.410 227.300 36.705 ;
        POLYGON 227.300 36.705 227.520 36.410 227.300 36.410 ;
        POLYGON 235.565 36.705 235.765 36.705 235.765 36.515 ;
        RECT 235.765 36.605 241.480 36.705 ;
        POLYGON 241.480 36.735 241.710 36.605 241.480 36.605 ;
        POLYGON 256.875 36.735 256.875 36.650 256.720 36.650 ;
        RECT 256.875 36.650 261.070 36.735 ;
        POLYGON 256.720 36.650 256.720 36.605 256.635 36.605 ;
        RECT 256.720 36.605 261.070 36.650 ;
        RECT 235.765 36.515 241.710 36.605 ;
        POLYGON 235.765 36.515 235.885 36.515 235.885 36.410 ;
        RECT 235.885 36.420 241.710 36.515 ;
        POLYGON 241.710 36.605 242.050 36.420 241.710 36.420 ;
        POLYGON 256.635 36.605 256.635 36.555 256.540 36.555 ;
        RECT 256.635 36.555 261.070 36.605 ;
        POLYGON 256.540 36.555 256.540 36.455 256.360 36.455 ;
        RECT 256.540 36.455 261.070 36.555 ;
        POLYGON 256.360 36.455 256.360 36.450 256.355 36.450 ;
        RECT 256.360 36.450 261.070 36.455 ;
        POLYGON 256.355 36.450 256.355 36.420 256.290 36.420 ;
        RECT 256.355 36.420 261.070 36.450 ;
        RECT 235.885 36.410 242.050 36.420 ;
        RECT 212.275 36.000 227.520 36.410 ;
        POLYGON 227.520 36.410 227.830 36.000 227.520 36.000 ;
        POLYGON 235.885 36.410 236.005 36.410 236.005 36.305 ;
        RECT 236.005 36.305 242.050 36.410 ;
        POLYGON 236.005 36.305 236.345 36.305 236.345 36.000 ;
        RECT 236.345 36.255 242.050 36.305 ;
        POLYGON 242.050 36.420 242.380 36.255 242.050 36.255 ;
        POLYGON 256.290 36.420 256.290 36.405 256.255 36.405 ;
        RECT 256.290 36.405 261.070 36.420 ;
        POLYGON 256.255 36.405 256.255 36.255 255.935 36.255 ;
        RECT 256.255 36.255 261.070 36.405 ;
        RECT 236.345 36.230 242.385 36.255 ;
        POLYGON 242.385 36.255 242.440 36.230 242.385 36.230 ;
        POLYGON 255.935 36.255 255.935 36.230 255.880 36.230 ;
        RECT 255.935 36.230 261.070 36.255 ;
        RECT 236.345 36.060 242.440 36.230 ;
        POLYGON 242.440 36.230 242.785 36.060 242.440 36.060 ;
        POLYGON 255.880 36.230 255.880 36.180 255.775 36.180 ;
        RECT 255.880 36.210 261.070 36.230 ;
        POLYGON 261.070 36.810 261.690 36.810 261.070 36.210 ;
        POLYGON 267.705 36.810 267.705 36.710 267.645 36.710 ;
        RECT 267.705 36.710 276.115 36.810 ;
        POLYGON 267.645 36.710 267.645 36.210 267.295 36.210 ;
        RECT 267.645 36.435 276.115 36.710 ;
        POLYGON 276.115 37.205 276.380 37.205 276.115 36.435 ;
        POLYGON 287.425 37.205 287.425 36.440 287.385 36.440 ;
        RECT 287.425 36.440 303.120 37.215 ;
        RECT 267.645 36.210 275.725 36.435 ;
        RECT 255.880 36.180 260.970 36.210 ;
        POLYGON 255.775 36.180 255.775 36.155 255.720 36.155 ;
        RECT 255.775 36.155 260.970 36.180 ;
        POLYGON 255.720 36.155 255.720 36.115 255.630 36.115 ;
        RECT 255.720 36.125 260.970 36.155 ;
        POLYGON 260.970 36.210 261.070 36.210 260.970 36.125 ;
        POLYGON 267.295 36.210 267.295 36.165 267.265 36.165 ;
        RECT 267.295 36.165 275.725 36.210 ;
        POLYGON 267.265 36.165 267.265 36.125 267.235 36.125 ;
        RECT 267.265 36.125 275.725 36.165 ;
        RECT 255.720 36.115 260.585 36.125 ;
        POLYGON 255.630 36.115 255.630 36.060 255.495 36.060 ;
        RECT 255.630 36.060 260.585 36.115 ;
        RECT 236.345 36.020 242.785 36.060 ;
        POLYGON 242.785 36.060 242.885 36.020 242.785 36.020 ;
        POLYGON 255.495 36.060 255.495 36.020 255.395 36.020 ;
        RECT 255.495 36.020 260.585 36.060 ;
        RECT 236.345 36.000 242.885 36.020 ;
        RECT 212.275 35.925 227.830 36.000 ;
        POLYGON 227.830 36.000 227.890 35.925 227.830 35.925 ;
        POLYGON 236.345 36.000 236.390 36.000 236.390 35.960 ;
        RECT 236.390 35.960 242.885 36.000 ;
        POLYGON 236.390 35.960 236.430 35.960 236.430 35.925 ;
        RECT 236.430 35.925 242.885 35.960 ;
        RECT 212.275 35.690 227.890 35.925 ;
        POLYGON 212.275 35.690 212.325 35.690 212.325 35.600 ;
        RECT 212.325 35.600 227.890 35.690 ;
        POLYGON 212.325 35.600 212.395 35.600 212.395 35.485 ;
        RECT 212.395 35.485 227.890 35.600 ;
        RECT 180.810 35.320 197.510 35.485 ;
        POLYGON 180.685 35.320 180.685 35.220 180.645 35.220 ;
        RECT 180.685 35.220 197.510 35.320 ;
        POLYGON 180.645 35.220 180.645 35.090 180.585 35.090 ;
        RECT 180.645 35.090 197.510 35.220 ;
        RECT 164.845 35.045 171.285 35.090 ;
        RECT 117.885 35.000 156.975 35.045 ;
        POLYGON 156.975 35.045 157.270 35.045 156.975 35.000 ;
        POLYGON 164.750 35.045 164.750 35.000 164.690 35.000 ;
        RECT 164.750 35.000 171.285 35.045 ;
        RECT 117.885 34.925 156.490 35.000 ;
        POLYGON 156.490 35.000 156.975 35.000 156.490 34.925 ;
        POLYGON 164.690 35.000 164.690 34.925 164.590 34.925 ;
        RECT 164.690 34.925 171.285 35.000 ;
        RECT 117.885 34.900 156.240 34.925 ;
        POLYGON 156.240 34.925 156.445 34.925 156.240 34.900 ;
        POLYGON 164.590 34.925 164.590 34.900 164.555 34.900 ;
        RECT 164.590 34.915 171.285 34.925 ;
        POLYGON 171.285 35.090 171.435 35.090 171.285 34.915 ;
        POLYGON 180.585 35.085 180.585 34.920 180.510 34.920 ;
        RECT 180.585 34.950 197.510 35.090 ;
        POLYGON 197.510 35.485 197.580 35.485 197.510 34.950 ;
        POLYGON 212.395 35.485 212.410 35.485 212.410 35.460 ;
        RECT 212.410 35.455 227.890 35.485 ;
        POLYGON 227.890 35.925 228.270 35.455 227.890 35.455 ;
        POLYGON 236.430 35.925 236.610 35.925 236.610 35.780 ;
        RECT 236.610 35.890 242.885 35.925 ;
        POLYGON 242.885 36.020 243.190 35.890 242.885 35.890 ;
        POLYGON 255.395 36.020 255.395 35.980 255.295 35.980 ;
        RECT 255.395 35.980 260.585 36.020 ;
        POLYGON 255.290 35.980 255.290 35.975 255.280 35.975 ;
        RECT 255.290 35.975 260.585 35.980 ;
        POLYGON 255.280 35.975 255.280 35.890 255.070 35.890 ;
        RECT 255.280 35.890 260.585 35.975 ;
        RECT 236.610 35.780 243.190 35.890 ;
        POLYGON 236.610 35.780 236.875 35.780 236.875 35.560 ;
        RECT 236.875 35.775 243.190 35.780 ;
        POLYGON 243.190 35.890 243.455 35.775 243.190 35.775 ;
        POLYGON 255.070 35.890 255.070 35.815 254.885 35.815 ;
        RECT 255.070 35.815 260.585 35.890 ;
        POLYGON 254.885 35.815 254.885 35.810 254.870 35.810 ;
        RECT 254.885 35.810 260.585 35.815 ;
        POLYGON 254.870 35.810 254.870 35.780 254.770 35.780 ;
        RECT 254.870 35.790 260.585 35.810 ;
        POLYGON 260.585 36.125 260.970 36.125 260.585 35.790 ;
        POLYGON 267.235 36.125 267.235 35.835 267.015 35.835 ;
        RECT 267.235 35.835 275.725 36.125 ;
        POLYGON 267.015 35.835 267.015 35.790 266.980 35.790 ;
        RECT 267.015 35.790 275.725 35.835 ;
        RECT 254.870 35.780 260.195 35.790 ;
        POLYGON 254.770 35.780 254.770 35.775 254.755 35.775 ;
        RECT 254.770 35.775 260.195 35.780 ;
        RECT 236.875 35.740 243.455 35.775 ;
        POLYGON 243.455 35.775 243.540 35.740 243.455 35.740 ;
        POLYGON 254.755 35.775 254.755 35.740 254.650 35.740 ;
        RECT 254.755 35.740 260.195 35.775 ;
        RECT 236.875 35.700 243.540 35.740 ;
        POLYGON 243.540 35.740 243.640 35.700 243.540 35.700 ;
        POLYGON 254.650 35.740 254.650 35.700 254.535 35.700 ;
        RECT 254.650 35.700 260.195 35.740 ;
        RECT 236.875 35.585 243.645 35.700 ;
        POLYGON 243.645 35.700 243.960 35.585 243.645 35.585 ;
        POLYGON 254.535 35.700 254.535 35.595 254.225 35.595 ;
        RECT 254.535 35.595 260.195 35.700 ;
        POLYGON 254.225 35.595 254.225 35.585 254.200 35.585 ;
        RECT 254.225 35.585 260.195 35.595 ;
        RECT 236.875 35.560 243.960 35.585 ;
        POLYGON 236.875 35.560 237.000 35.560 237.000 35.455 ;
        RECT 237.000 35.455 243.960 35.560 ;
        POLYGON 243.960 35.585 244.310 35.455 243.960 35.455 ;
        POLYGON 254.200 35.585 254.200 35.545 254.090 35.545 ;
        RECT 254.200 35.545 260.195 35.585 ;
        POLYGON 254.090 35.545 254.090 35.535 254.045 35.535 ;
        RECT 254.090 35.535 260.195 35.545 ;
        POLYGON 254.045 35.535 254.045 35.455 253.760 35.455 ;
        RECT 254.045 35.455 260.195 35.535 ;
        POLYGON 260.195 35.790 260.585 35.790 260.195 35.455 ;
        POLYGON 266.980 35.785 266.980 35.780 266.975 35.780 ;
        RECT 266.980 35.780 275.725 35.790 ;
        POLYGON 266.975 35.780 266.975 35.645 266.870 35.645 ;
        RECT 266.975 35.645 275.725 35.780 ;
        POLYGON 266.870 35.645 266.870 35.595 266.830 35.595 ;
        RECT 266.870 35.595 275.725 35.645 ;
        POLYGON 266.830 35.595 266.830 35.485 266.740 35.485 ;
        RECT 266.830 35.485 275.725 35.595 ;
        POLYGON 266.740 35.485 266.740 35.470 266.725 35.470 ;
        RECT 266.740 35.470 275.725 35.485 ;
        POLYGON 266.725 35.470 266.725 35.455 266.715 35.455 ;
        RECT 266.725 35.455 275.725 35.470 ;
        POLYGON 275.725 36.435 276.115 36.435 275.725 35.460 ;
        POLYGON 287.385 36.435 287.385 35.485 287.335 35.485 ;
        RECT 287.385 35.485 303.120 36.440 ;
        POLYGON 212.410 35.455 212.530 35.455 212.530 35.260 ;
        RECT 212.530 35.315 228.270 35.455 ;
        POLYGON 228.270 35.455 228.385 35.315 228.270 35.315 ;
        POLYGON 237.000 35.455 237.025 35.455 237.025 35.435 ;
        RECT 237.025 35.435 244.310 35.455 ;
        POLYGON 237.025 35.435 237.180 35.435 237.180 35.315 ;
        RECT 237.180 35.415 244.310 35.435 ;
        POLYGON 244.310 35.455 244.440 35.415 244.310 35.415 ;
        POLYGON 253.760 35.455 253.760 35.415 253.615 35.415 ;
        RECT 253.760 35.415 260.145 35.455 ;
        RECT 237.180 35.390 244.440 35.415 ;
        POLYGON 244.440 35.415 244.525 35.390 244.440 35.390 ;
        POLYGON 253.615 35.415 253.615 35.390 253.530 35.390 ;
        RECT 253.615 35.410 260.145 35.415 ;
        POLYGON 260.145 35.455 260.195 35.455 260.145 35.410 ;
        POLYGON 266.715 35.455 266.715 35.430 266.695 35.430 ;
        RECT 266.715 35.430 275.645 35.455 ;
        POLYGON 266.695 35.430 266.695 35.410 266.680 35.410 ;
        RECT 266.695 35.410 275.645 35.430 ;
        RECT 253.615 35.390 259.955 35.410 ;
        RECT 237.180 35.340 244.530 35.390 ;
        POLYGON 244.530 35.390 244.675 35.340 244.530 35.340 ;
        POLYGON 253.530 35.390 253.530 35.385 253.510 35.385 ;
        RECT 253.530 35.385 259.955 35.390 ;
        POLYGON 253.505 35.385 253.505 35.340 253.355 35.340 ;
        RECT 253.505 35.340 259.955 35.385 ;
        RECT 237.180 35.320 244.675 35.340 ;
        POLYGON 244.675 35.340 244.750 35.320 244.675 35.320 ;
        POLYGON 253.355 35.340 253.355 35.320 253.285 35.320 ;
        RECT 253.355 35.320 259.955 35.340 ;
        RECT 237.180 35.315 244.750 35.320 ;
        RECT 212.530 35.260 228.385 35.315 ;
        POLYGON 228.385 35.315 228.430 35.260 228.385 35.260 ;
        POLYGON 237.180 35.315 237.250 35.315 237.250 35.260 ;
        RECT 237.250 35.260 244.750 35.315 ;
        POLYGON 244.750 35.320 244.955 35.260 244.750 35.260 ;
        POLYGON 253.285 35.320 253.285 35.310 253.235 35.310 ;
        RECT 253.285 35.310 259.955 35.320 ;
        POLYGON 253.235 35.310 253.235 35.300 253.195 35.300 ;
        RECT 253.235 35.300 259.955 35.310 ;
        POLYGON 253.190 35.300 253.190 35.290 253.155 35.290 ;
        RECT 253.190 35.290 259.955 35.300 ;
        POLYGON 253.150 35.290 253.150 35.260 253.015 35.260 ;
        RECT 253.150 35.260 259.955 35.290 ;
        POLYGON 259.955 35.410 260.145 35.410 259.955 35.260 ;
        POLYGON 266.680 35.410 266.680 35.365 266.645 35.365 ;
        RECT 266.680 35.365 275.645 35.410 ;
        POLYGON 266.645 35.365 266.645 35.275 266.570 35.275 ;
        RECT 266.645 35.275 275.645 35.365 ;
        POLYGON 266.570 35.275 266.570 35.265 266.560 35.265 ;
        RECT 266.570 35.265 275.645 35.275 ;
        RECT 266.560 35.260 275.645 35.265 ;
        POLYGON 275.645 35.455 275.725 35.455 275.645 35.260 ;
        POLYGON 287.335 35.455 287.335 35.260 287.325 35.260 ;
        RECT 287.335 35.260 303.120 35.485 ;
        POLYGON 212.530 35.260 212.720 35.260 212.720 34.950 ;
        RECT 212.720 35.150 228.430 35.260 ;
        POLYGON 228.430 35.260 228.525 35.150 228.430 35.150 ;
        POLYGON 237.250 35.260 237.395 35.260 237.395 35.150 ;
        RECT 237.395 35.235 244.955 35.260 ;
        POLYGON 244.955 35.260 245.045 35.235 244.955 35.235 ;
        POLYGON 253.015 35.260 253.015 35.250 252.970 35.250 ;
        RECT 253.015 35.250 259.820 35.260 ;
        POLYGON 252.970 35.250 252.970 35.235 252.905 35.235 ;
        RECT 252.970 35.235 259.820 35.250 ;
        RECT 237.395 35.225 245.045 35.235 ;
        POLYGON 245.045 35.235 245.095 35.225 245.045 35.225 ;
        POLYGON 252.905 35.235 252.905 35.225 252.860 35.225 ;
        RECT 252.905 35.225 259.820 35.235 ;
        RECT 237.395 35.150 245.095 35.225 ;
        POLYGON 245.095 35.225 245.385 35.150 245.095 35.150 ;
        POLYGON 252.860 35.225 252.860 35.190 252.710 35.190 ;
        RECT 252.860 35.190 259.820 35.225 ;
        POLYGON 252.705 35.190 252.705 35.150 252.540 35.150 ;
        RECT 252.705 35.155 259.820 35.190 ;
        POLYGON 259.820 35.260 259.955 35.260 259.820 35.155 ;
        POLYGON 266.560 35.260 266.560 35.160 266.475 35.160 ;
        RECT 266.560 35.235 275.635 35.260 ;
        POLYGON 275.635 35.260 275.645 35.260 275.635 35.235 ;
        POLYGON 287.325 35.260 287.325 35.235 287.320 35.235 ;
        RECT 287.325 35.235 303.120 35.260 ;
        RECT 266.560 35.160 275.495 35.235 ;
        POLYGON 266.475 35.160 266.475 35.155 266.470 35.155 ;
        RECT 266.475 35.155 275.495 35.160 ;
        RECT 252.705 35.150 259.530 35.155 ;
        RECT 212.720 34.950 228.525 35.150 ;
        RECT 180.585 34.920 197.100 34.950 ;
        RECT 164.590 34.900 171.065 34.915 ;
        RECT 117.885 34.885 156.115 34.900 ;
        POLYGON 156.115 34.900 156.235 34.900 156.115 34.885 ;
        POLYGON 164.555 34.900 164.555 34.885 164.535 34.885 ;
        RECT 164.555 34.885 171.065 34.900 ;
        RECT 117.885 34.830 155.685 34.885 ;
        POLYGON 155.685 34.885 156.115 34.885 155.685 34.840 ;
        POLYGON 164.535 34.885 164.535 34.875 164.520 34.875 ;
        RECT 164.535 34.875 171.065 34.885 ;
        POLYGON 164.520 34.875 164.520 34.860 164.505 34.860 ;
        RECT 164.520 34.860 171.065 34.875 ;
        POLYGON 164.505 34.860 164.505 34.840 164.475 34.840 ;
        RECT 164.505 34.840 171.065 34.860 ;
        POLYGON 164.475 34.840 164.475 34.835 164.470 34.835 ;
        RECT 164.475 34.835 171.065 34.840 ;
        POLYGON 155.685 34.835 155.690 34.830 155.685 34.830 ;
        POLYGON 164.470 34.835 164.470 34.830 164.460 34.830 ;
        RECT 164.470 34.830 171.065 34.835 ;
        RECT 117.885 34.815 155.690 34.830 ;
        POLYGON 155.690 34.830 155.700 34.815 155.690 34.815 ;
        POLYGON 164.460 34.830 164.460 34.815 164.440 34.815 ;
        RECT 164.460 34.815 171.065 34.830 ;
        RECT 117.885 34.790 155.700 34.815 ;
        POLYGON 155.700 34.815 155.715 34.790 155.700 34.790 ;
        POLYGON 164.440 34.815 164.440 34.790 164.400 34.790 ;
        RECT 164.440 34.790 171.065 34.815 ;
        RECT 117.885 34.780 155.715 34.790 ;
        POLYGON 155.715 34.790 155.720 34.780 155.715 34.780 ;
        RECT 60.990 34.600 117.775 34.780 ;
        POLYGON 117.775 34.780 117.885 34.600 117.775 34.600 ;
        POLYGON 117.885 34.780 117.910 34.780 117.910 34.610 ;
        RECT 117.910 34.655 155.720 34.780 ;
        POLYGON 164.400 34.790 164.400 34.775 164.380 34.775 ;
        RECT 164.400 34.775 171.065 34.790 ;
        POLYGON 155.720 34.775 155.795 34.655 155.720 34.655 ;
        RECT 117.910 34.640 155.795 34.655 ;
        POLYGON 164.380 34.775 164.380 34.650 164.195 34.650 ;
        RECT 164.380 34.665 171.065 34.775 ;
        POLYGON 171.065 34.915 171.285 34.915 171.065 34.665 ;
        POLYGON 180.510 34.915 180.510 34.720 180.420 34.720 ;
        RECT 180.510 34.720 197.100 34.920 ;
        POLYGON 180.420 34.720 180.420 34.665 180.395 34.665 ;
        RECT 180.420 34.665 197.100 34.720 ;
        RECT 164.380 34.650 170.455 34.665 ;
        POLYGON 155.795 34.650 155.805 34.640 155.795 34.640 ;
        POLYGON 164.195 34.650 164.195 34.640 164.180 34.640 ;
        RECT 164.195 34.640 170.455 34.650 ;
        RECT 117.910 34.605 155.805 34.640 ;
        POLYGON 155.805 34.640 155.825 34.605 155.805 34.605 ;
        POLYGON 164.180 34.640 164.180 34.605 164.130 34.605 ;
        RECT 164.180 34.605 170.455 34.640 ;
        RECT 117.910 34.600 155.825 34.605 ;
        RECT 60.990 34.560 117.885 34.600 ;
        POLYGON 117.885 34.600 117.910 34.560 117.885 34.560 ;
        POLYGON 117.910 34.600 117.915 34.600 117.915 34.570 ;
        RECT 60.990 34.550 117.910 34.560 ;
        POLYGON 117.910 34.560 117.915 34.550 117.910 34.550 ;
        RECT 117.915 34.550 155.825 34.600 ;
        RECT 60.990 34.520 155.825 34.550 ;
        POLYGON 155.825 34.605 155.875 34.520 155.825 34.520 ;
        RECT 60.990 34.485 155.875 34.520 ;
        POLYGON 164.130 34.605 164.130 34.515 164.000 34.515 ;
        RECT 164.130 34.515 170.455 34.605 ;
        POLYGON 155.875 34.515 155.895 34.485 155.875 34.485 ;
        POLYGON 164.000 34.515 164.000 34.485 163.950 34.485 ;
        RECT 164.000 34.485 170.455 34.515 ;
        RECT 60.990 34.480 155.895 34.485 ;
        POLYGON 155.895 34.485 155.900 34.480 155.895 34.480 ;
        RECT 60.990 34.445 155.900 34.480 ;
        POLYGON 163.950 34.485 163.950 34.475 163.940 34.475 ;
        RECT 163.950 34.475 170.455 34.485 ;
        POLYGON 155.900 34.475 155.920 34.445 155.900 34.445 ;
        RECT 60.990 34.380 155.920 34.445 ;
        POLYGON 163.940 34.475 163.940 34.440 163.885 34.440 ;
        RECT 163.940 34.440 170.455 34.475 ;
        POLYGON 155.920 34.440 155.960 34.380 155.920 34.380 ;
        POLYGON 163.885 34.440 163.885 34.380 163.790 34.380 ;
        RECT 163.885 34.380 170.455 34.440 ;
        RECT 60.990 34.235 155.960 34.380 ;
        POLYGON 155.960 34.380 156.045 34.235 155.960 34.235 ;
        RECT 60.990 34.200 156.045 34.235 ;
        POLYGON 163.790 34.380 163.790 34.230 163.555 34.230 ;
        RECT 163.790 34.230 170.455 34.380 ;
        POLYGON 60.990 34.200 62.050 34.200 62.050 32.460 ;
        RECT 62.050 34.125 156.045 34.200 ;
        POLYGON 156.045 34.230 156.110 34.125 156.045 34.125 ;
        POLYGON 163.555 34.230 163.555 34.125 163.390 34.125 ;
        RECT 163.555 34.125 170.455 34.230 ;
        RECT 62.050 34.120 156.110 34.125 ;
        POLYGON 156.110 34.125 156.115 34.120 156.110 34.120 ;
        POLYGON 163.390 34.125 163.390 34.120 163.380 34.120 ;
        RECT 163.390 34.120 170.455 34.125 ;
        RECT 62.050 34.100 156.115 34.120 ;
        POLYGON 156.115 34.120 156.125 34.100 156.115 34.100 ;
        POLYGON 163.380 34.120 163.380 34.110 163.365 34.110 ;
        RECT 163.380 34.110 170.455 34.120 ;
        POLYGON 163.365 34.110 163.365 34.100 163.350 34.100 ;
        RECT 163.365 34.100 170.455 34.110 ;
        RECT 62.050 33.965 156.125 34.100 ;
        POLYGON 156.125 34.100 156.215 33.965 156.125 33.965 ;
        RECT 62.050 33.855 156.215 33.965 ;
        POLYGON 163.350 34.100 163.350 33.960 163.105 33.960 ;
        RECT 163.350 33.970 170.455 34.100 ;
        POLYGON 170.455 34.665 171.065 34.665 170.455 33.970 ;
        POLYGON 180.395 34.665 180.395 34.040 180.110 34.040 ;
        RECT 180.395 34.040 197.100 34.665 ;
        POLYGON 180.110 34.040 180.110 33.995 180.085 33.995 ;
        RECT 180.110 33.995 197.100 34.040 ;
        POLYGON 180.085 33.995 180.085 33.970 180.070 33.970 ;
        RECT 180.085 33.970 197.100 33.995 ;
        RECT 163.350 33.960 169.875 33.970 ;
        POLYGON 156.215 33.960 156.285 33.855 156.215 33.855 ;
        POLYGON 163.105 33.960 163.105 33.855 162.930 33.855 ;
        RECT 163.105 33.855 169.875 33.960 ;
        RECT 62.050 33.850 156.285 33.855 ;
        POLYGON 156.285 33.855 156.290 33.850 156.285 33.850 ;
        POLYGON 162.930 33.855 162.930 33.850 162.920 33.850 ;
        RECT 162.930 33.850 169.875 33.855 ;
        RECT 62.050 33.790 156.290 33.850 ;
        POLYGON 156.290 33.850 156.330 33.790 156.290 33.790 ;
        RECT 62.050 33.750 156.330 33.790 ;
        POLYGON 162.920 33.850 162.920 33.785 162.810 33.785 ;
        RECT 162.920 33.785 169.875 33.850 ;
        POLYGON 156.330 33.785 156.355 33.750 156.330 33.750 ;
        POLYGON 162.810 33.785 162.810 33.750 162.740 33.750 ;
        RECT 162.810 33.750 169.875 33.785 ;
        RECT 62.050 33.615 156.355 33.750 ;
        POLYGON 156.355 33.750 156.445 33.615 156.355 33.615 ;
        POLYGON 162.740 33.750 162.740 33.615 162.490 33.615 ;
        RECT 162.740 33.615 169.875 33.750 ;
        RECT 62.050 33.590 156.445 33.615 ;
        POLYGON 162.490 33.615 162.490 33.610 162.480 33.610 ;
        RECT 162.490 33.610 169.875 33.615 ;
        POLYGON 156.445 33.610 156.460 33.590 156.445 33.590 ;
        RECT 62.050 33.505 156.460 33.590 ;
        POLYGON 162.480 33.610 162.480 33.585 162.435 33.585 ;
        RECT 162.480 33.585 169.875 33.610 ;
        POLYGON 156.460 33.585 156.515 33.505 156.460 33.505 ;
        POLYGON 162.435 33.585 162.435 33.505 162.285 33.505 ;
        RECT 162.435 33.505 169.875 33.585 ;
        RECT 62.050 33.470 156.515 33.505 ;
        POLYGON 156.515 33.505 156.540 33.470 156.515 33.470 ;
        POLYGON 162.285 33.505 162.285 33.470 162.220 33.470 ;
        RECT 162.285 33.470 169.875 33.505 ;
        RECT 62.050 33.425 156.540 33.470 ;
        POLYGON 156.540 33.470 156.570 33.425 156.540 33.425 ;
        RECT 62.050 33.385 156.570 33.425 ;
        POLYGON 162.220 33.470 162.220 33.420 162.120 33.420 ;
        RECT 162.220 33.420 169.875 33.470 ;
        POLYGON 156.570 33.420 156.595 33.385 156.570 33.385 ;
        POLYGON 162.120 33.420 162.120 33.385 162.055 33.385 ;
        RECT 162.120 33.385 169.875 33.420 ;
        RECT 62.050 33.380 156.595 33.385 ;
        POLYGON 156.595 33.385 156.600 33.380 156.595 33.380 ;
        RECT 62.050 33.265 156.600 33.380 ;
        POLYGON 162.055 33.385 162.055 33.375 162.035 33.375 ;
        RECT 162.055 33.375 169.875 33.385 ;
        POLYGON 156.600 33.375 156.675 33.265 156.600 33.265 ;
        POLYGON 162.035 33.375 162.035 33.265 161.805 33.265 ;
        RECT 162.035 33.365 169.875 33.375 ;
        POLYGON 169.875 33.970 170.455 33.970 169.875 33.365 ;
        POLYGON 180.070 33.965 180.070 33.370 179.760 33.370 ;
        RECT 180.070 33.370 197.100 33.970 ;
        RECT 162.035 33.265 169.375 33.365 ;
        RECT 62.050 33.205 156.675 33.265 ;
        POLYGON 156.675 33.265 156.715 33.205 156.675 33.205 ;
        RECT 62.050 33.175 156.715 33.205 ;
        POLYGON 161.805 33.265 161.805 33.200 161.670 33.200 ;
        RECT 161.805 33.200 169.375 33.265 ;
        POLYGON 156.715 33.200 156.735 33.175 156.715 33.175 ;
        POLYGON 161.670 33.200 161.670 33.175 161.620 33.175 ;
        RECT 161.670 33.175 169.375 33.200 ;
        RECT 62.050 33.115 156.735 33.175 ;
        POLYGON 156.735 33.175 156.775 33.115 156.735 33.115 ;
        POLYGON 161.620 33.175 161.620 33.145 161.555 33.145 ;
        RECT 161.620 33.145 169.375 33.175 ;
        POLYGON 161.555 33.145 161.555 33.115 161.485 33.115 ;
        RECT 161.555 33.115 169.375 33.145 ;
        RECT 62.050 32.975 156.775 33.115 ;
        POLYGON 156.775 33.115 156.865 32.975 156.775 32.975 ;
        POLYGON 161.485 33.115 161.485 32.975 161.175 32.975 ;
        RECT 161.485 32.975 169.375 33.115 ;
        RECT 62.050 32.940 156.865 32.975 ;
        POLYGON 156.865 32.975 156.890 32.940 156.865 32.940 ;
        RECT 62.050 32.900 156.890 32.940 ;
        POLYGON 161.175 32.975 161.175 32.935 161.085 32.935 ;
        RECT 161.175 32.935 169.375 32.975 ;
        POLYGON 156.890 32.935 156.915 32.900 156.890 32.900 ;
        POLYGON 161.085 32.935 161.085 32.900 161.010 32.900 ;
        RECT 161.085 32.900 169.375 32.935 ;
        RECT 62.050 32.895 156.915 32.900 ;
        POLYGON 156.915 32.900 156.920 32.895 156.915 32.895 ;
        RECT 62.050 32.885 156.920 32.895 ;
        POLYGON 161.010 32.900 161.010 32.890 160.985 32.890 ;
        RECT 161.010 32.890 169.375 32.900 ;
        POLYGON 156.920 32.890 156.925 32.885 156.920 32.885 ;
        POLYGON 160.985 32.890 160.985 32.885 160.970 32.885 ;
        RECT 160.985 32.885 169.375 32.890 ;
        RECT 62.050 32.825 156.925 32.885 ;
        POLYGON 156.925 32.885 156.965 32.825 156.925 32.825 ;
        POLYGON 160.970 32.885 160.970 32.825 160.830 32.825 ;
        RECT 160.970 32.845 169.375 32.885 ;
        POLYGON 169.375 33.365 169.875 33.365 169.375 32.845 ;
        POLYGON 179.760 33.365 179.760 32.885 179.510 32.885 ;
        RECT 179.760 32.885 197.100 33.370 ;
        POLYGON 179.510 32.885 179.510 32.845 179.485 32.845 ;
        RECT 179.510 32.845 197.100 32.885 ;
        RECT 160.970 32.825 168.875 32.845 ;
        RECT 62.050 32.800 156.965 32.825 ;
        POLYGON 156.965 32.825 156.980 32.800 156.965 32.800 ;
        POLYGON 160.830 32.825 160.830 32.800 160.770 32.800 ;
        RECT 160.830 32.800 168.875 32.825 ;
        RECT 62.050 32.705 156.980 32.800 ;
        POLYGON 156.980 32.800 157.045 32.705 156.980 32.705 ;
        RECT 62.050 32.645 157.045 32.705 ;
        POLYGON 160.770 32.800 160.770 32.700 160.520 32.700 ;
        RECT 160.770 32.700 168.875 32.800 ;
        POLYGON 157.045 32.700 157.085 32.645 157.045 32.645 ;
        POLYGON 160.520 32.700 160.520 32.645 160.390 32.645 ;
        RECT 160.520 32.645 168.875 32.700 ;
        RECT 62.050 32.630 157.085 32.645 ;
        POLYGON 157.085 32.645 157.095 32.630 157.085 32.630 ;
        RECT 62.050 32.560 157.095 32.630 ;
        POLYGON 160.390 32.645 160.390 32.625 160.335 32.625 ;
        RECT 160.390 32.625 168.875 32.645 ;
        POLYGON 157.095 32.625 157.140 32.560 157.095 32.560 ;
        POLYGON 160.335 32.625 160.335 32.560 160.160 32.560 ;
        RECT 160.335 32.560 168.875 32.625 ;
        RECT 62.050 32.555 157.140 32.560 ;
        POLYGON 157.140 32.560 157.145 32.555 157.140 32.555 ;
        RECT 62.050 32.530 157.145 32.555 ;
        POLYGON 160.160 32.560 160.160 32.550 160.130 32.550 ;
        RECT 160.160 32.550 168.875 32.560 ;
        POLYGON 157.145 32.550 157.160 32.530 157.145 32.530 ;
        RECT 62.050 32.470 157.160 32.530 ;
        POLYGON 160.130 32.550 160.130 32.525 160.065 32.525 ;
        RECT 160.130 32.525 168.875 32.550 ;
        POLYGON 157.160 32.525 157.200 32.470 157.160 32.470 ;
        POLYGON 160.065 32.525 160.065 32.470 159.910 32.470 ;
        RECT 160.065 32.470 168.875 32.525 ;
        RECT 62.050 32.460 157.200 32.470 ;
        POLYGON 62.050 32.460 63.450 32.460 63.450 30.405 ;
        RECT 63.450 32.455 157.200 32.460 ;
        POLYGON 157.200 32.470 157.210 32.455 157.200 32.455 ;
        POLYGON 159.910 32.470 159.910 32.455 159.870 32.455 ;
        RECT 159.910 32.455 168.875 32.470 ;
        RECT 63.450 32.445 157.210 32.455 ;
        POLYGON 157.210 32.450 157.215 32.445 157.210 32.445 ;
        POLYGON 159.865 32.450 159.865 32.445 159.845 32.445 ;
        RECT 159.865 32.445 168.875 32.455 ;
        RECT 63.450 32.415 157.215 32.445 ;
        POLYGON 157.215 32.445 157.235 32.415 157.215 32.415 ;
        POLYGON 159.845 32.445 159.845 32.415 159.760 32.415 ;
        RECT 159.845 32.415 168.875 32.445 ;
        RECT 63.450 32.380 157.235 32.415 ;
        POLYGON 157.235 32.415 157.260 32.380 157.235 32.380 ;
        RECT 63.450 32.320 157.260 32.380 ;
        POLYGON 159.760 32.415 159.760 32.375 159.640 32.375 ;
        RECT 159.760 32.375 168.875 32.415 ;
        POLYGON 157.260 32.375 157.300 32.320 157.260 32.320 ;
        POLYGON 159.640 32.375 159.640 32.320 159.470 32.320 ;
        RECT 159.640 32.365 168.875 32.375 ;
        POLYGON 168.875 32.845 169.375 32.845 168.875 32.365 ;
        POLYGON 179.485 32.840 179.485 32.710 179.410 32.710 ;
        RECT 179.485 32.710 197.100 32.845 ;
        POLYGON 179.410 32.710 179.410 32.365 179.210 32.365 ;
        RECT 179.410 32.700 197.100 32.710 ;
        POLYGON 197.100 34.950 197.510 34.950 197.100 32.700 ;
        POLYGON 212.720 34.950 212.730 34.950 212.730 34.935 ;
        RECT 212.730 34.940 228.525 34.950 ;
        POLYGON 228.525 35.150 228.705 34.940 228.525 34.940 ;
        POLYGON 237.395 35.150 237.670 35.150 237.670 34.940 ;
        RECT 237.670 35.140 245.385 35.150 ;
        POLYGON 245.385 35.150 245.425 35.140 245.385 35.140 ;
        POLYGON 252.540 35.150 252.540 35.140 252.500 35.140 ;
        RECT 252.540 35.140 259.530 35.150 ;
        RECT 237.670 35.115 245.425 35.140 ;
        POLYGON 245.425 35.140 245.555 35.115 245.425 35.115 ;
        POLYGON 252.500 35.140 252.500 35.130 252.460 35.130 ;
        RECT 252.500 35.130 259.530 35.140 ;
        POLYGON 252.435 35.130 252.435 35.115 252.365 35.115 ;
        RECT 252.435 35.115 259.530 35.130 ;
        RECT 237.670 35.105 245.560 35.115 ;
        POLYGON 245.560 35.115 245.605 35.105 245.560 35.105 ;
        POLYGON 252.365 35.115 252.365 35.110 252.340 35.110 ;
        RECT 252.365 35.110 259.530 35.115 ;
        POLYGON 252.335 35.110 252.335 35.105 252.310 35.105 ;
        RECT 252.335 35.105 259.530 35.110 ;
        RECT 237.670 35.090 245.605 35.105 ;
        POLYGON 245.605 35.105 245.665 35.090 245.605 35.090 ;
        POLYGON 252.310 35.105 252.310 35.090 252.230 35.090 ;
        RECT 252.310 35.090 259.530 35.105 ;
        RECT 237.670 35.060 245.665 35.090 ;
        POLYGON 245.665 35.090 245.810 35.060 245.665 35.060 ;
        POLYGON 252.230 35.090 252.230 35.075 252.155 35.075 ;
        RECT 252.230 35.075 259.530 35.090 ;
        POLYGON 252.150 35.075 252.150 35.065 252.080 35.065 ;
        RECT 252.150 35.065 259.530 35.075 ;
        POLYGON 252.080 35.065 252.080 35.060 252.050 35.060 ;
        RECT 252.080 35.060 259.530 35.065 ;
        RECT 237.670 35.035 245.810 35.060 ;
        POLYGON 245.810 35.060 245.940 35.035 245.810 35.035 ;
        POLYGON 252.050 35.060 252.050 35.035 251.910 35.035 ;
        RECT 252.050 35.035 259.530 35.060 ;
        RECT 237.670 34.990 245.940 35.035 ;
        POLYGON 245.940 35.035 246.215 34.990 245.940 34.990 ;
        POLYGON 251.910 35.035 251.910 35.025 251.855 35.025 ;
        RECT 251.910 35.025 259.530 35.035 ;
        POLYGON 251.855 35.025 251.855 34.990 251.675 34.990 ;
        RECT 251.855 34.990 259.530 35.025 ;
        RECT 237.670 34.960 246.220 34.990 ;
        POLYGON 246.220 34.990 246.375 34.960 246.220 34.960 ;
        POLYGON 251.675 34.990 251.675 34.980 251.625 34.980 ;
        RECT 251.675 34.980 259.530 34.990 ;
        POLYGON 251.625 34.980 251.625 34.970 251.530 34.970 ;
        RECT 251.625 34.970 259.530 34.980 ;
        POLYGON 251.530 34.970 251.530 34.965 251.480 34.965 ;
        RECT 251.530 34.965 259.530 34.970 ;
        POLYGON 251.480 34.965 251.480 34.960 251.445 34.960 ;
        RECT 251.480 34.960 259.530 34.965 ;
        RECT 237.670 34.940 246.380 34.960 ;
        POLYGON 246.380 34.960 246.500 34.940 246.380 34.940 ;
        POLYGON 251.445 34.960 251.445 34.940 251.295 34.940 ;
        RECT 251.445 34.940 259.530 34.960 ;
        RECT 212.730 34.930 228.705 34.940 ;
        POLYGON 228.705 34.940 228.710 34.930 228.705 34.930 ;
        POLYGON 237.670 34.940 237.680 34.940 237.680 34.930 ;
        RECT 237.680 34.930 246.505 34.940 ;
        POLYGON 246.505 34.940 246.570 34.930 246.505 34.930 ;
        POLYGON 251.295 34.940 251.295 34.930 251.220 34.930 ;
        RECT 251.295 34.930 259.530 34.940 ;
        POLYGON 259.530 35.155 259.820 35.155 259.530 34.930 ;
        POLYGON 266.470 35.155 266.470 35.105 266.430 35.105 ;
        RECT 266.470 35.105 275.495 35.155 ;
        POLYGON 266.430 35.105 266.430 35.025 266.365 35.025 ;
        RECT 266.430 35.025 275.495 35.105 ;
        POLYGON 266.365 35.025 266.365 34.930 266.280 34.930 ;
        RECT 266.365 34.930 275.495 35.025 ;
        POLYGON 275.495 35.235 275.635 35.235 275.495 34.930 ;
        POLYGON 287.320 35.225 287.320 34.950 287.280 34.950 ;
        RECT 287.320 34.950 303.120 35.235 ;
        POLYGON 212.730 34.930 213.040 34.930 213.040 34.430 ;
        RECT 213.040 34.650 228.710 34.930 ;
        POLYGON 228.710 34.930 228.955 34.650 228.710 34.650 ;
        POLYGON 237.680 34.930 237.775 34.930 237.775 34.865 ;
        RECT 237.775 34.925 246.570 34.930 ;
        POLYGON 246.570 34.930 246.605 34.925 246.570 34.925 ;
        POLYGON 251.220 34.930 251.220 34.925 251.180 34.925 ;
        RECT 251.220 34.925 259.455 34.930 ;
        RECT 237.775 34.915 246.605 34.925 ;
        POLYGON 246.605 34.925 246.685 34.915 246.605 34.915 ;
        POLYGON 251.180 34.925 251.180 34.915 251.110 34.915 ;
        RECT 251.180 34.915 259.455 34.925 ;
        RECT 237.775 34.900 246.685 34.915 ;
        POLYGON 246.685 34.915 246.795 34.900 246.685 34.900 ;
        POLYGON 251.110 34.915 251.110 34.900 251.000 34.900 ;
        RECT 251.110 34.900 259.455 34.915 ;
        RECT 237.775 34.865 246.805 34.900 ;
        POLYGON 246.805 34.900 247.130 34.865 246.805 34.865 ;
        POLYGON 250.990 34.900 250.990 34.870 250.780 34.870 ;
        RECT 250.990 34.870 259.455 34.900 ;
        POLYGON 259.455 34.930 259.530 34.930 259.455 34.870 ;
        POLYGON 266.280 34.930 266.280 34.875 266.230 34.875 ;
        RECT 266.280 34.875 275.095 34.930 ;
        POLYGON 266.230 34.875 266.230 34.870 266.225 34.870 ;
        RECT 266.230 34.870 275.095 34.875 ;
        POLYGON 250.780 34.870 250.780 34.865 250.705 34.865 ;
        RECT 250.780 34.865 259.210 34.870 ;
        POLYGON 237.775 34.865 237.940 34.865 237.940 34.750 ;
        RECT 237.940 34.855 247.130 34.865 ;
        POLYGON 247.130 34.865 247.210 34.855 247.130 34.855 ;
        POLYGON 250.705 34.865 250.705 34.860 250.625 34.860 ;
        RECT 250.705 34.860 259.210 34.865 ;
        POLYGON 250.620 34.860 250.620 34.855 250.570 34.855 ;
        RECT 250.620 34.855 259.210 34.860 ;
        RECT 237.940 34.830 247.210 34.855 ;
        POLYGON 247.210 34.855 247.415 34.830 247.210 34.830 ;
        POLYGON 250.570 34.855 250.570 34.835 250.365 34.835 ;
        RECT 250.570 34.835 259.210 34.855 ;
        POLYGON 250.360 34.835 250.360 34.830 250.300 34.830 ;
        RECT 250.360 34.830 259.210 34.835 ;
        RECT 237.940 34.825 247.415 34.830 ;
        POLYGON 247.415 34.830 247.485 34.825 247.415 34.825 ;
        POLYGON 250.300 34.830 250.300 34.825 250.235 34.825 ;
        RECT 250.300 34.825 259.210 34.830 ;
        RECT 237.940 34.810 247.485 34.825 ;
        POLYGON 247.485 34.825 247.760 34.810 247.485 34.810 ;
        POLYGON 250.235 34.825 250.235 34.810 250.055 34.810 ;
        RECT 250.235 34.810 259.210 34.825 ;
        RECT 237.940 34.790 247.760 34.810 ;
        POLYGON 247.760 34.810 248.050 34.790 247.760 34.790 ;
        POLYGON 250.055 34.810 250.055 34.800 249.930 34.800 ;
        RECT 250.055 34.800 259.210 34.810 ;
        POLYGON 249.920 34.800 249.920 34.795 249.860 34.795 ;
        RECT 249.920 34.795 259.210 34.800 ;
        POLYGON 249.850 34.795 249.850 34.790 249.690 34.790 ;
        RECT 249.850 34.790 259.210 34.795 ;
        RECT 237.940 34.780 248.055 34.790 ;
        POLYGON 248.055 34.790 248.245 34.780 248.055 34.780 ;
        POLYGON 249.685 34.790 249.685 34.780 249.385 34.780 ;
        RECT 249.685 34.780 259.210 34.790 ;
        RECT 237.940 34.770 248.315 34.780 ;
        POLYGON 248.315 34.780 248.835 34.770 248.315 34.770 ;
        POLYGON 249.385 34.780 249.385 34.770 249.085 34.770 ;
        RECT 249.385 34.770 259.210 34.780 ;
        RECT 237.940 34.750 259.210 34.770 ;
        POLYGON 237.940 34.750 238.080 34.750 238.080 34.650 ;
        RECT 238.080 34.685 259.210 34.750 ;
        POLYGON 259.210 34.870 259.455 34.870 259.210 34.685 ;
        POLYGON 266.225 34.870 266.225 34.700 266.075 34.700 ;
        RECT 266.225 34.700 275.095 34.870 ;
        POLYGON 266.075 34.700 266.075 34.685 266.060 34.685 ;
        RECT 266.075 34.685 275.095 34.700 ;
        RECT 238.080 34.650 258.750 34.685 ;
        RECT 213.040 34.430 228.955 34.650 ;
        POLYGON 213.040 34.430 213.125 34.430 213.125 34.300 ;
        RECT 213.125 34.400 228.955 34.430 ;
        POLYGON 228.955 34.650 229.190 34.400 228.955 34.400 ;
        POLYGON 238.080 34.650 238.320 34.650 238.320 34.480 ;
        RECT 238.320 34.480 258.750 34.650 ;
        POLYGON 238.320 34.480 238.440 34.480 238.440 34.400 ;
        RECT 238.440 34.400 258.750 34.480 ;
        RECT 213.125 34.380 229.190 34.400 ;
        POLYGON 229.190 34.400 229.205 34.380 229.190 34.380 ;
        POLYGON 238.440 34.400 238.475 34.400 238.475 34.380 ;
        RECT 238.475 34.380 258.750 34.400 ;
        RECT 213.125 34.330 229.205 34.380 ;
        POLYGON 229.205 34.380 229.250 34.330 229.205 34.330 ;
        POLYGON 238.475 34.380 238.550 34.380 238.550 34.330 ;
        RECT 238.550 34.355 258.750 34.380 ;
        POLYGON 258.750 34.685 259.210 34.685 258.750 34.355 ;
        POLYGON 266.060 34.685 266.060 34.555 265.950 34.555 ;
        RECT 266.060 34.555 275.095 34.685 ;
        POLYGON 265.950 34.555 265.950 34.445 265.850 34.445 ;
        RECT 265.950 34.445 275.095 34.555 ;
        POLYGON 265.850 34.445 265.850 34.355 265.775 34.355 ;
        RECT 265.850 34.355 275.095 34.445 ;
        RECT 238.550 34.330 258.660 34.355 ;
        RECT 213.125 34.300 229.250 34.330 ;
        POLYGON 213.125 34.300 213.790 34.300 213.790 33.285 ;
        RECT 213.790 34.270 229.250 34.300 ;
        POLYGON 229.250 34.330 229.305 34.270 229.250 34.270 ;
        POLYGON 238.550 34.330 238.645 34.330 238.645 34.270 ;
        RECT 238.645 34.300 258.660 34.330 ;
        POLYGON 258.660 34.355 258.750 34.355 258.660 34.300 ;
        POLYGON 265.775 34.355 265.775 34.300 265.725 34.300 ;
        RECT 265.775 34.300 275.095 34.355 ;
        RECT 238.645 34.270 258.300 34.300 ;
        RECT 213.790 34.080 229.305 34.270 ;
        POLYGON 229.305 34.270 229.485 34.080 229.305 34.080 ;
        POLYGON 238.645 34.270 238.710 34.270 238.710 34.230 ;
        RECT 238.710 34.230 258.300 34.270 ;
        POLYGON 238.710 34.230 238.935 34.230 238.935 34.080 ;
        RECT 238.935 34.080 258.300 34.230 ;
        RECT 213.790 34.005 229.485 34.080 ;
        POLYGON 229.485 34.080 229.550 34.005 229.485 34.005 ;
        POLYGON 238.935 34.080 238.965 34.080 238.965 34.060 ;
        RECT 238.965 34.060 258.300 34.080 ;
        POLYGON 258.300 34.300 258.660 34.300 258.300 34.060 ;
        POLYGON 265.725 34.300 265.725 34.275 265.705 34.275 ;
        RECT 265.725 34.275 275.095 34.300 ;
        POLYGON 265.705 34.275 265.705 34.060 265.515 34.060 ;
        RECT 265.705 34.060 275.095 34.275 ;
        POLYGON 275.095 34.930 275.495 34.930 275.095 34.060 ;
        POLYGON 287.280 34.930 287.280 34.060 287.160 34.060 ;
        RECT 287.280 34.060 303.120 34.950 ;
        POLYGON 238.965 34.060 239.055 34.060 239.055 34.005 ;
        RECT 239.055 34.005 257.850 34.060 ;
        RECT 213.790 33.790 229.550 34.005 ;
        POLYGON 229.550 34.005 229.765 33.790 229.550 33.790 ;
        POLYGON 239.055 34.005 239.300 34.005 239.300 33.865 ;
        RECT 239.300 33.865 257.850 34.005 ;
        POLYGON 239.300 33.865 239.430 33.865 239.430 33.790 ;
        RECT 239.430 33.790 257.850 33.865 ;
        POLYGON 257.850 34.060 258.295 34.060 257.850 33.790 ;
        POLYGON 265.515 34.060 265.515 34.030 265.490 34.030 ;
        RECT 265.515 34.030 274.500 34.060 ;
        POLYGON 265.490 34.030 265.490 33.990 265.450 33.990 ;
        RECT 265.490 33.990 274.500 34.030 ;
        POLYGON 265.450 33.990 265.450 33.790 265.265 33.790 ;
        RECT 265.450 33.790 274.500 33.990 ;
        RECT 213.790 33.640 229.765 33.790 ;
        POLYGON 229.765 33.790 229.910 33.640 229.765 33.640 ;
        POLYGON 239.430 33.790 239.615 33.790 239.615 33.685 ;
        RECT 239.615 33.685 257.495 33.790 ;
        POLYGON 239.615 33.685 239.670 33.685 239.670 33.655 ;
        RECT 239.670 33.655 257.495 33.685 ;
        POLYGON 239.670 33.655 239.695 33.655 239.695 33.640 ;
        RECT 239.695 33.640 257.495 33.655 ;
        RECT 213.790 33.385 229.910 33.640 ;
        POLYGON 229.910 33.640 230.165 33.385 229.910 33.385 ;
        POLYGON 239.695 33.640 240.195 33.640 240.195 33.385 ;
        RECT 240.195 33.605 257.495 33.640 ;
        POLYGON 257.495 33.790 257.850 33.790 257.495 33.605 ;
        POLYGON 265.265 33.790 265.265 33.780 265.255 33.780 ;
        RECT 265.265 33.780 274.500 33.790 ;
        POLYGON 265.255 33.780 265.255 33.605 265.085 33.605 ;
        RECT 265.255 33.605 274.500 33.780 ;
        RECT 240.195 33.560 257.415 33.605 ;
        POLYGON 257.415 33.605 257.495 33.605 257.415 33.560 ;
        POLYGON 265.085 33.605 265.085 33.560 265.040 33.560 ;
        RECT 265.085 33.560 274.500 33.605 ;
        RECT 240.195 33.415 257.115 33.560 ;
        POLYGON 257.115 33.560 257.415 33.560 257.115 33.415 ;
        POLYGON 265.040 33.560 265.040 33.515 264.995 33.515 ;
        RECT 265.040 33.515 274.500 33.560 ;
        POLYGON 264.995 33.515 264.995 33.415 264.900 33.415 ;
        RECT 264.995 33.415 274.500 33.515 ;
        RECT 240.195 33.385 256.360 33.415 ;
        RECT 213.790 33.285 230.165 33.385 ;
        POLYGON 213.790 33.285 214.030 33.285 214.030 32.950 ;
        RECT 214.030 33.270 230.165 33.285 ;
        POLYGON 230.165 33.385 230.285 33.270 230.165 33.270 ;
        POLYGON 240.195 33.385 240.255 33.385 240.255 33.355 ;
        RECT 240.255 33.355 256.360 33.385 ;
        POLYGON 240.255 33.355 240.440 33.355 240.440 33.270 ;
        RECT 240.440 33.270 256.360 33.355 ;
        RECT 214.030 33.235 230.285 33.270 ;
        POLYGON 230.285 33.270 230.320 33.235 230.285 33.235 ;
        POLYGON 240.440 33.270 240.515 33.270 240.515 33.235 ;
        RECT 240.515 33.235 256.360 33.270 ;
        RECT 214.030 33.060 230.320 33.235 ;
        POLYGON 230.320 33.235 230.505 33.060 230.320 33.060 ;
        POLYGON 240.515 33.235 240.660 33.235 240.660 33.170 ;
        RECT 240.660 33.170 256.360 33.235 ;
        POLYGON 240.660 33.170 240.745 33.170 240.745 33.135 ;
        RECT 240.745 33.135 256.360 33.170 ;
        POLYGON 240.745 33.135 240.905 33.135 240.905 33.060 ;
        RECT 240.905 33.060 256.360 33.135 ;
        POLYGON 256.360 33.415 257.115 33.415 256.360 33.060 ;
        POLYGON 264.900 33.415 264.900 33.360 264.850 33.360 ;
        RECT 264.900 33.360 274.500 33.415 ;
        POLYGON 264.850 33.360 264.850 33.225 264.720 33.225 ;
        RECT 264.850 33.225 274.500 33.360 ;
        POLYGON 264.720 33.225 264.720 33.060 264.560 33.060 ;
        RECT 264.720 33.060 274.500 33.225 ;
        RECT 214.030 33.020 230.505 33.060 ;
        POLYGON 230.505 33.060 230.545 33.020 230.505 33.020 ;
        POLYGON 240.905 33.060 240.995 33.060 240.995 33.020 ;
        RECT 240.995 33.045 256.330 33.060 ;
        POLYGON 256.330 33.060 256.360 33.060 256.330 33.045 ;
        POLYGON 264.560 33.060 264.560 33.045 264.545 33.045 ;
        RECT 264.560 33.045 274.500 33.060 ;
        RECT 240.995 33.020 255.905 33.045 ;
        RECT 214.030 32.950 230.545 33.020 ;
        POLYGON 214.030 32.950 214.200 32.950 214.200 32.705 ;
        RECT 214.200 32.835 230.545 32.950 ;
        POLYGON 230.545 33.020 230.745 32.835 230.545 32.835 ;
        POLYGON 240.995 33.020 241.315 33.020 241.315 32.875 ;
        RECT 241.315 32.875 255.905 33.020 ;
        POLYGON 255.905 33.045 256.330 33.045 255.905 32.875 ;
        POLYGON 264.545 33.045 264.545 32.915 264.420 32.915 ;
        RECT 264.545 32.915 274.500 33.045 ;
        POLYGON 264.420 32.915 264.420 32.875 264.385 32.875 ;
        RECT 264.420 32.905 274.500 32.915 ;
        POLYGON 274.500 34.060 275.095 34.060 274.500 32.905 ;
        POLYGON 287.160 34.055 287.160 32.905 287.000 32.905 ;
        RECT 287.160 32.905 303.120 34.060 ;
        RECT 264.420 32.875 274.380 32.905 ;
        POLYGON 241.315 32.875 241.420 32.875 241.420 32.835 ;
        RECT 241.420 32.835 255.485 32.875 ;
        RECT 214.200 32.785 230.745 32.835 ;
        POLYGON 230.745 32.835 230.795 32.785 230.745 32.785 ;
        POLYGON 241.420 32.835 241.555 32.835 241.555 32.785 ;
        RECT 241.555 32.785 255.485 32.835 ;
        RECT 214.200 32.700 230.795 32.785 ;
        POLYGON 230.795 32.785 230.890 32.700 230.795 32.700 ;
        POLYGON 241.555 32.785 241.680 32.785 241.680 32.740 ;
        RECT 241.680 32.740 255.485 32.785 ;
        POLYGON 241.680 32.740 241.780 32.740 241.780 32.700 ;
        RECT 241.780 32.700 255.485 32.740 ;
        POLYGON 255.485 32.875 255.905 32.875 255.485 32.700 ;
        POLYGON 264.385 32.875 264.385 32.865 264.375 32.865 ;
        RECT 264.385 32.865 274.380 32.875 ;
        POLYGON 264.375 32.865 264.375 32.850 264.355 32.850 ;
        RECT 264.375 32.850 274.380 32.865 ;
        POLYGON 264.355 32.850 264.355 32.700 264.200 32.700 ;
        RECT 264.355 32.700 274.380 32.850 ;
        POLYGON 274.380 32.905 274.500 32.905 274.380 32.700 ;
        POLYGON 287.000 32.890 287.000 32.710 286.975 32.710 ;
        RECT 287.000 32.710 303.120 32.905 ;
        RECT 179.410 32.365 196.580 32.700 ;
        RECT 159.640 32.320 168.445 32.365 ;
        RECT 63.450 32.240 157.300 32.320 ;
        POLYGON 157.300 32.320 157.350 32.240 157.300 32.240 ;
        POLYGON 159.470 32.320 159.470 32.240 159.235 32.240 ;
        RECT 159.470 32.240 168.445 32.320 ;
        RECT 63.450 32.210 157.350 32.240 ;
        POLYGON 157.350 32.240 157.370 32.210 157.350 32.210 ;
        POLYGON 159.235 32.240 159.235 32.210 159.145 32.210 ;
        RECT 159.235 32.210 168.445 32.240 ;
        RECT 63.450 32.205 157.370 32.210 ;
        POLYGON 157.370 32.210 157.375 32.205 157.370 32.205 ;
        POLYGON 159.145 32.210 159.145 32.205 159.120 32.205 ;
        RECT 159.145 32.205 168.445 32.210 ;
        RECT 63.450 32.165 157.375 32.205 ;
        POLYGON 157.375 32.205 157.400 32.165 157.375 32.165 ;
        POLYGON 159.120 32.205 159.120 32.165 158.980 32.165 ;
        RECT 159.120 32.165 168.445 32.205 ;
        RECT 63.450 32.100 157.400 32.165 ;
        POLYGON 157.400 32.165 157.445 32.100 157.400 32.100 ;
        POLYGON 158.980 32.165 158.980 32.100 158.755 32.100 ;
        RECT 158.980 32.100 168.445 32.165 ;
        RECT 63.450 32.075 157.445 32.100 ;
        POLYGON 158.755 32.100 158.755 32.095 158.740 32.095 ;
        RECT 158.755 32.095 168.445 32.100 ;
        POLYGON 157.445 32.095 157.460 32.075 157.445 32.075 ;
        POLYGON 158.740 32.095 158.740 32.075 158.675 32.075 ;
        RECT 158.740 32.075 168.445 32.095 ;
        RECT 63.450 32.040 157.460 32.075 ;
        POLYGON 157.460 32.075 157.485 32.040 157.460 32.040 ;
        RECT 63.450 32.015 157.485 32.040 ;
        POLYGON 158.675 32.075 158.675 32.035 158.545 32.035 ;
        RECT 158.675 32.035 168.445 32.075 ;
        POLYGON 157.485 32.035 157.500 32.015 157.485 32.015 ;
        POLYGON 158.545 32.035 158.545 32.015 158.475 32.015 ;
        RECT 158.545 32.015 168.445 32.035 ;
        RECT 63.450 32.005 157.500 32.015 ;
        POLYGON 157.500 32.015 157.505 32.005 157.500 32.005 ;
        POLYGON 158.475 32.015 158.475 32.005 158.430 32.005 ;
        RECT 158.475 32.005 168.445 32.015 ;
        RECT 63.450 31.970 157.505 32.005 ;
        POLYGON 157.505 32.005 157.530 31.970 157.505 31.970 ;
        POLYGON 158.430 32.005 158.430 31.970 158.290 31.970 ;
        RECT 158.430 31.970 168.445 32.005 ;
        RECT 63.450 31.910 157.530 31.970 ;
        POLYGON 157.530 31.970 157.570 31.910 157.530 31.910 ;
        POLYGON 158.290 31.970 158.290 31.940 158.165 31.940 ;
        RECT 158.290 31.950 168.445 31.970 ;
        POLYGON 168.445 32.365 168.875 32.365 168.445 31.950 ;
        POLYGON 179.210 32.360 179.210 32.345 179.200 32.345 ;
        RECT 179.210 32.345 196.580 32.365 ;
        POLYGON 179.200 32.345 179.200 32.190 179.105 32.190 ;
        RECT 179.200 32.190 196.580 32.345 ;
        POLYGON 179.105 32.190 179.105 31.950 178.965 31.950 ;
        RECT 179.105 31.950 196.580 32.190 ;
        RECT 158.290 31.940 168.255 31.950 ;
        RECT 63.450 31.855 157.570 31.910 ;
        POLYGON 158.165 31.940 158.165 31.905 158.025 31.905 ;
        RECT 158.165 31.905 168.255 31.940 ;
        POLYGON 157.570 31.905 157.605 31.855 157.570 31.855 ;
        POLYGON 158.020 31.905 158.020 31.855 157.825 31.855 ;
        RECT 158.020 31.855 168.255 31.905 ;
        RECT 63.450 31.835 157.605 31.855 ;
        POLYGON 157.605 31.855 157.620 31.835 157.605 31.835 ;
        POLYGON 157.825 31.855 157.825 31.835 157.735 31.835 ;
        RECT 157.825 31.835 168.255 31.855 ;
        RECT 63.450 31.820 157.620 31.835 ;
        POLYGON 157.735 31.835 157.735 31.830 157.710 31.830 ;
        RECT 157.735 31.830 168.255 31.835 ;
        POLYGON 157.620 31.830 157.630 31.820 157.620 31.820 ;
        POLYGON 157.705 31.830 157.705 31.820 157.665 31.820 ;
        RECT 157.705 31.820 168.255 31.830 ;
        RECT 63.450 31.815 157.630 31.820 ;
        POLYGON 157.665 31.820 157.665 31.815 157.640 31.815 ;
        RECT 157.665 31.815 168.255 31.820 ;
        RECT 63.450 31.770 168.255 31.815 ;
        POLYGON 168.255 31.950 168.445 31.950 168.255 31.770 ;
        POLYGON 178.965 31.950 178.965 31.770 178.860 31.770 ;
        RECT 178.965 31.770 196.580 31.950 ;
        RECT 63.450 30.785 167.135 31.770 ;
        POLYGON 167.135 31.770 168.255 31.770 167.135 30.785 ;
        POLYGON 178.860 31.765 178.860 31.750 178.850 31.750 ;
        RECT 178.860 31.750 196.580 31.770 ;
        POLYGON 178.850 31.750 178.850 31.455 178.660 31.455 ;
        RECT 178.850 31.455 196.580 31.750 ;
        POLYGON 178.660 31.455 178.660 30.785 178.230 30.785 ;
        RECT 178.660 30.785 196.580 31.455 ;
        RECT 63.450 30.670 166.995 30.785 ;
        POLYGON 166.995 30.785 167.135 30.785 166.995 30.670 ;
        POLYGON 178.230 30.785 178.230 30.670 178.155 30.670 ;
        RECT 178.230 30.670 196.580 30.785 ;
        RECT 63.450 30.405 166.620 30.670 ;
        POLYGON 63.450 30.405 64.025 30.405 64.025 29.560 ;
        RECT 64.025 30.365 166.620 30.405 ;
        POLYGON 166.620 30.670 166.995 30.670 166.620 30.365 ;
        POLYGON 178.155 30.670 178.155 30.630 178.130 30.630 ;
        RECT 178.155 30.630 196.580 30.670 ;
        POLYGON 178.130 30.630 178.130 30.375 177.945 30.375 ;
        RECT 178.130 30.475 196.580 30.630 ;
        POLYGON 196.580 32.700 197.100 32.700 196.580 30.475 ;
        POLYGON 214.200 32.700 214.575 32.700 214.575 32.170 ;
        RECT 214.575 32.600 230.890 32.700 ;
        POLYGON 230.890 32.700 231.005 32.600 230.890 32.600 ;
        POLYGON 241.780 32.700 242.040 32.700 242.040 32.600 ;
        RECT 242.040 32.620 255.295 32.700 ;
        POLYGON 255.295 32.700 255.485 32.700 255.295 32.620 ;
        POLYGON 264.200 32.700 264.200 32.620 264.120 32.620 ;
        RECT 264.200 32.620 274.070 32.700 ;
        RECT 242.040 32.600 255.160 32.620 ;
        RECT 214.575 32.550 231.005 32.600 ;
        POLYGON 231.005 32.600 231.060 32.550 231.005 32.550 ;
        POLYGON 242.040 32.600 242.165 32.600 242.165 32.550 ;
        RECT 242.165 32.575 255.160 32.600 ;
        POLYGON 255.160 32.620 255.295 32.620 255.160 32.575 ;
        POLYGON 264.120 32.620 264.120 32.575 264.075 32.575 ;
        RECT 264.120 32.575 274.070 32.620 ;
        RECT 242.165 32.550 254.670 32.575 ;
        RECT 214.575 32.475 231.060 32.550 ;
        POLYGON 231.060 32.550 231.140 32.475 231.060 32.475 ;
        POLYGON 242.165 32.550 242.310 32.550 242.310 32.495 ;
        RECT 242.310 32.495 254.670 32.550 ;
        POLYGON 242.310 32.495 242.360 32.495 242.360 32.475 ;
        RECT 242.360 32.475 254.670 32.495 ;
        RECT 214.575 32.350 231.140 32.475 ;
        POLYGON 231.140 32.475 231.280 32.350 231.140 32.350 ;
        POLYGON 242.360 32.475 242.385 32.475 242.385 32.465 ;
        RECT 242.385 32.465 254.670 32.475 ;
        POLYGON 242.385 32.465 242.720 32.465 242.720 32.360 ;
        RECT 242.720 32.405 254.670 32.465 ;
        POLYGON 254.670 32.575 255.160 32.575 254.670 32.405 ;
        POLYGON 264.075 32.575 264.075 32.405 263.895 32.405 ;
        RECT 264.075 32.405 274.070 32.575 ;
        RECT 242.720 32.360 254.225 32.405 ;
        POLYGON 242.720 32.360 242.750 32.360 242.750 32.350 ;
        RECT 242.750 32.350 254.225 32.360 ;
        RECT 214.575 32.295 231.280 32.350 ;
        POLYGON 231.280 32.350 231.345 32.295 231.280 32.295 ;
        POLYGON 242.750 32.350 242.915 32.350 242.915 32.295 ;
        RECT 242.915 32.295 254.225 32.350 ;
        RECT 214.575 32.205 231.350 32.295 ;
        POLYGON 231.350 32.295 231.445 32.205 231.350 32.205 ;
        POLYGON 242.915 32.295 243.190 32.295 243.190 32.205 ;
        RECT 243.190 32.250 254.225 32.295 ;
        POLYGON 254.225 32.405 254.670 32.405 254.225 32.250 ;
        POLYGON 263.895 32.405 263.895 32.335 263.820 32.335 ;
        RECT 263.895 32.335 274.070 32.405 ;
        POLYGON 263.820 32.330 263.820 32.250 263.735 32.250 ;
        RECT 263.820 32.250 274.070 32.335 ;
        RECT 243.190 32.205 253.990 32.250 ;
        RECT 214.575 32.165 231.445 32.205 ;
        POLYGON 231.445 32.205 231.490 32.165 231.445 32.165 ;
        POLYGON 243.190 32.205 243.315 32.205 243.315 32.165 ;
        RECT 243.315 32.185 253.990 32.205 ;
        POLYGON 253.990 32.250 254.225 32.250 253.990 32.185 ;
        POLYGON 263.735 32.250 263.735 32.185 263.665 32.185 ;
        RECT 263.735 32.185 274.070 32.250 ;
        RECT 243.315 32.165 253.915 32.185 ;
        POLYGON 253.915 32.185 253.985 32.185 253.915 32.165 ;
        POLYGON 263.665 32.185 263.665 32.165 263.645 32.165 ;
        RECT 263.665 32.165 274.070 32.185 ;
        POLYGON 274.070 32.700 274.380 32.700 274.070 32.165 ;
        POLYGON 286.975 32.700 286.975 32.165 286.900 32.165 ;
        RECT 286.975 32.165 303.120 32.710 ;
        POLYGON 214.575 32.165 214.980 32.165 214.980 31.630 ;
        RECT 214.980 32.095 231.490 32.165 ;
        POLYGON 231.490 32.165 231.580 32.095 231.490 32.095 ;
        POLYGON 243.315 32.165 243.455 32.165 243.455 32.120 ;
        RECT 243.455 32.120 253.410 32.165 ;
        POLYGON 243.455 32.120 243.545 32.120 243.545 32.095 ;
        RECT 243.545 32.095 253.410 32.120 ;
        RECT 214.980 32.005 231.580 32.095 ;
        POLYGON 231.580 32.095 231.685 32.005 231.580 32.005 ;
        POLYGON 243.545 32.095 243.775 32.095 243.775 32.035 ;
        RECT 243.775 32.035 253.410 32.095 ;
        POLYGON 243.780 32.035 243.900 32.035 243.900 32.005 ;
        RECT 243.900 32.020 253.410 32.035 ;
        POLYGON 253.410 32.165 253.915 32.165 253.410 32.020 ;
        POLYGON 263.645 32.165 263.645 32.025 263.495 32.025 ;
        RECT 263.645 32.025 273.840 32.165 ;
        POLYGON 263.495 32.025 263.495 32.020 263.490 32.020 ;
        RECT 263.495 32.020 273.840 32.025 ;
        RECT 243.900 32.005 253.155 32.020 ;
        RECT 214.980 31.830 231.685 32.005 ;
        POLYGON 231.685 32.005 231.900 31.830 231.685 31.830 ;
        POLYGON 243.900 32.005 244.040 32.005 244.040 31.970 ;
        RECT 244.040 31.970 253.155 32.005 ;
        POLYGON 244.040 31.970 244.530 31.970 244.530 31.840 ;
        RECT 244.530 31.945 253.155 31.970 ;
        POLYGON 253.155 32.020 253.405 32.020 253.155 31.945 ;
        POLYGON 263.490 32.020 263.490 31.945 263.410 31.945 ;
        RECT 263.490 31.945 273.840 32.020 ;
        RECT 244.530 31.870 252.820 31.945 ;
        POLYGON 252.820 31.945 253.155 31.945 252.820 31.870 ;
        POLYGON 263.410 31.945 263.410 31.870 263.335 31.870 ;
        RECT 263.410 31.870 273.840 31.945 ;
        RECT 244.530 31.840 252.120 31.870 ;
        POLYGON 244.530 31.840 244.580 31.840 244.580 31.830 ;
        RECT 244.580 31.830 252.120 31.840 ;
        RECT 214.980 31.685 231.900 31.830 ;
        POLYGON 231.900 31.830 232.075 31.685 231.900 31.685 ;
        POLYGON 244.580 31.830 244.860 31.830 244.860 31.775 ;
        RECT 244.860 31.775 252.120 31.830 ;
        POLYGON 244.860 31.775 245.305 31.775 245.305 31.685 ;
        RECT 245.305 31.715 252.120 31.775 ;
        POLYGON 252.120 31.870 252.820 31.870 252.120 31.715 ;
        POLYGON 263.335 31.870 263.335 31.790 263.250 31.790 ;
        RECT 263.335 31.790 273.840 31.870 ;
        POLYGON 263.250 31.790 263.250 31.780 263.240 31.780 ;
        RECT 263.250 31.780 273.840 31.790 ;
        POLYGON 263.240 31.780 263.240 31.715 263.165 31.715 ;
        RECT 263.240 31.770 273.840 31.780 ;
        POLYGON 273.840 32.165 274.070 32.165 273.840 31.770 ;
        POLYGON 286.900 32.165 286.900 31.770 286.845 31.770 ;
        RECT 286.900 31.770 303.120 32.165 ;
        RECT 263.240 31.715 273.535 31.770 ;
        RECT 245.305 31.705 252.080 31.715 ;
        POLYGON 252.080 31.715 252.120 31.715 252.080 31.705 ;
        POLYGON 263.165 31.715 263.165 31.705 263.155 31.705 ;
        RECT 263.165 31.705 273.535 31.715 ;
        RECT 245.305 31.685 251.655 31.705 ;
        RECT 214.980 31.650 232.075 31.685 ;
        POLYGON 232.075 31.685 232.115 31.650 232.075 31.650 ;
        POLYGON 245.305 31.685 245.480 31.685 245.480 31.650 ;
        RECT 245.480 31.650 251.655 31.685 ;
        RECT 214.980 31.630 232.115 31.650 ;
        POLYGON 214.980 31.630 215.390 31.630 215.390 31.080 ;
        RECT 215.390 31.555 232.115 31.630 ;
        POLYGON 232.115 31.650 232.240 31.555 232.115 31.555 ;
        POLYGON 245.480 31.650 245.605 31.650 245.605 31.625 ;
        RECT 245.605 31.635 251.655 31.650 ;
        POLYGON 251.655 31.705 252.080 31.705 251.655 31.635 ;
        POLYGON 263.155 31.705 263.155 31.695 263.145 31.695 ;
        RECT 263.155 31.695 273.535 31.705 ;
        POLYGON 263.145 31.695 263.145 31.635 263.075 31.635 ;
        RECT 263.145 31.635 273.535 31.695 ;
        RECT 245.605 31.625 251.105 31.635 ;
        POLYGON 245.605 31.625 245.955 31.625 245.955 31.575 ;
        RECT 245.955 31.575 251.105 31.625 ;
        POLYGON 245.960 31.575 246.105 31.575 246.105 31.555 ;
        RECT 246.105 31.555 251.105 31.575 ;
        RECT 215.390 31.435 232.240 31.555 ;
        POLYGON 232.240 31.555 232.390 31.435 232.240 31.435 ;
        POLYGON 246.105 31.555 246.585 31.555 246.585 31.490 ;
        RECT 246.585 31.545 251.105 31.555 ;
        POLYGON 251.105 31.635 251.655 31.635 251.105 31.545 ;
        POLYGON 263.075 31.635 263.075 31.545 262.975 31.545 ;
        RECT 263.075 31.545 273.535 31.635 ;
        RECT 246.585 31.530 251.000 31.545 ;
        POLYGON 251.000 31.545 251.105 31.545 251.000 31.530 ;
        POLYGON 262.975 31.545 262.975 31.530 262.960 31.530 ;
        RECT 262.975 31.530 273.535 31.545 ;
        RECT 246.585 31.490 250.495 31.530 ;
        POLYGON 246.585 31.490 246.685 31.490 246.685 31.475 ;
        RECT 246.685 31.475 250.495 31.490 ;
        POLYGON 250.495 31.530 251.000 31.530 250.495 31.475 ;
        POLYGON 262.960 31.530 262.960 31.475 262.895 31.475 ;
        RECT 262.960 31.475 273.535 31.530 ;
        POLYGON 246.685 31.475 247.065 31.475 247.065 31.445 ;
        RECT 247.065 31.445 250.195 31.475 ;
        POLYGON 250.195 31.475 250.495 31.475 250.195 31.445 ;
        POLYGON 262.895 31.475 262.895 31.445 262.860 31.445 ;
        RECT 262.895 31.445 273.535 31.475 ;
        POLYGON 247.075 31.445 247.195 31.445 247.195 31.435 ;
        RECT 247.195 31.435 249.920 31.445 ;
        RECT 215.390 31.350 232.390 31.435 ;
        POLYGON 232.390 31.435 232.500 31.350 232.390 31.350 ;
        POLYGON 247.195 31.435 247.760 31.435 247.760 31.390 ;
        RECT 247.760 31.415 249.920 31.435 ;
        POLYGON 249.920 31.445 250.195 31.445 249.920 31.415 ;
        POLYGON 262.860 31.445 262.860 31.415 262.825 31.415 ;
        RECT 262.860 31.415 273.535 31.445 ;
        RECT 247.760 31.395 249.345 31.415 ;
        POLYGON 249.345 31.415 249.920 31.415 249.345 31.395 ;
        POLYGON 262.825 31.415 262.825 31.395 262.805 31.395 ;
        RECT 262.825 31.395 273.535 31.415 ;
        RECT 247.760 31.390 248.840 31.395 ;
        POLYGON 247.760 31.390 248.160 31.390 248.160 31.385 ;
        RECT 248.160 31.385 248.840 31.390 ;
        POLYGON 248.205 31.385 248.445 31.385 248.445 31.380 ;
        RECT 248.445 31.380 248.840 31.385 ;
        POLYGON 248.495 31.380 248.840 31.380 248.840 31.370 ;
        POLYGON 248.840 31.395 249.345 31.395 248.840 31.370 ;
        POLYGON 262.805 31.395 262.805 31.370 262.775 31.370 ;
        RECT 262.805 31.370 273.535 31.395 ;
        POLYGON 262.775 31.370 262.775 31.350 262.755 31.350 ;
        RECT 262.775 31.350 273.535 31.370 ;
        RECT 215.390 31.115 232.500 31.350 ;
        POLYGON 232.500 31.350 232.805 31.115 232.500 31.115 ;
        POLYGON 262.755 31.350 262.755 31.115 262.485 31.115 ;
        RECT 262.755 31.300 273.535 31.350 ;
        POLYGON 273.535 31.770 273.840 31.770 273.535 31.300 ;
        POLYGON 286.845 31.770 286.845 31.300 286.780 31.300 ;
        RECT 286.845 31.300 303.120 31.770 ;
        RECT 262.755 31.115 273.120 31.300 ;
        RECT 215.390 31.080 232.805 31.115 ;
        POLYGON 215.390 31.080 215.875 31.080 215.875 30.475 ;
        RECT 215.875 31.040 232.805 31.080 ;
        POLYGON 232.805 31.115 232.910 31.040 232.805 31.040 ;
        POLYGON 262.485 31.115 262.485 31.040 262.400 31.040 ;
        RECT 262.485 31.040 273.120 31.115 ;
        RECT 215.875 30.995 232.910 31.040 ;
        POLYGON 232.910 31.040 232.970 30.995 232.910 30.995 ;
        POLYGON 262.400 31.040 262.400 30.995 262.350 30.995 ;
        RECT 262.400 30.995 273.120 31.040 ;
        RECT 215.875 30.630 232.970 30.995 ;
        POLYGON 232.970 30.995 233.475 30.630 232.970 30.630 ;
        POLYGON 262.350 30.995 262.350 30.805 262.135 30.805 ;
        RECT 262.350 30.805 273.120 30.995 ;
        POLYGON 262.135 30.805 262.135 30.790 262.115 30.790 ;
        RECT 262.135 30.790 273.120 30.805 ;
        POLYGON 262.115 30.790 262.115 30.660 261.955 30.660 ;
        RECT 262.115 30.660 273.120 30.790 ;
        POLYGON 261.950 30.660 261.950 30.630 261.915 30.630 ;
        RECT 261.950 30.655 273.120 30.660 ;
        POLYGON 273.120 31.300 273.535 31.300 273.120 30.655 ;
        POLYGON 286.780 31.300 286.780 30.655 286.690 30.655 ;
        RECT 286.780 30.655 303.120 31.300 ;
        RECT 261.950 30.630 272.985 30.655 ;
        RECT 215.875 30.605 233.475 30.630 ;
        POLYGON 233.475 30.630 233.505 30.605 233.475 30.605 ;
        POLYGON 261.915 30.630 261.915 30.605 261.885 30.605 ;
        RECT 261.915 30.605 272.985 30.630 ;
        RECT 215.875 30.530 233.505 30.605 ;
        POLYGON 233.505 30.605 233.620 30.530 233.505 30.530 ;
        POLYGON 261.885 30.605 261.885 30.530 261.795 30.530 ;
        RECT 261.885 30.530 272.985 30.605 ;
        RECT 215.875 30.475 233.620 30.530 ;
        RECT 178.130 30.375 195.955 30.475 ;
        POLYGON 177.945 30.375 177.945 30.370 177.940 30.370 ;
        RECT 177.945 30.370 195.955 30.375 ;
        RECT 64.025 30.345 166.595 30.365 ;
        POLYGON 166.595 30.365 166.620 30.365 166.595 30.345 ;
        POLYGON 177.940 30.365 177.940 30.345 177.925 30.345 ;
        RECT 177.940 30.345 195.955 30.370 ;
        RECT 64.025 29.950 166.070 30.345 ;
        POLYGON 166.070 30.345 166.595 30.345 166.070 29.950 ;
        POLYGON 177.925 30.345 177.925 30.220 177.840 30.220 ;
        RECT 177.925 30.220 195.955 30.345 ;
        POLYGON 177.840 30.220 177.840 29.950 177.650 29.950 ;
        RECT 177.840 29.950 195.955 30.220 ;
        RECT 64.025 29.600 165.575 29.950 ;
        POLYGON 165.575 29.950 166.070 29.950 165.575 29.600 ;
        POLYGON 177.650 29.950 177.650 29.600 177.400 29.600 ;
        RECT 177.650 29.600 195.955 29.950 ;
        RECT 64.025 29.570 165.525 29.600 ;
        POLYGON 165.525 29.600 165.575 29.600 165.525 29.570 ;
        POLYGON 177.400 29.600 177.400 29.570 177.380 29.570 ;
        RECT 177.400 29.570 195.955 29.600 ;
        RECT 64.025 29.560 165.115 29.570 ;
        RECT 16.145 28.180 23.480 29.560 ;
        POLYGON 23.480 29.560 23.730 28.180 23.480 28.180 ;
        POLYGON 64.025 29.560 64.845 29.560 64.845 28.360 ;
        RECT 64.845 29.310 165.115 29.560 ;
        POLYGON 165.115 29.570 165.525 29.570 165.115 29.310 ;
        POLYGON 177.380 29.570 177.380 29.530 177.350 29.530 ;
        RECT 177.380 29.530 195.955 29.570 ;
        POLYGON 177.350 29.530 177.350 29.350 177.210 29.350 ;
        RECT 177.350 29.350 195.955 29.530 ;
        POLYGON 177.210 29.350 177.210 29.310 177.180 29.310 ;
        RECT 177.210 29.310 195.955 29.350 ;
        RECT 64.845 28.855 164.295 29.310 ;
        POLYGON 164.295 29.310 165.115 29.310 164.295 28.855 ;
        POLYGON 177.180 29.310 177.180 29.005 176.940 29.005 ;
        RECT 177.180 29.005 195.955 29.310 ;
        POLYGON 176.940 29.005 176.940 28.855 176.825 28.855 ;
        RECT 176.940 28.855 195.955 29.005 ;
        RECT 64.845 28.775 164.145 28.855 ;
        POLYGON 164.145 28.855 164.295 28.855 164.145 28.775 ;
        POLYGON 176.825 28.855 176.825 28.775 176.765 28.775 ;
        RECT 176.825 28.775 195.955 28.855 ;
        RECT 64.845 28.765 164.130 28.775 ;
        POLYGON 164.130 28.775 164.145 28.775 164.130 28.765 ;
        POLYGON 176.765 28.775 176.765 28.765 176.755 28.765 ;
        RECT 176.765 28.765 195.955 28.775 ;
        RECT 64.845 28.360 163.105 28.765 ;
        POLYGON 64.845 28.360 64.980 28.360 64.980 28.180 ;
        RECT 64.980 28.265 163.105 28.360 ;
        POLYGON 163.105 28.765 164.130 28.765 163.105 28.265 ;
        POLYGON 176.755 28.760 176.755 28.650 176.670 28.650 ;
        RECT 176.755 28.650 195.955 28.765 ;
        POLYGON 176.670 28.650 176.670 28.435 176.500 28.435 ;
        RECT 176.670 28.435 195.955 28.650 ;
        POLYGON 176.500 28.435 176.500 28.265 176.355 28.265 ;
        RECT 176.500 28.270 195.955 28.435 ;
        POLYGON 195.955 30.475 196.580 30.475 195.955 28.270 ;
        POLYGON 215.875 30.475 215.885 30.475 215.885 30.465 ;
        RECT 215.885 30.465 233.620 30.475 ;
        POLYGON 233.620 30.530 233.715 30.465 233.620 30.465 ;
        POLYGON 261.795 30.530 261.795 30.465 261.715 30.465 ;
        RECT 261.795 30.465 272.985 30.530 ;
        POLYGON 272.985 30.655 273.120 30.655 272.985 30.465 ;
        POLYGON 286.690 30.655 286.690 30.475 286.665 30.475 ;
        RECT 286.690 30.475 303.120 30.655 ;
        POLYGON 215.885 30.465 216.240 30.465 216.240 30.025 ;
        RECT 216.240 30.355 233.715 30.465 ;
        POLYGON 233.715 30.465 233.880 30.355 233.715 30.355 ;
        POLYGON 261.715 30.465 261.715 30.445 261.690 30.445 ;
        RECT 261.715 30.445 272.340 30.465 ;
        POLYGON 261.690 30.445 261.690 30.355 261.570 30.355 ;
        RECT 261.690 30.355 272.340 30.445 ;
        RECT 216.240 30.270 233.880 30.355 ;
        POLYGON 233.880 30.355 234.005 30.270 233.880 30.270 ;
        POLYGON 261.570 30.355 261.570 30.270 261.460 30.270 ;
        RECT 261.570 30.270 272.340 30.355 ;
        RECT 216.240 30.120 234.010 30.270 ;
        POLYGON 234.010 30.270 234.230 30.120 234.010 30.120 ;
        POLYGON 261.460 30.270 261.460 30.120 261.265 30.120 ;
        RECT 261.460 30.120 272.340 30.270 ;
        RECT 216.240 30.025 234.230 30.120 ;
        POLYGON 234.230 30.120 234.375 30.025 234.230 30.025 ;
        POLYGON 261.265 30.120 261.265 30.025 261.140 30.025 ;
        RECT 261.265 30.025 272.340 30.120 ;
        POLYGON 216.240 30.025 216.790 30.025 216.790 29.380 ;
        RECT 216.790 29.905 234.380 30.025 ;
        POLYGON 234.380 30.025 234.570 29.905 234.380 29.905 ;
        POLYGON 261.140 30.025 261.140 29.970 261.070 29.970 ;
        RECT 261.140 29.970 272.340 30.025 ;
        POLYGON 261.070 29.970 261.070 29.905 260.975 29.905 ;
        RECT 261.070 29.905 272.340 29.970 ;
        RECT 216.790 29.655 234.570 29.905 ;
        POLYGON 234.570 29.905 234.965 29.655 234.570 29.655 ;
        POLYGON 260.975 29.905 260.975 29.900 260.970 29.900 ;
        RECT 260.975 29.900 272.340 29.905 ;
        POLYGON 260.970 29.900 260.970 29.655 260.620 29.655 ;
        RECT 260.970 29.655 272.340 29.900 ;
        RECT 216.790 29.545 234.965 29.655 ;
        POLYGON 234.965 29.655 235.160 29.545 234.965 29.545 ;
        POLYGON 260.620 29.655 260.620 29.630 260.585 29.630 ;
        RECT 260.620 29.630 272.340 29.655 ;
        POLYGON 260.585 29.630 260.585 29.625 260.575 29.625 ;
        RECT 260.585 29.625 272.340 29.630 ;
        POLYGON 260.575 29.625 260.575 29.545 260.450 29.545 ;
        RECT 260.575 29.550 272.340 29.625 ;
        POLYGON 272.340 30.465 272.985 30.465 272.340 29.550 ;
        POLYGON 286.665 30.465 286.665 29.560 286.540 29.560 ;
        RECT 286.665 29.560 303.120 30.475 ;
        RECT 260.575 29.545 272.205 29.550 ;
        RECT 216.790 29.535 235.160 29.545 ;
        POLYGON 235.160 29.545 235.175 29.535 235.160 29.535 ;
        POLYGON 260.450 29.545 260.450 29.535 260.430 29.535 ;
        RECT 260.450 29.535 272.205 29.545 ;
        RECT 216.790 29.480 235.175 29.535 ;
        POLYGON 235.175 29.535 235.275 29.480 235.175 29.480 ;
        POLYGON 260.430 29.535 260.430 29.480 260.345 29.480 ;
        RECT 260.430 29.480 272.205 29.535 ;
        RECT 216.790 29.380 235.275 29.480 ;
        POLYGON 235.275 29.480 235.445 29.380 235.275 29.380 ;
        POLYGON 260.345 29.480 260.345 29.380 260.185 29.380 ;
        RECT 260.345 29.380 272.205 29.480 ;
        POLYGON 272.205 29.550 272.340 29.550 272.205 29.380 ;
        POLYGON 286.540 29.550 286.540 29.380 286.515 29.380 ;
        RECT 286.540 29.380 303.120 29.560 ;
        POLYGON 216.790 29.380 217.025 29.380 217.025 29.110 ;
        RECT 217.025 29.220 235.445 29.380 ;
        POLYGON 235.445 29.380 235.720 29.220 235.445 29.220 ;
        POLYGON 260.185 29.380 260.185 29.355 260.145 29.355 ;
        RECT 260.185 29.375 272.205 29.380 ;
        RECT 260.185 29.355 271.490 29.375 ;
        POLYGON 260.145 29.355 260.145 29.335 260.115 29.335 ;
        RECT 260.145 29.335 271.490 29.355 ;
        POLYGON 260.115 29.335 260.115 29.220 259.910 29.220 ;
        RECT 260.115 29.220 271.490 29.335 ;
        RECT 217.025 29.195 235.720 29.220 ;
        POLYGON 235.720 29.220 235.765 29.195 235.720 29.195 ;
        POLYGON 259.910 29.220 259.910 29.195 259.865 29.195 ;
        RECT 259.910 29.195 271.490 29.220 ;
        RECT 217.025 29.110 235.765 29.195 ;
        POLYGON 217.025 29.110 217.120 29.110 217.120 28.995 ;
        RECT 217.120 29.070 235.765 29.110 ;
        POLYGON 235.765 29.195 236.005 29.070 235.765 29.070 ;
        POLYGON 259.865 29.195 259.865 29.070 259.640 29.070 ;
        RECT 259.865 29.070 271.490 29.195 ;
        RECT 217.120 28.995 236.005 29.070 ;
        POLYGON 217.120 28.995 217.790 28.995 217.790 28.270 ;
        RECT 217.790 28.860 236.005 28.995 ;
        POLYGON 236.005 29.070 236.390 28.860 236.005 28.860 ;
        POLYGON 259.640 29.070 259.640 28.970 259.455 28.970 ;
        RECT 259.640 28.970 271.490 29.070 ;
        POLYGON 259.455 28.970 259.455 28.860 259.255 28.860 ;
        RECT 259.455 28.860 271.490 28.970 ;
        RECT 217.790 28.620 236.390 28.860 ;
        POLYGON 236.390 28.860 236.870 28.620 236.390 28.620 ;
        POLYGON 259.255 28.860 259.255 28.835 259.210 28.835 ;
        RECT 259.255 28.835 271.490 28.860 ;
        POLYGON 259.210 28.835 259.210 28.790 259.130 28.790 ;
        RECT 259.210 28.790 271.490 28.835 ;
        POLYGON 259.130 28.790 259.130 28.620 258.790 28.620 ;
        RECT 259.130 28.620 271.490 28.790 ;
        RECT 217.790 28.545 236.875 28.620 ;
        POLYGON 236.875 28.620 237.025 28.545 236.875 28.545 ;
        POLYGON 258.790 28.620 258.790 28.600 258.750 28.600 ;
        RECT 258.790 28.600 271.490 28.620 ;
        POLYGON 258.750 28.600 258.750 28.560 258.665 28.560 ;
        RECT 258.750 28.560 271.490 28.600 ;
        POLYGON 258.660 28.560 258.660 28.545 258.630 28.545 ;
        RECT 258.660 28.545 271.490 28.560 ;
        RECT 217.790 28.425 237.025 28.545 ;
        POLYGON 237.025 28.545 237.270 28.425 237.025 28.425 ;
        POLYGON 258.630 28.545 258.630 28.425 258.390 28.425 ;
        RECT 258.630 28.460 271.490 28.545 ;
        POLYGON 271.490 29.375 272.205 29.375 271.490 28.460 ;
        POLYGON 286.515 29.380 286.515 28.460 286.345 28.460 ;
        RECT 286.515 28.460 303.120 29.380 ;
        RECT 258.630 28.425 271.315 28.460 ;
        RECT 217.790 28.270 237.270 28.425 ;
        RECT 176.500 28.265 195.225 28.270 ;
        RECT 64.980 28.180 162.565 28.265 ;
        RECT 16.145 23.645 23.730 28.180 ;
        POLYGON 23.730 28.180 24.555 23.645 23.730 23.645 ;
        POLYGON 64.980 28.180 66.125 28.180 66.125 26.670 ;
        RECT 66.125 28.035 162.565 28.180 ;
        POLYGON 162.565 28.265 163.105 28.265 162.565 28.035 ;
        POLYGON 176.355 28.265 176.355 28.035 176.160 28.035 ;
        RECT 176.355 28.035 195.225 28.265 ;
        RECT 66.125 27.815 162.055 28.035 ;
        POLYGON 162.055 28.035 162.565 28.035 162.055 27.815 ;
        POLYGON 176.160 28.035 176.160 27.815 175.975 27.815 ;
        RECT 176.160 27.815 195.225 28.035 ;
        RECT 66.125 27.760 161.905 27.815 ;
        POLYGON 161.905 27.815 162.055 27.815 161.905 27.760 ;
        POLYGON 175.975 27.815 175.975 27.810 175.970 27.810 ;
        RECT 175.975 27.810 195.225 27.815 ;
        POLYGON 175.970 27.810 175.970 27.760 175.930 27.760 ;
        RECT 175.970 27.760 195.225 27.810 ;
        RECT 66.125 27.505 161.215 27.760 ;
        POLYGON 161.215 27.760 161.905 27.760 161.215 27.505 ;
        POLYGON 175.930 27.760 175.930 27.505 175.715 27.505 ;
        RECT 175.930 27.505 195.225 27.760 ;
        RECT 66.125 27.415 160.970 27.505 ;
        POLYGON 160.970 27.505 161.215 27.505 160.970 27.415 ;
        POLYGON 175.715 27.505 175.715 27.485 175.700 27.485 ;
        RECT 175.715 27.485 195.225 27.505 ;
        POLYGON 175.700 27.485 175.700 27.465 175.685 27.465 ;
        RECT 175.700 27.465 195.225 27.485 ;
        POLYGON 175.685 27.465 175.685 27.415 175.640 27.415 ;
        RECT 175.685 27.415 195.225 27.465 ;
        RECT 66.125 27.375 160.850 27.415 ;
        POLYGON 160.850 27.415 160.970 27.415 160.850 27.375 ;
        POLYGON 175.640 27.415 175.640 27.375 175.605 27.375 ;
        RECT 175.640 27.375 195.225 27.415 ;
        RECT 66.125 27.345 160.750 27.375 ;
        POLYGON 160.750 27.375 160.850 27.375 160.750 27.345 ;
        POLYGON 175.605 27.370 175.605 27.345 175.580 27.345 ;
        RECT 175.605 27.345 195.225 27.375 ;
        RECT 66.125 27.335 160.745 27.345 ;
        POLYGON 175.580 27.345 175.580 27.340 175.575 27.340 ;
        RECT 175.580 27.340 195.225 27.345 ;
        POLYGON 160.745 27.340 160.750 27.335 160.745 27.335 ;
        POLYGON 175.575 27.340 175.575 27.335 175.570 27.335 ;
        RECT 175.575 27.335 195.225 27.340 ;
        RECT 66.125 27.290 160.750 27.335 ;
        POLYGON 160.750 27.335 160.785 27.290 160.750 27.290 ;
        POLYGON 175.570 27.335 175.570 27.290 175.530 27.290 ;
        RECT 175.570 27.290 195.225 27.335 ;
        RECT 66.125 27.230 160.785 27.290 ;
        POLYGON 160.785 27.290 160.830 27.230 160.785 27.230 ;
        RECT 66.125 27.205 160.830 27.230 ;
        POLYGON 175.530 27.290 175.530 27.225 175.470 27.225 ;
        RECT 175.530 27.225 195.225 27.290 ;
        POLYGON 160.830 27.225 160.850 27.205 160.830 27.205 ;
        POLYGON 175.470 27.225 175.470 27.210 175.455 27.210 ;
        RECT 175.470 27.210 195.225 27.225 ;
        RECT 66.125 27.105 160.850 27.205 ;
        POLYGON 160.850 27.205 160.925 27.105 160.850 27.105 ;
        POLYGON 175.455 27.205 175.455 27.145 175.400 27.145 ;
        RECT 175.455 27.145 195.225 27.210 ;
        POLYGON 175.400 27.145 175.400 27.105 175.360 27.105 ;
        RECT 175.400 27.105 195.225 27.145 ;
        RECT 66.125 27.070 160.925 27.105 ;
        POLYGON 160.925 27.105 160.950 27.070 160.925 27.070 ;
        POLYGON 175.360 27.105 175.360 27.070 175.330 27.070 ;
        RECT 175.360 27.070 195.225 27.105 ;
        RECT 66.125 27.065 160.950 27.070 ;
        POLYGON 160.950 27.070 160.955 27.065 160.950 27.065 ;
        POLYGON 175.330 27.070 175.330 27.065 175.325 27.065 ;
        RECT 175.330 27.065 195.225 27.070 ;
        RECT 66.125 27.055 160.955 27.065 ;
        POLYGON 160.955 27.065 160.960 27.055 160.955 27.055 ;
        POLYGON 175.325 27.065 175.325 27.055 175.315 27.055 ;
        RECT 175.325 27.055 195.225 27.065 ;
        RECT 66.125 26.965 160.960 27.055 ;
        POLYGON 160.960 27.055 161.030 26.965 160.960 26.965 ;
        POLYGON 175.315 27.055 175.315 26.965 175.235 26.965 ;
        RECT 175.315 26.965 195.225 27.055 ;
        RECT 66.125 26.955 161.030 26.965 ;
        POLYGON 161.030 26.965 161.035 26.955 161.030 26.955 ;
        POLYGON 175.235 26.965 175.235 26.955 175.225 26.955 ;
        RECT 175.235 26.955 195.225 26.965 ;
        RECT 66.125 26.850 161.035 26.955 ;
        POLYGON 161.035 26.955 161.115 26.850 161.035 26.850 ;
        POLYGON 175.225 26.955 175.225 26.850 175.130 26.850 ;
        RECT 175.225 26.850 195.225 26.955 ;
        RECT 66.125 26.830 161.115 26.850 ;
        POLYGON 161.115 26.850 161.130 26.830 161.115 26.830 ;
        POLYGON 175.130 26.850 175.130 26.830 175.110 26.830 ;
        RECT 175.130 26.830 195.225 26.850 ;
        RECT 66.125 26.765 161.130 26.830 ;
        POLYGON 161.130 26.830 161.180 26.765 161.130 26.765 ;
        RECT 66.125 26.720 161.180 26.765 ;
        POLYGON 175.110 26.830 175.110 26.760 175.045 26.760 ;
        RECT 175.110 26.760 195.225 26.830 ;
        POLYGON 161.180 26.760 161.215 26.720 161.180 26.720 ;
        POLYGON 175.045 26.760 175.045 26.720 175.010 26.720 ;
        RECT 175.045 26.720 195.225 26.760 ;
        RECT 66.125 26.670 161.215 26.720 ;
        POLYGON 66.125 26.670 67.385 26.670 67.385 25.000 ;
        RECT 67.385 26.545 161.215 26.670 ;
        POLYGON 161.215 26.720 161.345 26.545 161.215 26.545 ;
        RECT 67.385 26.510 161.345 26.545 ;
        POLYGON 175.010 26.720 175.010 26.540 174.845 26.540 ;
        RECT 175.010 26.540 195.225 26.720 ;
        POLYGON 161.345 26.540 161.370 26.510 161.345 26.510 ;
        POLYGON 174.845 26.540 174.845 26.510 174.820 26.510 ;
        RECT 174.845 26.510 195.225 26.540 ;
        RECT 67.385 26.465 161.370 26.510 ;
        POLYGON 161.370 26.510 161.405 26.465 161.370 26.465 ;
        RECT 67.385 26.435 161.405 26.465 ;
        POLYGON 174.820 26.510 174.820 26.460 174.775 26.460 ;
        RECT 174.820 26.460 195.225 26.510 ;
        POLYGON 161.405 26.460 161.425 26.435 161.405 26.435 ;
        POLYGON 174.775 26.460 174.775 26.435 174.750 26.435 ;
        RECT 174.775 26.435 195.225 26.460 ;
        RECT 67.385 26.315 161.425 26.435 ;
        POLYGON 161.425 26.435 161.515 26.315 161.425 26.315 ;
        POLYGON 174.750 26.435 174.750 26.315 174.640 26.315 ;
        RECT 174.750 26.315 195.225 26.435 ;
        RECT 67.385 26.285 161.515 26.315 ;
        POLYGON 161.515 26.315 161.540 26.285 161.515 26.285 ;
        POLYGON 174.640 26.315 174.640 26.285 174.615 26.285 ;
        RECT 174.640 26.285 195.225 26.315 ;
        RECT 67.385 26.035 161.540 26.285 ;
        POLYGON 161.540 26.285 161.725 26.035 161.540 26.035 ;
        POLYGON 174.615 26.285 174.615 26.035 174.365 26.035 ;
        RECT 174.615 26.095 195.225 26.285 ;
        POLYGON 195.225 28.270 195.955 28.270 195.225 26.095 ;
        POLYGON 217.790 28.270 217.800 28.270 217.800 28.255 ;
        RECT 217.800 28.255 237.270 28.270 ;
        POLYGON 237.270 28.425 237.645 28.255 237.270 28.255 ;
        POLYGON 258.390 28.425 258.390 28.380 258.300 28.380 ;
        RECT 258.390 28.380 271.315 28.425 ;
        POLYGON 258.295 28.380 258.295 28.290 258.110 28.290 ;
        RECT 258.295 28.290 271.315 28.380 ;
        POLYGON 258.110 28.290 258.110 28.255 258.025 28.255 ;
        RECT 258.110 28.255 271.315 28.290 ;
        POLYGON 271.315 28.460 271.490 28.460 271.315 28.255 ;
        POLYGON 286.345 28.460 286.345 28.270 286.310 28.270 ;
        RECT 286.345 28.270 303.120 28.460 ;
        POLYGON 217.800 28.255 217.975 28.255 217.975 28.065 ;
        RECT 217.975 28.245 237.645 28.255 ;
        POLYGON 237.645 28.255 237.670 28.245 237.645 28.245 ;
        POLYGON 258.025 28.255 258.025 28.245 258.005 28.245 ;
        RECT 258.025 28.250 271.315 28.255 ;
        RECT 258.025 28.245 271.155 28.250 ;
        RECT 217.975 28.195 237.670 28.245 ;
        POLYGON 237.670 28.245 237.775 28.195 237.670 28.195 ;
        POLYGON 258.005 28.245 258.005 28.195 257.885 28.195 ;
        RECT 258.005 28.195 271.155 28.245 ;
        RECT 217.975 28.125 237.775 28.195 ;
        POLYGON 237.775 28.195 237.940 28.125 237.775 28.125 ;
        POLYGON 257.885 28.195 257.885 28.180 257.850 28.180 ;
        RECT 257.885 28.180 271.155 28.195 ;
        POLYGON 257.845 28.180 257.845 28.125 257.715 28.125 ;
        RECT 257.845 28.125 271.155 28.180 ;
        RECT 217.975 28.065 237.940 28.125 ;
        POLYGON 237.940 28.125 238.070 28.065 237.940 28.065 ;
        POLYGON 257.715 28.125 257.715 28.065 257.575 28.065 ;
        RECT 257.715 28.065 271.155 28.125 ;
        POLYGON 271.155 28.250 271.315 28.250 271.155 28.065 ;
        POLYGON 286.310 28.255 286.310 28.065 286.275 28.065 ;
        RECT 286.310 28.065 303.120 28.270 ;
        POLYGON 217.975 28.065 218.035 28.065 218.035 28.005 ;
        RECT 218.035 28.005 238.070 28.065 ;
        POLYGON 218.035 28.005 218.975 28.005 218.975 27.040 ;
        RECT 218.975 27.965 238.070 28.005 ;
        POLYGON 238.070 28.065 238.315 27.965 238.070 27.965 ;
        POLYGON 257.575 28.065 257.575 27.995 257.415 27.995 ;
        RECT 257.575 28.060 271.155 28.065 ;
        RECT 257.575 27.995 270.585 28.060 ;
        POLYGON 257.415 27.995 257.415 27.965 257.345 27.965 ;
        RECT 257.415 27.965 270.585 27.995 ;
        RECT 218.975 27.805 238.320 27.965 ;
        POLYGON 238.320 27.965 238.705 27.805 238.320 27.805 ;
        POLYGON 257.345 27.965 257.345 27.865 257.115 27.865 ;
        RECT 257.345 27.865 270.585 27.965 ;
        POLYGON 257.115 27.865 257.115 27.840 257.055 27.840 ;
        RECT 257.115 27.840 270.585 27.865 ;
        POLYGON 257.055 27.840 257.055 27.805 256.960 27.805 ;
        RECT 257.055 27.805 270.585 27.840 ;
        RECT 218.975 27.730 238.710 27.805 ;
        POLYGON 238.710 27.805 238.880 27.730 238.710 27.730 ;
        POLYGON 256.960 27.805 256.960 27.730 256.760 27.730 ;
        RECT 256.960 27.730 270.585 27.805 ;
        RECT 218.975 27.700 238.880 27.730 ;
        POLYGON 238.880 27.730 238.965 27.700 238.880 27.700 ;
        POLYGON 256.760 27.730 256.760 27.700 256.680 27.700 ;
        RECT 256.760 27.700 270.585 27.730 ;
        RECT 218.975 27.575 238.965 27.700 ;
        POLYGON 238.965 27.700 239.300 27.575 238.965 27.575 ;
        POLYGON 256.680 27.700 256.680 27.580 256.360 27.580 ;
        RECT 256.680 27.580 270.585 27.700 ;
        POLYGON 256.360 27.580 256.360 27.575 256.345 27.575 ;
        RECT 256.360 27.575 270.585 27.580 ;
        RECT 218.975 27.460 239.300 27.575 ;
        POLYGON 239.300 27.575 239.615 27.460 239.300 27.460 ;
        POLYGON 256.345 27.575 256.345 27.570 256.330 27.570 ;
        RECT 256.345 27.570 270.585 27.575 ;
        POLYGON 256.330 27.570 256.330 27.460 256.030 27.460 ;
        RECT 256.330 27.460 270.585 27.570 ;
        RECT 218.975 27.440 239.615 27.460 ;
        POLYGON 239.615 27.460 239.670 27.440 239.615 27.440 ;
        POLYGON 256.030 27.460 256.030 27.440 255.975 27.440 ;
        RECT 256.030 27.440 270.585 27.460 ;
        RECT 218.975 27.425 239.670 27.440 ;
        POLYGON 239.670 27.440 239.710 27.425 239.670 27.425 ;
        POLYGON 255.975 27.440 255.975 27.425 255.935 27.425 ;
        RECT 255.975 27.425 270.585 27.440 ;
        RECT 218.975 27.245 239.710 27.425 ;
        POLYGON 239.710 27.425 240.250 27.245 239.710 27.245 ;
        POLYGON 255.935 27.425 255.935 27.415 255.905 27.415 ;
        RECT 255.935 27.415 270.585 27.425 ;
        POLYGON 255.905 27.415 255.905 27.245 255.360 27.245 ;
        RECT 255.905 27.385 270.585 27.415 ;
        POLYGON 270.585 28.060 271.155 28.060 270.585 27.385 ;
        POLYGON 286.275 28.065 286.275 27.385 286.150 27.385 ;
        RECT 286.275 27.385 303.120 28.065 ;
        RECT 255.905 27.245 269.610 27.385 ;
        RECT 218.975 27.145 240.255 27.245 ;
        POLYGON 240.255 27.245 240.545 27.145 240.255 27.145 ;
        POLYGON 255.360 27.245 255.360 27.225 255.295 27.225 ;
        RECT 255.360 27.225 269.610 27.245 ;
        POLYGON 255.295 27.225 255.295 27.180 255.160 27.180 ;
        RECT 255.295 27.180 269.610 27.225 ;
        POLYGON 255.160 27.180 255.160 27.145 255.045 27.145 ;
        RECT 255.160 27.145 269.610 27.180 ;
        RECT 218.975 27.115 240.545 27.145 ;
        POLYGON 240.545 27.145 240.660 27.115 240.545 27.115 ;
        POLYGON 255.045 27.145 255.045 27.115 254.950 27.115 ;
        RECT 255.045 27.115 269.610 27.145 ;
        RECT 218.975 27.090 240.660 27.115 ;
        POLYGON 240.660 27.115 240.740 27.090 240.660 27.090 ;
        POLYGON 254.950 27.115 254.950 27.090 254.870 27.090 ;
        RECT 254.950 27.090 269.610 27.115 ;
        RECT 218.975 27.040 240.745 27.090 ;
        POLYGON 218.975 27.040 219.265 27.040 219.265 26.765 ;
        RECT 219.265 26.920 240.745 27.040 ;
        POLYGON 240.745 27.090 241.315 26.920 240.745 26.920 ;
        POLYGON 254.870 27.090 254.870 27.035 254.670 27.035 ;
        RECT 254.870 27.035 269.610 27.090 ;
        POLYGON 254.670 27.035 254.670 26.920 254.245 26.920 ;
        RECT 254.670 26.920 269.610 27.035 ;
        RECT 219.265 26.895 241.315 26.920 ;
        POLYGON 241.315 26.920 241.400 26.895 241.315 26.895 ;
        POLYGON 254.245 26.920 254.245 26.895 254.145 26.895 ;
        RECT 254.245 26.895 269.610 26.920 ;
        RECT 219.265 26.825 241.400 26.895 ;
        POLYGON 241.400 26.895 241.675 26.825 241.400 26.825 ;
        POLYGON 254.145 26.895 254.145 26.855 253.990 26.855 ;
        RECT 254.145 26.855 269.610 26.895 ;
        POLYGON 253.985 26.855 253.985 26.825 253.875 26.825 ;
        RECT 253.985 26.825 269.610 26.855 ;
        RECT 219.265 26.765 241.680 26.825 ;
        POLYGON 219.265 26.765 219.950 26.765 219.950 26.110 ;
        RECT 219.950 26.675 241.680 26.765 ;
        POLYGON 241.680 26.825 242.260 26.675 241.680 26.675 ;
        POLYGON 253.875 26.825 253.875 26.790 253.750 26.790 ;
        RECT 253.875 26.790 269.610 26.825 ;
        POLYGON 253.750 26.790 253.750 26.715 253.405 26.715 ;
        RECT 253.750 26.715 269.610 26.790 ;
        POLYGON 253.405 26.715 253.405 26.675 253.225 26.675 ;
        RECT 253.405 26.675 269.610 26.715 ;
        RECT 219.950 26.665 242.260 26.675 ;
        POLYGON 242.260 26.675 242.305 26.665 242.260 26.665 ;
        POLYGON 253.225 26.675 253.225 26.665 253.180 26.665 ;
        RECT 253.225 26.665 269.610 26.675 ;
        RECT 219.950 26.650 242.310 26.665 ;
        POLYGON 242.310 26.665 242.380 26.650 242.310 26.650 ;
        POLYGON 253.180 26.665 253.180 26.660 253.155 26.660 ;
        RECT 253.180 26.660 269.610 26.665 ;
        POLYGON 253.155 26.660 253.155 26.650 253.110 26.650 ;
        RECT 253.155 26.650 269.610 26.660 ;
        RECT 219.950 26.580 242.385 26.650 ;
        POLYGON 242.385 26.650 242.720 26.580 242.385 26.580 ;
        POLYGON 253.110 26.650 253.110 26.585 252.820 26.585 ;
        RECT 253.110 26.585 269.610 26.650 ;
        POLYGON 252.820 26.585 252.820 26.580 252.795 26.580 ;
        RECT 252.820 26.580 269.610 26.585 ;
        RECT 219.950 26.440 242.720 26.580 ;
        POLYGON 242.720 26.580 243.370 26.440 242.720 26.440 ;
        POLYGON 252.795 26.580 252.795 26.540 252.610 26.540 ;
        RECT 252.795 26.540 269.610 26.580 ;
        POLYGON 252.610 26.540 252.610 26.455 252.120 26.455 ;
        RECT 252.610 26.455 269.610 26.540 ;
        POLYGON 252.120 26.455 252.120 26.450 252.080 26.450 ;
        RECT 252.120 26.450 269.610 26.455 ;
        POLYGON 252.080 26.450 252.080 26.440 252.025 26.440 ;
        RECT 252.080 26.440 269.610 26.450 ;
        RECT 219.950 26.430 243.370 26.440 ;
        POLYGON 243.370 26.440 243.450 26.430 243.370 26.430 ;
        POLYGON 252.025 26.440 252.025 26.430 251.965 26.430 ;
        RECT 252.025 26.430 269.610 26.440 ;
        RECT 219.950 26.375 243.455 26.430 ;
        POLYGON 243.455 26.430 243.780 26.375 243.455 26.375 ;
        POLYGON 251.965 26.430 251.965 26.375 251.655 26.375 ;
        RECT 251.965 26.375 269.610 26.430 ;
        RECT 219.950 26.335 243.780 26.375 ;
        POLYGON 243.780 26.375 244.040 26.335 243.780 26.335 ;
        POLYGON 251.655 26.375 251.655 26.340 251.455 26.340 ;
        RECT 251.655 26.340 269.610 26.375 ;
        POLYGON 251.455 26.340 251.455 26.335 251.415 26.335 ;
        RECT 251.455 26.335 269.610 26.340 ;
        RECT 219.950 26.265 244.040 26.335 ;
        POLYGON 244.040 26.335 244.500 26.265 244.040 26.265 ;
        POLYGON 251.415 26.335 251.415 26.295 251.105 26.295 ;
        RECT 251.415 26.315 269.610 26.335 ;
        POLYGON 269.610 27.385 270.585 27.385 269.610 26.315 ;
        POLYGON 286.150 27.380 286.150 26.315 285.955 26.315 ;
        RECT 286.150 26.315 303.120 27.385 ;
        RECT 251.415 26.295 269.390 26.315 ;
        POLYGON 251.105 26.295 251.105 26.285 251.000 26.285 ;
        RECT 251.105 26.285 269.390 26.295 ;
        POLYGON 251.000 26.285 251.000 26.265 250.845 26.265 ;
        RECT 251.000 26.265 269.390 26.285 ;
        RECT 219.950 26.260 244.500 26.265 ;
        POLYGON 244.500 26.265 244.520 26.260 244.500 26.260 ;
        POLYGON 250.845 26.265 250.845 26.260 250.805 26.260 ;
        RECT 250.845 26.260 269.390 26.265 ;
        RECT 219.950 26.225 244.530 26.260 ;
        POLYGON 244.530 26.260 244.860 26.225 244.530 26.225 ;
        POLYGON 250.805 26.260 250.805 26.225 250.535 26.225 ;
        RECT 250.805 26.225 269.390 26.260 ;
        RECT 219.950 26.145 244.860 26.225 ;
        POLYGON 244.860 26.225 245.600 26.145 244.860 26.145 ;
        POLYGON 250.535 26.225 250.535 26.195 250.295 26.195 ;
        RECT 250.535 26.195 269.390 26.225 ;
        POLYGON 250.295 26.195 250.295 26.185 250.195 26.185 ;
        RECT 250.295 26.185 269.390 26.195 ;
        POLYGON 250.195 26.185 250.195 26.165 249.925 26.165 ;
        RECT 250.195 26.165 269.390 26.185 ;
        POLYGON 249.920 26.165 249.920 26.145 249.665 26.145 ;
        RECT 249.920 26.145 269.390 26.165 ;
        RECT 219.950 26.140 245.605 26.145 ;
        POLYGON 245.605 26.145 245.645 26.140 245.605 26.140 ;
        POLYGON 249.665 26.145 249.665 26.140 249.600 26.140 ;
        RECT 249.665 26.140 269.390 26.145 ;
        RECT 219.950 26.125 245.645 26.140 ;
        POLYGON 245.645 26.140 245.950 26.125 245.645 26.125 ;
        POLYGON 249.600 26.140 249.600 26.125 249.410 26.125 ;
        RECT 249.600 26.125 269.390 26.140 ;
        RECT 219.950 26.110 245.960 26.125 ;
        POLYGON 219.950 26.110 219.965 26.110 219.965 26.095 ;
        RECT 219.965 26.095 245.960 26.110 ;
        RECT 174.615 26.035 195.130 26.095 ;
        RECT 67.385 25.685 161.725 26.035 ;
        POLYGON 161.725 26.035 161.990 25.685 161.725 25.685 ;
        POLYGON 174.365 26.035 174.365 25.685 174.025 25.685 ;
        RECT 174.365 25.850 195.130 26.035 ;
        POLYGON 195.130 26.095 195.225 26.095 195.130 25.850 ;
        POLYGON 219.965 26.095 219.970 26.095 219.970 26.090 ;
        RECT 219.970 26.090 245.960 26.095 ;
        POLYGON 245.960 26.125 246.500 26.090 245.960 26.090 ;
        POLYGON 249.410 26.125 249.410 26.120 249.345 26.120 ;
        RECT 249.410 26.120 269.390 26.125 ;
        POLYGON 249.340 26.120 249.340 26.100 249.130 26.100 ;
        RECT 249.340 26.100 269.390 26.120 ;
        POLYGON 249.130 26.100 249.130 26.090 248.820 26.090 ;
        RECT 249.130 26.090 269.390 26.100 ;
        POLYGON 269.390 26.315 269.610 26.315 269.390 26.090 ;
        POLYGON 285.955 26.315 285.955 26.095 285.915 26.095 ;
        RECT 285.955 26.095 303.120 26.315 ;
        POLYGON 219.970 26.090 220.240 26.090 220.240 25.850 ;
        RECT 220.240 26.085 246.500 26.090 ;
        POLYGON 246.500 26.090 246.580 26.085 246.500 26.085 ;
        POLYGON 248.820 26.090 248.820 26.085 248.660 26.085 ;
        RECT 248.820 26.085 269.150 26.090 ;
        RECT 220.240 26.080 246.585 26.085 ;
        POLYGON 246.585 26.085 246.685 26.080 246.585 26.080 ;
        POLYGON 248.660 26.085 248.660 26.080 248.505 26.080 ;
        RECT 248.660 26.080 269.150 26.085 ;
        RECT 220.240 26.075 246.685 26.080 ;
        POLYGON 246.685 26.080 246.800 26.075 246.685 26.075 ;
        POLYGON 248.495 26.080 248.495 26.075 248.360 26.075 ;
        RECT 248.495 26.075 269.150 26.080 ;
        RECT 220.240 26.070 246.800 26.075 ;
        POLYGON 246.800 26.075 247.070 26.070 246.800 26.070 ;
        POLYGON 248.360 26.075 248.360 26.070 248.220 26.070 ;
        RECT 248.360 26.070 269.150 26.075 ;
        RECT 220.240 26.065 247.075 26.070 ;
        POLYGON 247.075 26.070 247.695 26.065 247.075 26.065 ;
        POLYGON 248.205 26.070 248.205 26.065 248.085 26.065 ;
        RECT 248.205 26.065 269.150 26.070 ;
        RECT 220.240 26.060 247.760 26.065 ;
        POLYGON 247.760 26.065 247.965 26.060 247.760 26.060 ;
        POLYGON 248.085 26.065 248.085 26.060 247.965 26.060 ;
        RECT 248.085 26.060 269.150 26.065 ;
        RECT 220.240 25.850 269.150 26.060 ;
        RECT 174.365 25.685 194.395 25.850 ;
        RECT 67.385 25.575 161.990 25.685 ;
        POLYGON 161.990 25.685 162.070 25.575 161.990 25.575 ;
        POLYGON 174.025 25.685 174.025 25.575 173.920 25.575 ;
        RECT 174.025 25.575 194.395 25.685 ;
        RECT 67.385 25.365 162.070 25.575 ;
        POLYGON 162.070 25.575 162.230 25.365 162.070 25.365 ;
        POLYGON 173.920 25.575 173.920 25.365 173.715 25.365 ;
        RECT 173.920 25.365 194.395 25.575 ;
        RECT 67.385 25.295 162.230 25.365 ;
        POLYGON 162.230 25.365 162.280 25.295 162.230 25.295 ;
        POLYGON 173.715 25.365 173.715 25.295 173.640 25.295 ;
        RECT 173.715 25.295 194.395 25.365 ;
        RECT 67.385 25.190 162.280 25.295 ;
        POLYGON 162.280 25.295 162.360 25.190 162.280 25.190 ;
        POLYGON 173.640 25.295 173.640 25.190 173.530 25.190 ;
        RECT 173.640 25.190 194.395 25.295 ;
        RECT 67.385 25.065 162.360 25.190 ;
        POLYGON 162.360 25.190 162.455 25.065 162.360 25.065 ;
        RECT 67.385 25.000 162.455 25.065 ;
        POLYGON 173.530 25.190 173.530 25.060 173.390 25.060 ;
        RECT 173.530 25.060 194.395 25.190 ;
        RECT 65.000 24.870 162.455 25.000 ;
        POLYGON 162.455 25.060 162.600 24.870 162.455 24.870 ;
        POLYGON 173.390 25.060 173.390 24.870 173.185 24.870 ;
        RECT 173.390 24.870 194.395 25.060 ;
        RECT 65.000 24.605 162.600 24.870 ;
        POLYGON 162.600 24.870 162.800 24.605 162.600 24.605 ;
        POLYGON 173.185 24.870 173.185 24.605 172.905 24.605 ;
        RECT 173.185 24.605 194.395 24.870 ;
        RECT 65.000 24.490 162.800 24.605 ;
        POLYGON 162.800 24.605 162.885 24.490 162.800 24.490 ;
        POLYGON 172.905 24.605 172.905 24.490 172.785 24.490 ;
        RECT 172.905 24.490 194.395 24.605 ;
        RECT 65.000 24.385 162.885 24.490 ;
        POLYGON 162.885 24.490 162.965 24.385 162.885 24.385 ;
        POLYGON 172.785 24.490 172.785 24.385 172.665 24.385 ;
        RECT 172.785 24.385 194.395 24.490 ;
        RECT 65.000 24.365 162.965 24.385 ;
        POLYGON 162.965 24.385 162.980 24.365 162.965 24.365 ;
        POLYGON 172.665 24.385 172.665 24.365 172.645 24.365 ;
        RECT 172.665 24.365 194.395 24.385 ;
        RECT 65.000 24.340 162.980 24.365 ;
        POLYGON 162.980 24.365 163.000 24.340 162.980 24.340 ;
        POLYGON 172.645 24.365 172.645 24.340 172.615 24.340 ;
        RECT 172.645 24.340 194.395 24.365 ;
        RECT 65.000 24.330 163.000 24.340 ;
        POLYGON 163.000 24.340 163.010 24.330 163.000 24.330 ;
        POLYGON 172.615 24.340 172.615 24.330 172.605 24.330 ;
        RECT 172.615 24.330 194.395 24.340 ;
        RECT 65.000 24.200 163.010 24.330 ;
        POLYGON 163.010 24.330 163.125 24.200 163.010 24.200 ;
        RECT 65.000 24.140 163.125 24.200 ;
        POLYGON 172.605 24.330 172.605 24.195 172.450 24.195 ;
        RECT 172.605 24.195 194.395 24.330 ;
        POLYGON 163.125 24.195 163.175 24.140 163.125 24.140 ;
        POLYGON 172.450 24.195 172.450 24.140 172.390 24.140 ;
        RECT 172.450 24.140 194.395 24.195 ;
        RECT 65.000 24.120 163.175 24.140 ;
        POLYGON 163.175 24.140 163.195 24.120 163.175 24.120 ;
        RECT 65.000 24.035 163.195 24.120 ;
        POLYGON 172.390 24.140 172.390 24.115 172.360 24.115 ;
        RECT 172.390 24.115 194.395 24.140 ;
        POLYGON 163.195 24.115 163.270 24.035 163.195 24.035 ;
        POLYGON 172.360 24.115 172.360 24.035 172.270 24.035 ;
        RECT 172.360 24.035 194.395 24.115 ;
        RECT 65.000 23.960 163.270 24.035 ;
        POLYGON 163.270 24.035 163.335 23.960 163.270 23.960 ;
        POLYGON 172.270 24.035 172.270 23.960 172.185 23.960 ;
        RECT 172.270 23.960 194.395 24.035 ;
        RECT 65.000 23.870 163.335 23.960 ;
        POLYGON 163.335 23.960 163.415 23.870 163.335 23.870 ;
        POLYGON 172.185 23.960 172.185 23.870 172.080 23.870 ;
        RECT 172.185 23.955 194.395 23.960 ;
        POLYGON 194.395 25.850 195.130 25.850 194.395 23.955 ;
        POLYGON 220.240 25.850 220.245 25.850 220.245 25.845 ;
        RECT 220.245 25.845 269.150 25.850 ;
        POLYGON 269.150 26.090 269.390 26.090 269.150 25.845 ;
        POLYGON 285.915 26.090 285.915 25.850 285.870 25.850 ;
        RECT 285.915 25.850 303.120 26.095 ;
        POLYGON 220.245 25.845 220.950 25.845 220.950 25.220 ;
        RECT 220.950 25.395 268.705 25.845 ;
        POLYGON 268.705 25.845 269.150 25.845 268.705 25.395 ;
        POLYGON 285.870 25.845 285.870 25.405 285.790 25.405 ;
        RECT 285.870 25.405 303.120 25.850 ;
        RECT 220.950 25.220 267.780 25.395 ;
        POLYGON 220.950 25.220 221.690 25.220 221.690 24.600 ;
        RECT 221.690 24.600 267.780 25.220 ;
        POLYGON 221.690 24.600 221.980 24.600 221.980 24.360 ;
        RECT 221.980 24.520 267.780 24.600 ;
        POLYGON 267.780 25.395 268.705 25.395 267.780 24.520 ;
        POLYGON 285.790 25.395 285.790 24.530 285.630 24.530 ;
        RECT 285.790 24.530 303.120 25.405 ;
        RECT 221.980 24.360 267.135 24.520 ;
        POLYGON 221.980 24.360 222.500 24.360 222.500 23.955 ;
        RECT 222.500 23.955 267.135 24.360 ;
        POLYGON 267.135 24.520 267.780 24.520 267.135 23.955 ;
        POLYGON 285.630 24.520 285.630 23.955 285.525 23.955 ;
        RECT 285.630 23.955 303.120 24.530 ;
        RECT 172.185 23.870 193.465 23.955 ;
        RECT 65.000 23.855 163.415 23.870 ;
        POLYGON 163.415 23.870 163.425 23.855 163.415 23.855 ;
        POLYGON 172.080 23.870 172.080 23.855 172.065 23.855 ;
        RECT 172.080 23.855 193.465 23.870 ;
        RECT 65.000 23.730 163.425 23.855 ;
        POLYGON 163.425 23.855 163.535 23.730 163.425 23.730 ;
        RECT 65.000 23.655 163.535 23.730 ;
        POLYGON 172.065 23.855 172.065 23.725 171.915 23.725 ;
        RECT 172.065 23.725 193.465 23.855 ;
        POLYGON 163.535 23.725 163.600 23.655 163.535 23.655 ;
        POLYGON 171.915 23.725 171.915 23.655 171.835 23.655 ;
        RECT 171.915 23.655 193.465 23.725 ;
        RECT 16.145 21.130 24.555 23.645 ;
        POLYGON 16.145 21.130 18.180 21.130 18.180 12.670 ;
        RECT 18.180 17.825 24.555 21.130 ;
        POLYGON 24.555 23.645 25.870 17.825 24.555 17.825 ;
        RECT 65.000 23.565 163.600 23.655 ;
        POLYGON 163.600 23.655 163.675 23.565 163.600 23.565 ;
        POLYGON 171.835 23.655 171.835 23.565 171.725 23.565 ;
        RECT 171.835 23.565 193.465 23.655 ;
        RECT 65.000 23.560 163.675 23.565 ;
        POLYGON 163.675 23.565 163.680 23.560 163.675 23.560 ;
        POLYGON 171.725 23.565 171.725 23.560 171.720 23.560 ;
        RECT 171.725 23.560 193.465 23.565 ;
        RECT 65.000 23.515 163.680 23.560 ;
        POLYGON 163.680 23.560 163.720 23.515 163.680 23.515 ;
        RECT 65.000 23.475 163.720 23.515 ;
        POLYGON 171.720 23.560 171.720 23.510 171.655 23.510 ;
        RECT 171.720 23.510 193.465 23.560 ;
        POLYGON 163.720 23.510 163.755 23.475 163.720 23.475 ;
        POLYGON 171.655 23.510 171.655 23.475 171.610 23.475 ;
        RECT 171.655 23.475 193.465 23.510 ;
        RECT 65.000 23.365 163.755 23.475 ;
        POLYGON 163.755 23.475 163.850 23.365 163.755 23.365 ;
        POLYGON 171.610 23.475 171.610 23.365 171.475 23.365 ;
        RECT 171.610 23.365 193.465 23.475 ;
        RECT 65.000 23.335 163.850 23.365 ;
        POLYGON 163.850 23.365 163.875 23.335 163.850 23.335 ;
        POLYGON 171.475 23.365 171.475 23.335 171.440 23.335 ;
        RECT 171.475 23.335 193.465 23.365 ;
        RECT 65.000 23.325 163.875 23.335 ;
        POLYGON 163.875 23.335 163.885 23.325 163.875 23.325 ;
        POLYGON 171.435 23.335 171.435 23.325 171.425 23.325 ;
        RECT 171.435 23.325 193.465 23.335 ;
        RECT 65.000 23.210 163.885 23.325 ;
        POLYGON 163.885 23.325 163.985 23.210 163.885 23.210 ;
        POLYGON 171.425 23.325 171.425 23.210 171.285 23.210 ;
        RECT 171.425 23.210 193.465 23.325 ;
        RECT 65.000 23.150 163.985 23.210 ;
        POLYGON 163.985 23.210 164.035 23.150 163.985 23.150 ;
        POLYGON 171.285 23.210 171.285 23.150 171.210 23.150 ;
        RECT 171.285 23.150 193.465 23.210 ;
        RECT 65.000 23.085 164.035 23.150 ;
        POLYGON 164.035 23.150 164.090 23.085 164.035 23.085 ;
        POLYGON 171.210 23.150 171.210 23.085 171.130 23.085 ;
        RECT 171.210 23.085 193.465 23.150 ;
        RECT 65.000 23.035 164.090 23.085 ;
        POLYGON 164.090 23.085 164.135 23.035 164.090 23.035 ;
        POLYGON 171.130 23.085 171.130 23.035 171.065 23.035 ;
        RECT 171.130 23.035 193.465 23.085 ;
        RECT 65.000 22.915 164.135 23.035 ;
        POLYGON 164.135 23.035 164.240 22.915 164.135 22.915 ;
        POLYGON 171.065 23.035 171.065 22.915 170.920 22.915 ;
        RECT 171.065 22.915 193.465 23.035 ;
        RECT 65.000 22.860 164.240 22.915 ;
        POLYGON 164.240 22.915 164.285 22.860 164.240 22.860 ;
        POLYGON 170.920 22.915 170.920 22.860 170.855 22.860 ;
        RECT 170.920 22.860 193.465 22.915 ;
        RECT 65.000 22.725 164.285 22.860 ;
        POLYGON 164.285 22.860 164.405 22.725 164.285 22.725 ;
        POLYGON 170.855 22.860 170.855 22.725 170.675 22.725 ;
        RECT 170.855 22.725 193.465 22.860 ;
        RECT 65.000 22.670 164.405 22.725 ;
        POLYGON 164.405 22.725 164.450 22.670 164.405 22.670 ;
        POLYGON 170.675 22.725 170.675 22.670 170.600 22.670 ;
        RECT 170.675 22.670 193.465 22.725 ;
        RECT 65.000 22.565 164.450 22.670 ;
        POLYGON 164.450 22.670 164.545 22.565 164.450 22.565 ;
        RECT 65.000 22.550 164.545 22.565 ;
        POLYGON 170.600 22.670 170.600 22.560 170.455 22.560 ;
        RECT 170.600 22.560 193.465 22.670 ;
        POLYGON 164.545 22.560 164.555 22.550 164.545 22.550 ;
        POLYGON 170.455 22.560 170.455 22.550 170.440 22.550 ;
        RECT 170.455 22.550 193.465 22.560 ;
        RECT 65.000 22.415 164.555 22.550 ;
        POLYGON 164.555 22.550 164.675 22.415 164.555 22.415 ;
        POLYGON 170.440 22.550 170.440 22.415 170.260 22.415 ;
        RECT 170.440 22.415 193.465 22.550 ;
        RECT 65.000 22.270 164.675 22.415 ;
        POLYGON 164.675 22.415 164.800 22.270 164.675 22.270 ;
        POLYGON 170.260 22.415 170.260 22.270 170.065 22.270 ;
        RECT 170.260 22.270 193.465 22.415 ;
        RECT 65.000 22.150 164.800 22.270 ;
        POLYGON 164.800 22.270 164.905 22.150 164.800 22.150 ;
        POLYGON 170.065 22.270 170.065 22.150 169.900 22.150 ;
        RECT 170.065 22.150 193.465 22.270 ;
        RECT 65.000 22.130 164.905 22.150 ;
        POLYGON 164.905 22.150 164.920 22.130 164.905 22.130 ;
        POLYGON 169.900 22.150 169.900 22.130 169.875 22.130 ;
        RECT 169.900 22.130 193.465 22.150 ;
        RECT 65.000 22.110 164.920 22.130 ;
        POLYGON 164.920 22.130 164.940 22.110 164.920 22.110 ;
        POLYGON 169.875 22.130 169.875 22.110 169.855 22.110 ;
        RECT 169.875 22.110 193.465 22.130 ;
        RECT 65.000 21.975 164.940 22.110 ;
        POLYGON 164.940 22.110 165.055 21.975 164.940 21.975 ;
        POLYGON 169.855 22.110 169.855 21.975 169.655 21.975 ;
        RECT 169.855 21.975 193.465 22.110 ;
        RECT 65.000 21.880 165.055 21.975 ;
        POLYGON 165.055 21.975 165.140 21.880 165.055 21.880 ;
        RECT 65.000 21.785 165.140 21.880 ;
        POLYGON 169.655 21.975 169.655 21.875 169.510 21.875 ;
        RECT 169.655 21.875 193.465 21.975 ;
        POLYGON 165.140 21.875 165.220 21.785 165.140 21.785 ;
        POLYGON 169.510 21.875 169.510 21.785 169.375 21.785 ;
        RECT 169.510 21.845 193.465 21.875 ;
        POLYGON 193.465 23.955 194.395 23.955 193.465 21.845 ;
        POLYGON 222.500 23.955 223.020 23.955 223.020 23.550 ;
        RECT 223.020 23.685 266.830 23.955 ;
        POLYGON 266.830 23.955 267.135 23.955 266.830 23.685 ;
        POLYGON 285.525 23.955 285.525 23.685 285.475 23.685 ;
        RECT 285.525 23.685 303.120 23.955 ;
        RECT 223.020 23.550 266.665 23.685 ;
        POLYGON 266.665 23.685 266.830 23.685 266.665 23.550 ;
        POLYGON 285.475 23.685 285.475 23.550 285.450 23.550 ;
        RECT 285.475 23.550 303.120 23.685 ;
        POLYGON 223.020 23.550 223.035 23.550 223.035 23.540 ;
        RECT 223.035 23.540 265.850 23.550 ;
        POLYGON 223.035 23.540 224.120 23.540 224.120 22.755 ;
        RECT 224.120 22.890 265.850 23.540 ;
        POLYGON 265.850 23.550 266.665 23.550 265.850 22.890 ;
        POLYGON 285.450 23.550 285.450 22.890 285.300 22.890 ;
        RECT 285.450 22.890 303.120 23.550 ;
        RECT 224.120 22.755 264.920 22.890 ;
        POLYGON 224.120 22.755 224.295 22.755 224.295 22.635 ;
        RECT 224.295 22.635 264.920 22.755 ;
        POLYGON 224.295 22.635 225.225 22.635 225.225 22.005 ;
        RECT 225.225 22.195 264.920 22.635 ;
        POLYGON 264.920 22.890 265.850 22.890 264.920 22.195 ;
        POLYGON 285.300 22.890 285.300 22.195 285.140 22.195 ;
        RECT 285.300 22.195 303.120 22.890 ;
        RECT 225.225 22.140 264.850 22.195 ;
        POLYGON 264.850 22.195 264.920 22.195 264.850 22.140 ;
        POLYGON 285.140 22.185 285.140 22.140 285.130 22.140 ;
        RECT 285.140 22.140 303.120 22.195 ;
        RECT 225.225 22.005 264.420 22.140 ;
        POLYGON 225.225 22.005 225.480 22.005 225.480 21.845 ;
        RECT 225.480 21.845 264.420 22.005 ;
        POLYGON 264.420 22.140 264.850 22.140 264.420 21.845 ;
        POLYGON 285.130 22.140 285.130 21.855 285.065 21.855 ;
        RECT 285.130 21.855 303.120 22.140 ;
        RECT 169.510 21.785 192.580 21.845 ;
        RECT 65.000 21.680 165.220 21.785 ;
        POLYGON 165.220 21.785 165.310 21.680 165.220 21.680 ;
        POLYGON 169.375 21.785 169.375 21.680 169.225 21.680 ;
        RECT 169.375 21.680 192.580 21.785 ;
        RECT 65.000 21.655 165.310 21.680 ;
        POLYGON 165.310 21.680 165.335 21.655 165.310 21.655 ;
        POLYGON 169.225 21.680 169.225 21.655 169.185 21.655 ;
        RECT 169.225 21.655 192.580 21.680 ;
        RECT 65.000 21.600 165.335 21.655 ;
        POLYGON 165.335 21.655 165.380 21.600 165.335 21.600 ;
        POLYGON 169.185 21.655 169.185 21.600 169.105 21.600 ;
        RECT 169.185 21.600 192.580 21.655 ;
        RECT 65.000 21.440 165.380 21.600 ;
        POLYGON 165.380 21.600 165.520 21.440 165.380 21.440 ;
        POLYGON 169.105 21.600 169.105 21.440 168.875 21.440 ;
        RECT 169.105 21.440 192.580 21.600 ;
        RECT 65.000 21.370 165.520 21.440 ;
        POLYGON 165.520 21.440 165.580 21.370 165.520 21.370 ;
        POLYGON 168.875 21.440 168.875 21.405 168.825 21.405 ;
        RECT 168.875 21.405 192.580 21.440 ;
        POLYGON 168.825 21.405 168.825 21.370 168.770 21.370 ;
        RECT 168.825 21.370 192.580 21.405 ;
        RECT 65.000 21.310 165.580 21.370 ;
        POLYGON 165.580 21.370 165.635 21.310 165.580 21.310 ;
        RECT 65.000 21.270 165.635 21.310 ;
        POLYGON 168.770 21.370 168.770 21.305 168.665 21.305 ;
        RECT 168.770 21.305 192.580 21.370 ;
        POLYGON 165.635 21.305 165.670 21.270 165.635 21.270 ;
        RECT 65.000 21.165 165.670 21.270 ;
        POLYGON 168.665 21.305 168.665 21.265 168.605 21.265 ;
        RECT 168.665 21.265 192.580 21.305 ;
        POLYGON 165.670 21.265 165.760 21.165 165.670 21.165 ;
        POLYGON 168.605 21.265 168.605 21.165 168.445 21.165 ;
        RECT 168.605 21.165 192.580 21.265 ;
        RECT 65.000 21.055 165.760 21.165 ;
        POLYGON 165.760 21.165 165.855 21.055 165.760 21.055 ;
        POLYGON 168.445 21.165 168.445 21.055 168.280 21.055 ;
        RECT 168.445 21.055 192.580 21.165 ;
        RECT 65.000 21.025 165.855 21.055 ;
        POLYGON 165.855 21.055 165.880 21.025 165.855 21.025 ;
        POLYGON 168.280 21.055 168.280 21.025 168.230 21.025 ;
        RECT 168.280 21.025 192.580 21.055 ;
        RECT 65.000 20.740 165.880 21.025 ;
        POLYGON 165.880 21.025 166.130 20.740 165.880 20.740 ;
        RECT 65.000 20.730 166.130 20.740 ;
        POLYGON 168.230 21.025 168.230 20.735 167.770 20.735 ;
        RECT 168.230 20.735 192.580 21.025 ;
        POLYGON 166.130 20.735 166.135 20.730 166.130 20.730 ;
        POLYGON 167.770 20.735 167.770 20.730 167.760 20.730 ;
        RECT 167.770 20.730 192.580 20.735 ;
        RECT 65.000 20.660 166.135 20.730 ;
        POLYGON 166.135 20.730 166.200 20.660 166.135 20.660 ;
        POLYGON 167.760 20.730 167.760 20.660 167.640 20.660 ;
        RECT 167.760 20.660 192.580 20.730 ;
        RECT 65.000 20.600 166.200 20.660 ;
        POLYGON 166.200 20.660 166.255 20.600 166.200 20.600 ;
        POLYGON 167.640 20.660 167.640 20.600 167.535 20.600 ;
        RECT 167.640 20.600 192.580 20.660 ;
        RECT 65.000 20.435 166.255 20.600 ;
        POLYGON 166.255 20.600 166.415 20.435 166.255 20.435 ;
        POLYGON 167.535 20.600 167.535 20.435 167.250 20.435 ;
        RECT 167.535 20.435 192.580 20.600 ;
        RECT 65.000 20.380 166.415 20.435 ;
        POLYGON 166.415 20.435 166.470 20.380 166.415 20.380 ;
        POLYGON 167.250 20.435 167.250 20.405 167.195 20.405 ;
        RECT 167.250 20.405 192.580 20.435 ;
        POLYGON 167.195 20.405 167.195 20.380 167.150 20.380 ;
        RECT 167.195 20.380 192.580 20.405 ;
        RECT 65.000 20.370 166.470 20.380 ;
        POLYGON 166.470 20.380 166.475 20.370 166.470 20.370 ;
        POLYGON 167.150 20.380 167.150 20.370 167.135 20.370 ;
        RECT 167.150 20.370 192.580 20.380 ;
        RECT 65.000 20.290 166.475 20.370 ;
        POLYGON 166.475 20.370 166.555 20.290 166.475 20.290 ;
        POLYGON 167.135 20.370 167.135 20.325 167.055 20.325 ;
        RECT 167.135 20.325 192.580 20.370 ;
        POLYGON 167.055 20.325 167.055 20.290 166.995 20.290 ;
        RECT 167.055 20.290 192.580 20.325 ;
        RECT 65.000 20.245 166.555 20.290 ;
        POLYGON 166.555 20.290 166.595 20.245 166.555 20.245 ;
        POLYGON 166.995 20.290 166.995 20.245 166.920 20.245 ;
        RECT 166.995 20.245 192.580 20.290 ;
        RECT 65.000 20.145 166.595 20.245 ;
        POLYGON 166.595 20.245 166.695 20.145 166.595 20.145 ;
        POLYGON 166.920 20.245 166.920 20.145 166.750 20.145 ;
        RECT 166.920 20.145 192.580 20.245 ;
        RECT 65.000 20.130 166.695 20.145 ;
        POLYGON 166.695 20.145 166.705 20.130 166.695 20.130 ;
        POLYGON 166.750 20.145 166.750 20.130 166.725 20.130 ;
        RECT 166.750 20.130 192.580 20.145 ;
        RECT 65.000 20.125 166.705 20.130 ;
        POLYGON 166.705 20.130 166.710 20.125 166.705 20.125 ;
        POLYGON 166.720 20.130 166.720 20.125 166.715 20.125 ;
        RECT 166.720 20.125 192.580 20.130 ;
        RECT 65.000 20.060 192.580 20.125 ;
        POLYGON 192.580 21.845 193.465 21.845 192.580 20.060 ;
        POLYGON 225.480 21.845 226.360 21.845 226.360 21.300 ;
        RECT 226.360 21.435 263.820 21.845 ;
        POLYGON 263.820 21.845 264.420 21.845 263.820 21.435 ;
        POLYGON 285.065 21.845 285.065 21.435 284.970 21.435 ;
        RECT 285.065 21.435 303.120 21.855 ;
        RECT 226.360 21.300 262.770 21.435 ;
        POLYGON 226.360 21.300 227.075 21.300 227.075 20.890 ;
        RECT 227.075 20.890 262.770 21.300 ;
        POLYGON 227.075 20.890 227.520 20.890 227.520 20.630 ;
        RECT 227.520 20.770 262.770 20.890 ;
        POLYGON 262.770 21.435 263.820 21.435 262.770 20.770 ;
        POLYGON 284.970 21.430 284.970 20.770 284.820 20.770 ;
        RECT 284.970 20.770 303.120 21.435 ;
        RECT 227.520 20.630 261.690 20.770 ;
        POLYGON 227.520 20.630 228.540 20.630 228.540 20.090 ;
        RECT 228.540 20.145 261.690 20.630 ;
        POLYGON 261.690 20.770 262.770 20.770 261.690 20.145 ;
        POLYGON 284.820 20.770 284.820 20.155 284.680 20.155 ;
        RECT 284.820 20.155 303.120 20.770 ;
        RECT 228.540 20.090 261.585 20.145 ;
        POLYGON 261.585 20.145 261.690 20.145 261.585 20.090 ;
        POLYGON 284.680 20.145 284.680 20.090 284.665 20.090 ;
        RECT 284.680 20.090 303.120 20.155 ;
        POLYGON 228.540 20.090 228.600 20.090 228.600 20.060 ;
        RECT 228.600 20.060 261.530 20.090 ;
        POLYGON 261.530 20.090 261.585 20.090 261.530 20.060 ;
        POLYGON 284.665 20.090 284.665 20.070 284.660 20.070 ;
        RECT 284.665 20.070 303.120 20.090 ;
        RECT 65.000 19.770 192.440 20.060 ;
        POLYGON 192.440 20.060 192.580 20.060 192.440 19.770 ;
        POLYGON 228.600 20.060 228.705 20.060 228.705 20.005 ;
        RECT 228.705 20.005 261.170 20.060 ;
        POLYGON 228.705 20.005 229.185 20.005 229.185 19.770 ;
        RECT 229.185 19.870 261.170 20.005 ;
        POLYGON 261.170 20.060 261.530 20.060 261.170 19.870 ;
        POLYGON 284.660 20.060 284.660 19.875 284.615 19.875 ;
        RECT 284.660 19.875 303.120 20.070 ;
        RECT 229.185 19.770 260.960 19.870 ;
        RECT 18.180 12.840 25.870 17.825 ;
        POLYGON 25.870 17.825 27.225 12.840 25.870 12.840 ;
        RECT 65.000 17.740 191.315 19.770 ;
        POLYGON 191.315 19.770 192.440 19.770 191.315 17.740 ;
        POLYGON 229.185 19.770 229.205 19.770 229.205 19.760 ;
        RECT 229.205 19.760 260.960 19.770 ;
        POLYGON 260.960 19.870 261.170 19.870 260.960 19.760 ;
        POLYGON 284.615 19.870 284.615 19.770 284.590 19.770 ;
        RECT 284.615 19.770 303.120 19.875 ;
        POLYGON 229.205 19.760 229.910 19.760 229.910 19.420 ;
        RECT 229.910 19.565 260.585 19.760 ;
        POLYGON 260.585 19.760 260.960 19.760 260.585 19.565 ;
        POLYGON 284.590 19.760 284.590 19.565 284.545 19.565 ;
        RECT 284.590 19.565 303.120 19.770 ;
        RECT 229.910 19.420 259.455 19.565 ;
        POLYGON 229.910 19.420 230.025 19.420 230.025 19.370 ;
        RECT 230.025 19.370 259.455 19.420 ;
        POLYGON 230.025 19.370 231.140 19.370 231.140 18.880 ;
        RECT 231.140 19.025 259.455 19.370 ;
        POLYGON 259.455 19.565 260.585 19.565 259.455 19.025 ;
        POLYGON 284.545 19.560 284.545 19.035 284.425 19.035 ;
        RECT 284.545 19.035 303.120 19.565 ;
        RECT 231.140 18.880 258.295 19.025 ;
        POLYGON 231.140 18.880 232.390 18.880 232.390 18.380 ;
        RECT 232.390 18.525 258.295 18.880 ;
        POLYGON 258.295 19.025 259.455 19.025 258.295 18.525 ;
        POLYGON 284.425 19.025 284.425 18.530 284.310 18.530 ;
        RECT 284.425 18.530 303.120 19.035 ;
        RECT 232.390 18.380 257.660 18.525 ;
        POLYGON 232.390 18.380 233.140 18.380 233.140 18.110 ;
        RECT 233.140 18.280 257.660 18.380 ;
        POLYGON 257.660 18.525 258.295 18.525 257.660 18.280 ;
        POLYGON 284.310 18.525 284.310 18.285 284.255 18.285 ;
        RECT 284.310 18.285 303.120 18.530 ;
        RECT 233.140 18.110 257.115 18.280 ;
        POLYGON 233.140 18.110 233.880 18.110 233.880 17.840 ;
        RECT 233.880 18.070 257.115 18.110 ;
        POLYGON 257.115 18.280 257.660 18.280 257.115 18.070 ;
        POLYGON 284.255 18.280 284.255 18.070 284.205 18.070 ;
        RECT 284.255 18.070 303.120 18.285 ;
        RECT 233.880 17.840 256.270 18.070 ;
        POLYGON 233.880 17.840 234.065 17.840 234.065 17.780 ;
        RECT 234.065 17.780 256.270 17.840 ;
        POLYGON 256.270 18.070 257.115 18.070 256.270 17.780 ;
        POLYGON 284.205 18.065 284.205 17.780 284.140 17.780 ;
        RECT 284.205 17.780 303.120 18.070 ;
        POLYGON 234.065 17.780 234.190 17.780 234.190 17.740 ;
        RECT 234.190 17.740 256.155 17.780 ;
        POLYGON 256.155 17.780 256.270 17.780 256.155 17.740 ;
        POLYGON 284.140 17.780 284.140 17.745 284.130 17.745 ;
        RECT 284.140 17.745 303.120 17.780 ;
        RECT 65.000 15.750 190.095 17.740 ;
        POLYGON 190.095 17.740 191.315 17.740 190.095 15.750 ;
        POLYGON 234.190 17.740 235.275 17.740 235.275 17.395 ;
        RECT 235.275 17.655 255.905 17.740 ;
        POLYGON 255.905 17.740 256.155 17.740 255.905 17.655 ;
        POLYGON 284.130 17.740 284.130 17.655 284.105 17.655 ;
        RECT 284.130 17.655 303.120 17.745 ;
        RECT 235.275 17.395 254.670 17.655 ;
        POLYGON 235.275 17.395 236.410 17.395 236.410 17.085 ;
        RECT 236.410 17.280 254.670 17.395 ;
        POLYGON 254.670 17.655 255.905 17.655 254.670 17.280 ;
        POLYGON 284.105 17.650 284.105 17.280 284.005 17.280 ;
        RECT 284.105 17.280 303.120 17.655 ;
        RECT 236.410 17.185 254.295 17.280 ;
        POLYGON 254.295 17.280 254.670 17.280 254.295 17.185 ;
        POLYGON 284.005 17.280 284.005 17.190 283.980 17.190 ;
        RECT 284.005 17.190 303.120 17.280 ;
        RECT 236.410 17.085 253.405 17.185 ;
        POLYGON 236.410 17.085 236.610 17.085 236.610 17.030 ;
        RECT 236.610 17.030 253.405 17.085 ;
        POLYGON 236.610 17.030 237.940 17.030 237.940 16.735 ;
        RECT 237.940 16.950 253.405 17.030 ;
        POLYGON 253.405 17.185 254.290 17.185 253.405 16.950 ;
        POLYGON 283.980 17.185 283.980 16.950 283.915 16.950 ;
        RECT 283.980 16.950 303.120 17.190 ;
        RECT 237.940 16.735 252.120 16.950 ;
        POLYGON 237.940 16.735 239.300 16.735 239.300 16.510 ;
        RECT 239.300 16.660 252.120 16.735 ;
        POLYGON 252.120 16.950 253.405 16.950 252.120 16.660 ;
        POLYGON 283.915 16.950 283.915 16.660 283.835 16.660 ;
        RECT 283.915 16.660 303.120 16.950 ;
        RECT 239.300 16.510 251.105 16.660 ;
        POLYGON 239.300 16.510 239.835 16.510 239.835 16.445 ;
        RECT 239.835 16.460 251.105 16.510 ;
        POLYGON 251.105 16.660 252.120 16.660 251.105 16.460 ;
        POLYGON 283.835 16.655 283.835 16.460 283.780 16.460 ;
        RECT 283.835 16.460 303.120 16.660 ;
        RECT 239.835 16.445 250.970 16.460 ;
        POLYGON 239.835 16.445 240.745 16.445 240.745 16.340 ;
        RECT 240.745 16.435 250.970 16.445 ;
        POLYGON 250.970 16.460 251.105 16.460 250.970 16.435 ;
        POLYGON 283.780 16.455 283.780 16.435 283.775 16.435 ;
        RECT 283.780 16.435 303.120 16.460 ;
        RECT 240.745 16.340 250.195 16.435 ;
        POLYGON 240.745 16.340 242.310 16.340 242.310 16.215 ;
        RECT 242.310 16.305 250.195 16.340 ;
        POLYGON 250.195 16.435 250.970 16.435 250.195 16.305 ;
        POLYGON 283.775 16.435 283.775 16.305 283.740 16.305 ;
        RECT 283.775 16.305 303.120 16.435 ;
        RECT 242.310 16.215 249.345 16.305 ;
        POLYGON 242.310 16.215 243.400 16.215 243.400 16.160 ;
        RECT 243.400 16.190 249.345 16.215 ;
        POLYGON 249.345 16.305 250.195 16.305 249.345 16.190 ;
        POLYGON 283.740 16.305 283.740 16.195 283.710 16.195 ;
        RECT 283.740 16.195 303.120 16.305 ;
        RECT 243.400 16.160 248.495 16.190 ;
        POLYGON 243.405 16.160 244.040 16.160 244.040 16.130 ;
        RECT 244.040 16.130 248.495 16.160 ;
        POLYGON 244.040 16.130 246.585 16.130 246.585 16.065 ;
        RECT 246.585 16.115 248.495 16.130 ;
        POLYGON 248.495 16.190 249.345 16.190 248.495 16.115 ;
        POLYGON 283.710 16.190 283.710 16.125 283.690 16.125 ;
        RECT 283.710 16.125 303.120 16.195 ;
        RECT 246.585 16.080 247.130 16.115 ;
        POLYGON 247.130 16.115 248.495 16.115 247.130 16.080 ;
        POLYGON 283.690 16.115 283.690 16.085 283.680 16.085 ;
        RECT 283.690 16.085 303.120 16.125 ;
        POLYGON 246.585 16.080 247.120 16.080 246.585 16.065 ;
        POLYGON 283.680 16.080 283.680 16.070 283.675 16.070 ;
        RECT 283.680 16.070 303.120 16.085 ;
        POLYGON 283.675 16.065 283.675 16.050 283.670 16.050 ;
        RECT 283.675 16.050 303.120 16.070 ;
        POLYGON 283.670 16.050 283.670 15.755 283.590 15.755 ;
        RECT 283.670 15.755 303.120 16.050 ;
        RECT 65.000 15.505 189.930 15.750 ;
        POLYGON 189.930 15.750 190.095 15.750 189.930 15.505 ;
        POLYGON 283.590 15.750 283.590 15.505 283.520 15.505 ;
        RECT 283.590 15.505 303.120 15.755 ;
        RECT 65.000 13.810 188.785 15.505 ;
        POLYGON 188.785 15.505 189.930 15.505 188.785 13.810 ;
        POLYGON 283.520 15.500 283.520 13.815 283.060 13.815 ;
        RECT 283.520 13.815 303.120 15.505 ;
        RECT 18.180 12.670 27.225 12.840 ;
        POLYGON 18.180 12.670 20.715 12.670 20.715 4.390 ;
        RECT 20.715 12.115 27.225 12.670 ;
        POLYGON 27.225 12.840 27.420 12.115 27.225 12.115 ;
        RECT 20.715 6.500 27.420 12.115 ;
        POLYGON 27.420 12.115 29.215 6.500 27.420 6.500 ;
        RECT 65.000 11.915 187.385 13.810 ;
        POLYGON 187.385 13.810 188.785 13.810 187.385 11.915 ;
        POLYGON 283.060 13.810 283.060 13.105 282.865 13.105 ;
        RECT 283.060 13.105 303.120 13.815 ;
        POLYGON 282.865 13.105 282.865 12.810 282.785 12.810 ;
        RECT 282.865 12.810 303.120 13.105 ;
        POLYGON 282.785 12.810 282.785 12.490 282.695 12.490 ;
        RECT 282.785 12.490 303.120 12.810 ;
        POLYGON 282.695 12.490 282.695 12.370 282.660 12.370 ;
        RECT 282.695 12.370 303.120 12.490 ;
        POLYGON 282.660 12.370 282.660 12.325 282.645 12.325 ;
        RECT 282.660 12.325 303.120 12.370 ;
        POLYGON 282.645 12.325 282.645 12.305 282.640 12.305 ;
        RECT 282.645 12.305 303.120 12.325 ;
        POLYGON 282.640 12.300 282.640 12.290 282.635 12.290 ;
        RECT 282.640 12.290 303.120 12.305 ;
        POLYGON 282.635 12.290 282.635 12.285 282.630 12.285 ;
        RECT 282.635 12.285 303.120 12.290 ;
        POLYGON 282.630 12.285 282.630 12.260 282.610 12.260 ;
        RECT 282.630 12.260 303.120 12.285 ;
        POLYGON 282.610 12.260 282.610 12.180 282.550 12.180 ;
        RECT 282.610 12.180 303.120 12.260 ;
        POLYGON 282.550 12.180 282.550 12.085 282.475 12.085 ;
        RECT 282.550 12.085 303.120 12.180 ;
        POLYGON 282.475 12.080 282.475 11.975 282.395 11.975 ;
        RECT 282.475 11.975 303.120 12.085 ;
        POLYGON 282.395 11.975 282.395 11.920 282.350 11.920 ;
        RECT 282.395 11.920 303.120 11.975 ;
        RECT 65.000 11.660 187.180 11.915 ;
        POLYGON 187.180 11.915 187.385 11.915 187.180 11.660 ;
        POLYGON 282.350 11.915 282.350 11.910 282.345 11.910 ;
        RECT 282.350 11.910 303.120 11.920 ;
        POLYGON 282.345 11.910 282.345 11.865 282.310 11.865 ;
        RECT 282.345 11.865 303.120 11.910 ;
        POLYGON 282.310 11.865 282.310 11.665 282.155 11.665 ;
        RECT 282.310 11.665 303.120 11.865 ;
        RECT 65.000 10.075 185.900 11.660 ;
        POLYGON 185.900 11.660 187.180 11.660 185.900 10.075 ;
        POLYGON 282.155 11.660 282.155 11.205 281.805 11.205 ;
        RECT 282.155 11.205 303.120 11.665 ;
        POLYGON 281.805 11.205 281.805 10.725 281.405 10.725 ;
        RECT 281.805 10.725 303.120 11.205 ;
        POLYGON 281.405 10.725 281.405 10.075 280.860 10.075 ;
        RECT 281.405 10.075 303.120 10.725 ;
        RECT 65.000 8.305 184.335 10.075 ;
        POLYGON 184.335 10.075 185.900 10.075 184.335 8.305 ;
        POLYGON 280.860 10.075 280.860 10.070 280.855 10.070 ;
        RECT 280.860 10.070 303.120 10.075 ;
        POLYGON 280.855 10.070 280.855 9.380 280.275 9.380 ;
        RECT 280.855 9.380 303.120 10.070 ;
        POLYGON 280.275 9.380 280.275 9.300 280.205 9.300 ;
        RECT 280.275 9.300 303.120 9.380 ;
        POLYGON 280.205 9.300 280.205 8.305 279.295 8.305 ;
        RECT 280.205 8.305 303.120 9.300 ;
        RECT 65.000 8.290 184.325 8.305 ;
        POLYGON 184.325 8.305 184.335 8.305 184.325 8.290 ;
        POLYGON 279.295 8.300 279.295 8.290 279.285 8.290 ;
        RECT 279.295 8.290 303.120 8.305 ;
        RECT 65.000 7.640 182.665 8.290 ;
        RECT 20.715 4.390 29.215 6.500 ;
        POLYGON 20.715 4.390 22.040 4.390 22.040 0.835 ;
        RECT 22.040 1.195 29.215 4.390 ;
        POLYGON 29.215 6.500 31.170 1.195 29.215 1.195 ;
        RECT 65.000 5.000 85.000 7.640 ;
        POLYGON 85.000 7.640 86.510 7.640 86.510 6.500 ;
        RECT 86.510 6.565 182.665 7.640 ;
        POLYGON 182.665 8.290 184.325 8.290 182.665 6.565 ;
        POLYGON 279.285 8.290 279.285 7.935 278.960 7.935 ;
        RECT 279.285 7.935 303.120 8.290 ;
        POLYGON 278.960 7.935 278.960 7.715 278.760 7.715 ;
        RECT 278.960 7.715 303.120 7.935 ;
        POLYGON 278.760 7.715 278.760 7.620 278.675 7.620 ;
        RECT 278.760 7.620 303.120 7.715 ;
        POLYGON 278.675 7.620 278.675 6.855 277.915 6.855 ;
        RECT 278.675 6.855 303.120 7.620 ;
        POLYGON 277.915 6.855 277.915 6.565 277.625 6.565 ;
        RECT 277.915 6.565 303.120 6.855 ;
        RECT 86.510 6.500 182.420 6.565 ;
        POLYGON 86.510 6.500 87.615 6.500 87.615 5.665 ;
        RECT 87.615 6.330 182.420 6.500 ;
        POLYGON 182.420 6.565 182.665 6.565 182.420 6.330 ;
        POLYGON 277.625 6.565 277.625 6.330 277.390 6.330 ;
        RECT 277.625 6.330 303.120 6.565 ;
        RECT 87.615 6.240 182.325 6.330 ;
        POLYGON 182.325 6.330 182.420 6.330 182.325 6.240 ;
        POLYGON 277.390 6.330 277.390 6.240 277.305 6.240 ;
        RECT 277.390 6.240 303.120 6.330 ;
        RECT 87.615 6.110 182.195 6.240 ;
        POLYGON 182.195 6.240 182.325 6.240 182.195 6.110 ;
        POLYGON 277.305 6.240 277.305 6.110 277.175 6.110 ;
        RECT 277.305 6.110 303.120 6.240 ;
        RECT 87.615 6.060 182.165 6.110 ;
        POLYGON 182.165 6.110 182.195 6.110 182.165 6.085 ;
        POLYGON 182.165 6.085 182.195 6.060 182.165 6.060 ;
        POLYGON 277.175 6.110 277.175 6.060 277.125 6.060 ;
        RECT 277.175 6.060 303.120 6.110 ;
        RECT 87.615 6.055 182.200 6.060 ;
        POLYGON 182.200 6.060 182.210 6.055 182.200 6.055 ;
        POLYGON 277.125 6.060 277.125 6.055 277.120 6.055 ;
        RECT 277.125 6.055 303.120 6.060 ;
        RECT 87.615 6.045 182.210 6.055 ;
        POLYGON 182.210 6.055 182.220 6.045 182.210 6.045 ;
        POLYGON 277.120 6.055 277.120 6.045 277.110 6.045 ;
        RECT 277.120 6.045 303.120 6.055 ;
        RECT 87.615 6.040 182.220 6.045 ;
        POLYGON 182.220 6.045 182.230 6.040 182.220 6.040 ;
        POLYGON 277.110 6.045 277.110 6.040 277.105 6.040 ;
        RECT 277.110 6.040 303.120 6.045 ;
        RECT 87.615 6.020 182.230 6.040 ;
        POLYGON 182.230 6.040 182.255 6.020 182.230 6.020 ;
        POLYGON 277.105 6.040 277.105 6.020 277.085 6.020 ;
        RECT 277.105 6.020 303.120 6.040 ;
        RECT 87.615 6.015 182.255 6.020 ;
        POLYGON 182.255 6.020 182.265 6.015 182.255 6.015 ;
        POLYGON 277.085 6.020 277.085 6.015 277.080 6.015 ;
        RECT 277.085 6.015 303.120 6.020 ;
        RECT 87.615 5.975 182.270 6.015 ;
        POLYGON 182.270 6.015 182.325 5.975 182.270 5.975 ;
        POLYGON 277.080 6.015 277.080 5.975 277.040 5.975 ;
        RECT 277.080 5.975 303.120 6.015 ;
        RECT 87.615 5.905 182.325 5.975 ;
        POLYGON 182.325 5.975 182.420 5.905 182.325 5.905 ;
        POLYGON 277.040 5.975 277.040 5.940 277.005 5.940 ;
        RECT 277.040 5.940 303.120 5.975 ;
        POLYGON 277.005 5.940 277.005 5.905 276.965 5.905 ;
        RECT 277.005 5.905 303.120 5.940 ;
        RECT 87.615 5.780 182.420 5.905 ;
        POLYGON 182.420 5.905 182.600 5.780 182.420 5.780 ;
        POLYGON 276.965 5.905 276.965 5.840 276.895 5.840 ;
        RECT 276.965 5.840 303.120 5.905 ;
        POLYGON 276.895 5.840 276.895 5.780 276.830 5.780 ;
        RECT 276.895 5.780 303.120 5.840 ;
        RECT 87.615 5.665 182.600 5.780 ;
        POLYGON 87.615 5.665 88.450 5.665 88.450 5.100 ;
        RECT 88.450 5.350 182.600 5.665 ;
        POLYGON 182.600 5.780 183.230 5.350 182.600 5.350 ;
        POLYGON 276.830 5.780 276.830 5.505 276.535 5.505 ;
        RECT 276.830 5.505 303.120 5.780 ;
        POLYGON 276.535 5.505 276.535 5.350 276.370 5.350 ;
        RECT 276.535 5.350 303.120 5.505 ;
        RECT 88.450 5.155 183.230 5.350 ;
        POLYGON 183.230 5.350 183.520 5.155 183.230 5.155 ;
        POLYGON 276.370 5.350 276.370 5.155 276.160 5.155 ;
        RECT 276.370 5.155 303.120 5.350 ;
        RECT 88.450 5.100 183.520 5.155 ;
        POLYGON 88.450 5.100 88.595 5.100 88.595 5.000 ;
        RECT 88.595 5.000 183.520 5.100 ;
        POLYGON 88.595 5.000 92.160 5.000 92.160 2.605 ;
        RECT 92.160 4.900 183.520 5.000 ;
        POLYGON 183.520 5.155 183.895 4.900 183.520 4.900 ;
        POLYGON 276.160 5.155 276.160 5.115 276.115 5.115 ;
        RECT 276.160 5.115 303.120 5.155 ;
        POLYGON 276.115 5.115 276.115 4.900 275.885 4.900 ;
        RECT 276.115 4.900 303.120 5.115 ;
        RECT 92.160 3.535 183.895 4.900 ;
        POLYGON 183.895 4.900 185.905 3.535 183.895 3.535 ;
        POLYGON 275.885 4.900 275.885 4.670 275.635 4.670 ;
        RECT 275.885 4.670 303.120 4.900 ;
        POLYGON 275.635 4.670 275.635 4.330 275.265 4.330 ;
        RECT 275.635 4.330 303.120 4.670 ;
        POLYGON 275.265 4.330 275.265 4.185 275.095 4.185 ;
        RECT 275.265 4.185 303.120 4.330 ;
        POLYGON 275.095 4.185 275.095 3.675 274.500 3.675 ;
        RECT 275.095 3.675 303.120 4.185 ;
        POLYGON 274.500 3.675 274.500 3.535 274.335 3.535 ;
        RECT 274.500 3.535 303.120 3.675 ;
        RECT 92.160 3.300 185.905 3.535 ;
        POLYGON 185.905 3.535 186.255 3.300 185.905 3.300 ;
        POLYGON 274.335 3.535 274.335 3.300 274.060 3.300 ;
        RECT 274.335 3.300 303.120 3.535 ;
        RECT 92.160 2.995 186.255 3.300 ;
        POLYGON 186.255 3.300 186.705 2.995 186.255 2.995 ;
        POLYGON 274.060 3.300 274.060 3.115 273.840 3.115 ;
        RECT 274.060 3.115 303.120 3.300 ;
        POLYGON 273.840 3.115 273.840 2.995 273.700 2.995 ;
        RECT 273.840 2.995 303.120 3.115 ;
        RECT 92.160 2.990 186.705 2.995 ;
        POLYGON 186.705 2.995 186.710 2.990 186.705 2.990 ;
        POLYGON 273.700 2.995 273.700 2.990 273.695 2.990 ;
        RECT 273.700 2.990 303.120 2.995 ;
        RECT 92.160 2.710 186.710 2.990 ;
        POLYGON 186.710 2.990 187.175 2.710 186.710 2.710 ;
        POLYGON 273.695 2.990 273.695 2.855 273.535 2.855 ;
        RECT 273.695 2.855 303.120 2.990 ;
        POLYGON 273.535 2.855 273.535 2.795 273.460 2.795 ;
        RECT 273.535 2.795 303.120 2.855 ;
        POLYGON 273.460 2.795 273.460 2.710 273.350 2.710 ;
        RECT 273.460 2.710 303.120 2.795 ;
        RECT 92.160 2.615 187.175 2.710 ;
        POLYGON 187.175 2.710 187.335 2.615 187.175 2.615 ;
        POLYGON 273.350 2.710 273.350 2.615 273.230 2.615 ;
        RECT 273.350 2.615 303.120 2.710 ;
        RECT 92.160 2.605 187.335 2.615 ;
        POLYGON 92.160 2.605 92.270 2.605 92.270 2.540 ;
        RECT 92.270 2.540 187.335 2.605 ;
        POLYGON 92.270 2.540 94.525 2.540 94.525 1.195 ;
        RECT 94.525 1.770 187.335 2.540 ;
        POLYGON 187.335 2.615 188.725 1.770 187.335 1.770 ;
        POLYGON 273.230 2.615 273.230 2.530 273.120 2.530 ;
        RECT 273.230 2.530 303.120 2.615 ;
        POLYGON 273.120 2.530 273.120 1.915 272.340 1.915 ;
        RECT 273.120 1.915 303.120 2.530 ;
        POLYGON 272.340 1.915 272.340 1.770 272.155 1.770 ;
        RECT 272.340 1.770 303.120 1.915 ;
        RECT 94.525 1.195 188.725 1.770 ;
        RECT 22.040 0.980 31.170 1.195 ;
        POLYGON 31.170 1.195 31.250 0.980 31.170 0.980 ;
        POLYGON 94.525 1.195 94.885 1.195 94.885 0.980 ;
        RECT 94.885 1.180 188.725 1.195 ;
        POLYGON 188.725 1.770 189.700 1.180 188.725 1.180 ;
        POLYGON 272.155 1.770 272.155 1.335 271.595 1.335 ;
        RECT 272.155 1.335 303.120 1.770 ;
        POLYGON 271.595 1.335 271.595 1.260 271.490 1.260 ;
        RECT 271.595 1.260 303.120 1.335 ;
        POLYGON 271.490 1.260 271.490 1.180 271.380 1.180 ;
        RECT 271.490 1.180 303.120 1.260 ;
        RECT 94.885 0.980 189.700 1.180 ;
        RECT 22.040 0.835 31.250 0.980 ;
        POLYGON 22.040 0.835 22.195 0.835 22.195 0.435 ;
        RECT 22.195 0.435 31.250 0.835 ;
        POLYGON 22.195 0.435 22.355 0.435 22.355 0.000 ;
        RECT 22.355 0.000 31.250 0.435 ;
        POLYGON 31.250 0.980 31.660 0.000 31.250 0.000 ;
        POLYGON 94.885 0.980 96.205 0.980 96.205 0.195 ;
        RECT 96.205 0.955 189.700 0.980 ;
        POLYGON 189.700 1.180 190.070 0.955 189.700 0.955 ;
        POLYGON 271.380 1.180 271.380 0.955 271.065 0.955 ;
        RECT 271.380 0.955 303.120 1.180 ;
        RECT 96.205 0.455 190.070 0.955 ;
        POLYGON 190.070 0.955 190.900 0.455 190.070 0.455 ;
        POLYGON 271.065 0.955 271.065 0.610 270.585 0.610 ;
        RECT 271.065 0.610 303.120 0.955 ;
        POLYGON 270.585 0.610 270.585 0.455 270.370 0.455 ;
        RECT 270.585 0.455 303.120 0.610 ;
        RECT 96.205 0.340 190.900 0.455 ;
        POLYGON 190.900 0.455 191.090 0.340 190.900 0.340 ;
        POLYGON 270.370 0.455 270.370 0.340 270.210 0.340 ;
        RECT 270.370 0.340 303.120 0.455 ;
        RECT 96.205 0.320 191.090 0.340 ;
        POLYGON 191.090 0.340 191.125 0.320 191.090 0.320 ;
        POLYGON 270.210 0.340 270.210 0.320 270.180 0.320 ;
        RECT 270.210 0.320 303.120 0.340 ;
        RECT 96.205 0.310 191.125 0.320 ;
        POLYGON 191.125 0.320 191.145 0.310 191.125 0.310 ;
        POLYGON 270.180 0.320 270.180 0.310 270.165 0.310 ;
        RECT 270.180 0.310 303.120 0.320 ;
        RECT 96.205 0.245 191.145 0.310 ;
        POLYGON 191.145 0.310 191.270 0.245 191.145 0.245 ;
        POLYGON 270.165 0.310 270.165 0.245 270.075 0.245 ;
        RECT 270.165 0.245 303.120 0.310 ;
        RECT 96.205 0.195 191.270 0.245 ;
        POLYGON 96.205 0.195 96.535 0.195 96.535 0.000 ;
        RECT 96.535 0.000 191.270 0.195 ;
        POLYGON 191.270 0.245 191.725 0.000 191.270 0.000 ;
        POLYGON 270.075 0.245 270.075 0.000 269.735 0.000 ;
        RECT 270.075 0.000 303.120 0.245 ;
      LAYER met4 ;
        RECT 0.200 0.000 1.800 750.000 ;
        RECT 5.000 60.000 25.000 70.000 ;
        RECT 85.000 30.000 105.000 40.000 ;
        RECT 85.000 5.000 105.000 25.000 ;
        RECT 298.200 0.000 299.800 750.000 ;
  END
END Art
END LIBRARY

