magic
tech sky130A
magscale 1 2
timestamp 1683882479
<< obsli1 >>
rect 1104 2159 58880 39729
<< obsm1 >>
rect 934 892 58880 41132
<< metal2 >>
rect 3882 41200 3938 42000
rect 11334 41200 11390 42000
rect 18786 41200 18842 42000
rect 26238 41200 26294 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48594 41200 48650 42000
rect 56046 41200 56102 42000
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57978 0 58034 800
<< obsm2 >>
rect 938 41144 3826 41200
rect 3994 41144 11278 41200
rect 11446 41144 18730 41200
rect 18898 41144 26182 41200
rect 26350 41144 33634 41200
rect 33802 41144 41086 41200
rect 41254 41144 48538 41200
rect 48706 41144 55990 41200
rect 56158 41144 58032 41200
rect 938 856 58032 41144
rect 938 711 1802 856
rect 1970 711 2262 856
rect 2430 711 2722 856
rect 2890 711 3182 856
rect 3350 711 3642 856
rect 3810 711 4102 856
rect 4270 711 4562 856
rect 4730 711 5022 856
rect 5190 711 5482 856
rect 5650 711 5942 856
rect 6110 711 6402 856
rect 6570 711 6862 856
rect 7030 711 7322 856
rect 7490 711 7782 856
rect 7950 711 8242 856
rect 8410 711 8702 856
rect 8870 711 9162 856
rect 9330 711 9622 856
rect 9790 711 10082 856
rect 10250 711 10542 856
rect 10710 711 11002 856
rect 11170 711 11462 856
rect 11630 711 11922 856
rect 12090 711 12382 856
rect 12550 711 12842 856
rect 13010 711 13302 856
rect 13470 711 13762 856
rect 13930 711 14222 856
rect 14390 711 14682 856
rect 14850 711 15142 856
rect 15310 711 15602 856
rect 15770 711 16062 856
rect 16230 711 16522 856
rect 16690 711 16982 856
rect 17150 711 17442 856
rect 17610 711 17902 856
rect 18070 711 18362 856
rect 18530 711 18822 856
rect 18990 711 19282 856
rect 19450 711 19742 856
rect 19910 711 20202 856
rect 20370 711 20662 856
rect 20830 711 21122 856
rect 21290 711 21582 856
rect 21750 711 22042 856
rect 22210 711 22502 856
rect 22670 711 22962 856
rect 23130 711 23422 856
rect 23590 711 23882 856
rect 24050 711 24342 856
rect 24510 711 24802 856
rect 24970 711 25262 856
rect 25430 711 25722 856
rect 25890 711 26182 856
rect 26350 711 26642 856
rect 26810 711 27102 856
rect 27270 711 27562 856
rect 27730 711 28022 856
rect 28190 711 28482 856
rect 28650 711 28942 856
rect 29110 711 29402 856
rect 29570 711 29862 856
rect 30030 711 30322 856
rect 30490 711 30782 856
rect 30950 711 31242 856
rect 31410 711 31702 856
rect 31870 711 32162 856
rect 32330 711 32622 856
rect 32790 711 33082 856
rect 33250 711 33542 856
rect 33710 711 34002 856
rect 34170 711 34462 856
rect 34630 711 34922 856
rect 35090 711 35382 856
rect 35550 711 35842 856
rect 36010 711 36302 856
rect 36470 711 36762 856
rect 36930 711 37222 856
rect 37390 711 37682 856
rect 37850 711 38142 856
rect 38310 711 38602 856
rect 38770 711 39062 856
rect 39230 711 39522 856
rect 39690 711 39982 856
rect 40150 711 40442 856
rect 40610 711 40902 856
rect 41070 711 41362 856
rect 41530 711 41822 856
rect 41990 711 42282 856
rect 42450 711 42742 856
rect 42910 711 43202 856
rect 43370 711 43662 856
rect 43830 711 44122 856
rect 44290 711 44582 856
rect 44750 711 45042 856
rect 45210 711 45502 856
rect 45670 711 45962 856
rect 46130 711 46422 856
rect 46590 711 46882 856
rect 47050 711 47342 856
rect 47510 711 47802 856
rect 47970 711 48262 856
rect 48430 711 48722 856
rect 48890 711 49182 856
rect 49350 711 49642 856
rect 49810 711 50102 856
rect 50270 711 50562 856
rect 50730 711 51022 856
rect 51190 711 51482 856
rect 51650 711 51942 856
rect 52110 711 52402 856
rect 52570 711 52862 856
rect 53030 711 53322 856
rect 53490 711 53782 856
rect 53950 711 54242 856
rect 54410 711 54702 856
rect 54870 711 55162 856
rect 55330 711 55622 856
rect 55790 711 56082 856
rect 56250 711 56542 856
rect 56710 711 57002 856
rect 57170 711 57462 856
rect 57630 711 57922 856
<< metal3 >>
rect 0 41080 800 41200
rect 0 40672 800 40792
rect 0 40264 800 40384
rect 0 39856 800 39976
rect 0 39448 800 39568
rect 0 39040 800 39160
rect 0 38632 800 38752
rect 0 38224 800 38344
rect 0 37816 800 37936
rect 0 37408 800 37528
rect 0 37000 800 37120
rect 0 36592 800 36712
rect 0 36184 800 36304
rect 0 35776 800 35896
rect 0 35368 800 35488
rect 0 34960 800 35080
rect 0 34552 800 34672
rect 0 34144 800 34264
rect 0 33736 800 33856
rect 0 33328 800 33448
rect 0 32920 800 33040
rect 0 32512 800 32632
rect 0 32104 800 32224
rect 0 31696 800 31816
rect 0 31288 800 31408
rect 0 30880 800 31000
rect 0 30472 800 30592
rect 0 30064 800 30184
rect 0 29656 800 29776
rect 0 29248 800 29368
rect 0 28840 800 28960
rect 0 28432 800 28552
rect 0 28024 800 28144
rect 0 27616 800 27736
rect 0 27208 800 27328
rect 0 26800 800 26920
rect 0 26392 800 26512
rect 0 25984 800 26104
rect 0 25576 800 25696
rect 0 25168 800 25288
rect 0 24760 800 24880
rect 0 24352 800 24472
rect 0 23944 800 24064
rect 0 23536 800 23656
rect 0 23128 800 23248
rect 0 22720 800 22840
rect 0 22312 800 22432
rect 0 21904 800 22024
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 0 20680 800 20800
rect 0 20272 800 20392
rect 0 19864 800 19984
rect 0 19456 800 19576
rect 0 19048 800 19168
rect 0 18640 800 18760
rect 0 18232 800 18352
rect 0 17824 800 17944
rect 0 17416 800 17536
rect 0 17008 800 17128
rect 0 16600 800 16720
rect 0 16192 800 16312
rect 0 15784 800 15904
rect 0 15376 800 15496
rect 0 14968 800 15088
rect 0 14560 800 14680
rect 0 14152 800 14272
rect 0 13744 800 13864
rect 0 13336 800 13456
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 12112 800 12232
rect 0 11704 800 11824
rect 0 11296 800 11416
rect 0 10888 800 11008
rect 0 10480 800 10600
rect 0 10072 800 10192
rect 0 9664 800 9784
rect 0 9256 800 9376
rect 0 8848 800 8968
rect 0 8440 800 8560
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6808 800 6928
rect 0 6400 800 6520
rect 0 5992 800 6112
rect 0 5584 800 5704
rect 0 5176 800 5296
rect 0 4768 800 4888
rect 0 4360 800 4480
rect 0 3952 800 4072
rect 0 3544 800 3664
rect 0 3136 800 3256
rect 0 2728 800 2848
rect 0 2320 800 2440
rect 0 1912 800 2032
rect 0 1504 800 1624
rect 0 1096 800 1216
rect 0 688 800 808
<< obsm3 >>
rect 880 41000 50606 41173
rect 800 40872 50606 41000
rect 880 40592 50606 40872
rect 800 40464 50606 40592
rect 880 40184 50606 40464
rect 800 40056 50606 40184
rect 880 39776 50606 40056
rect 800 39648 50606 39776
rect 880 39368 50606 39648
rect 800 39240 50606 39368
rect 880 38960 50606 39240
rect 800 38832 50606 38960
rect 880 38552 50606 38832
rect 800 38424 50606 38552
rect 880 38144 50606 38424
rect 800 38016 50606 38144
rect 880 37736 50606 38016
rect 800 37608 50606 37736
rect 880 37328 50606 37608
rect 800 37200 50606 37328
rect 880 36920 50606 37200
rect 800 36792 50606 36920
rect 880 36512 50606 36792
rect 800 36384 50606 36512
rect 880 36104 50606 36384
rect 800 35976 50606 36104
rect 880 35696 50606 35976
rect 800 35568 50606 35696
rect 880 35288 50606 35568
rect 800 35160 50606 35288
rect 880 34880 50606 35160
rect 800 34752 50606 34880
rect 880 34472 50606 34752
rect 800 34344 50606 34472
rect 880 34064 50606 34344
rect 800 33936 50606 34064
rect 880 33656 50606 33936
rect 800 33528 50606 33656
rect 880 33248 50606 33528
rect 800 33120 50606 33248
rect 880 32840 50606 33120
rect 800 32712 50606 32840
rect 880 32432 50606 32712
rect 800 32304 50606 32432
rect 880 32024 50606 32304
rect 800 31896 50606 32024
rect 880 31616 50606 31896
rect 800 31488 50606 31616
rect 880 31208 50606 31488
rect 800 31080 50606 31208
rect 880 30800 50606 31080
rect 800 30672 50606 30800
rect 880 30392 50606 30672
rect 800 30264 50606 30392
rect 880 29984 50606 30264
rect 800 29856 50606 29984
rect 880 29576 50606 29856
rect 800 29448 50606 29576
rect 880 29168 50606 29448
rect 800 29040 50606 29168
rect 880 28760 50606 29040
rect 800 28632 50606 28760
rect 880 28352 50606 28632
rect 800 28224 50606 28352
rect 880 27944 50606 28224
rect 800 27816 50606 27944
rect 880 27536 50606 27816
rect 800 27408 50606 27536
rect 880 27128 50606 27408
rect 800 27000 50606 27128
rect 880 26720 50606 27000
rect 800 26592 50606 26720
rect 880 26312 50606 26592
rect 800 26184 50606 26312
rect 880 25904 50606 26184
rect 800 25776 50606 25904
rect 880 25496 50606 25776
rect 800 25368 50606 25496
rect 880 25088 50606 25368
rect 800 24960 50606 25088
rect 880 24680 50606 24960
rect 800 24552 50606 24680
rect 880 24272 50606 24552
rect 800 24144 50606 24272
rect 880 23864 50606 24144
rect 800 23736 50606 23864
rect 880 23456 50606 23736
rect 800 23328 50606 23456
rect 880 23048 50606 23328
rect 800 22920 50606 23048
rect 880 22640 50606 22920
rect 800 22512 50606 22640
rect 880 22232 50606 22512
rect 800 22104 50606 22232
rect 880 21824 50606 22104
rect 800 21696 50606 21824
rect 880 21416 50606 21696
rect 800 21288 50606 21416
rect 880 21008 50606 21288
rect 800 20880 50606 21008
rect 880 20600 50606 20880
rect 800 20472 50606 20600
rect 880 20192 50606 20472
rect 800 20064 50606 20192
rect 880 19784 50606 20064
rect 800 19656 50606 19784
rect 880 19376 50606 19656
rect 800 19248 50606 19376
rect 880 18968 50606 19248
rect 800 18840 50606 18968
rect 880 18560 50606 18840
rect 800 18432 50606 18560
rect 880 18152 50606 18432
rect 800 18024 50606 18152
rect 880 17744 50606 18024
rect 800 17616 50606 17744
rect 880 17336 50606 17616
rect 800 17208 50606 17336
rect 880 16928 50606 17208
rect 800 16800 50606 16928
rect 880 16520 50606 16800
rect 800 16392 50606 16520
rect 880 16112 50606 16392
rect 800 15984 50606 16112
rect 880 15704 50606 15984
rect 800 15576 50606 15704
rect 880 15296 50606 15576
rect 800 15168 50606 15296
rect 880 14888 50606 15168
rect 800 14760 50606 14888
rect 880 14480 50606 14760
rect 800 14352 50606 14480
rect 880 14072 50606 14352
rect 800 13944 50606 14072
rect 880 13664 50606 13944
rect 800 13536 50606 13664
rect 880 13256 50606 13536
rect 800 13128 50606 13256
rect 880 12848 50606 13128
rect 800 12720 50606 12848
rect 880 12440 50606 12720
rect 800 12312 50606 12440
rect 880 12032 50606 12312
rect 800 11904 50606 12032
rect 880 11624 50606 11904
rect 800 11496 50606 11624
rect 880 11216 50606 11496
rect 800 11088 50606 11216
rect 880 10808 50606 11088
rect 800 10680 50606 10808
rect 880 10400 50606 10680
rect 800 10272 50606 10400
rect 880 9992 50606 10272
rect 800 9864 50606 9992
rect 880 9584 50606 9864
rect 800 9456 50606 9584
rect 880 9176 50606 9456
rect 800 9048 50606 9176
rect 880 8768 50606 9048
rect 800 8640 50606 8768
rect 880 8360 50606 8640
rect 800 8232 50606 8360
rect 880 7952 50606 8232
rect 800 7824 50606 7952
rect 880 7544 50606 7824
rect 800 7416 50606 7544
rect 880 7136 50606 7416
rect 800 7008 50606 7136
rect 880 6728 50606 7008
rect 800 6600 50606 6728
rect 880 6320 50606 6600
rect 800 6192 50606 6320
rect 880 5912 50606 6192
rect 800 5784 50606 5912
rect 880 5504 50606 5784
rect 800 5376 50606 5504
rect 880 5096 50606 5376
rect 800 4968 50606 5096
rect 880 4688 50606 4968
rect 800 4560 50606 4688
rect 880 4280 50606 4560
rect 800 4152 50606 4280
rect 880 3872 50606 4152
rect 800 3744 50606 3872
rect 880 3464 50606 3744
rect 800 3336 50606 3464
rect 880 3056 50606 3336
rect 800 2928 50606 3056
rect 880 2648 50606 2928
rect 800 2520 50606 2648
rect 880 2240 50606 2520
rect 800 2112 50606 2240
rect 880 1832 50606 2112
rect 800 1704 50606 1832
rect 880 1424 50606 1704
rect 800 1296 50606 1424
rect 880 1016 50606 1296
rect 800 888 50606 1016
rect 880 715 50606 888
<< metal4 >>
rect 4208 2128 4528 39760
rect 19568 2128 19888 39760
rect 34928 2128 35248 39760
rect 50288 2128 50608 39760
<< labels >>
rlabel metal2 s 3882 41200 3938 42000 6 flash_csb
port 1 nsew signal output
rlabel metal2 s 11334 41200 11390 42000 6 flash_io0_read
port 2 nsew signal input
rlabel metal2 s 18786 41200 18842 42000 6 flash_io0_we
port 3 nsew signal output
rlabel metal2 s 26238 41200 26294 42000 6 flash_io0_write
port 4 nsew signal output
rlabel metal2 s 33690 41200 33746 42000 6 flash_io1_read
port 5 nsew signal input
rlabel metal2 s 41142 41200 41198 42000 6 flash_io1_we
port 6 nsew signal output
rlabel metal2 s 48594 41200 48650 42000 6 flash_io1_write
port 7 nsew signal output
rlabel metal2 s 56046 41200 56102 42000 6 flash_sck
port 8 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 sram_addr0[0]
port 9 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 sram_addr0[1]
port 10 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 sram_addr0[2]
port 11 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 sram_addr0[3]
port 12 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 sram_addr0[4]
port 13 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 sram_addr0[5]
port 14 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 sram_addr0[6]
port 15 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 sram_addr0[7]
port 16 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 sram_addr0[8]
port 17 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 sram_addr1[0]
port 18 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 sram_addr1[1]
port 19 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 sram_addr1[2]
port 20 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 sram_addr1[3]
port 21 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 sram_addr1[4]
port 22 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 sram_addr1[5]
port 23 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 sram_addr1[6]
port 24 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 sram_addr1[7]
port 25 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 sram_addr1[8]
port 26 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 sram_clk0
port 27 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 sram_clk1
port 28 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 sram_csb0
port 29 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 sram_csb1
port 30 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 sram_din0[0]
port 31 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 sram_din0[10]
port 32 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 33 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 34 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 sram_din0[13]
port 35 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 sram_din0[14]
port 36 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 sram_din0[15]
port 37 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 sram_din0[16]
port 38 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 sram_din0[17]
port 39 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 sram_din0[18]
port 40 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 sram_din0[19]
port 41 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 sram_din0[1]
port 42 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 sram_din0[20]
port 43 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 sram_din0[21]
port 44 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 sram_din0[22]
port 45 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 sram_din0[23]
port 46 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 sram_din0[24]
port 47 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 sram_din0[25]
port 48 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 sram_din0[26]
port 49 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 sram_din0[27]
port 50 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 sram_din0[28]
port 51 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 sram_din0[29]
port 52 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 sram_din0[2]
port 53 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 sram_din0[30]
port 54 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 sram_din0[31]
port 55 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 sram_din0[3]
port 56 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 sram_din0[4]
port 57 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 sram_din0[5]
port 58 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 sram_din0[6]
port 59 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 sram_din0[7]
port 60 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 sram_din0[8]
port 61 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 sram_din0[9]
port 62 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 sram_dout0[0]
port 63 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 sram_dout0[10]
port 64 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 65 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 sram_dout0[12]
port 66 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 sram_dout0[13]
port 67 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 sram_dout0[14]
port 68 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 sram_dout0[15]
port 69 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 sram_dout0[16]
port 70 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 sram_dout0[17]
port 71 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 sram_dout0[18]
port 72 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 sram_dout0[19]
port 73 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 sram_dout0[1]
port 74 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 sram_dout0[20]
port 75 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 sram_dout0[21]
port 76 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 sram_dout0[22]
port 77 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout0[23]
port 78 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 sram_dout0[24]
port 79 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 sram_dout0[25]
port 80 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 sram_dout0[26]
port 81 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 sram_dout0[27]
port 82 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 sram_dout0[28]
port 83 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[29]
port 84 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 sram_dout0[2]
port 85 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 sram_dout0[30]
port 86 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 sram_dout0[31]
port 87 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 sram_dout0[3]
port 88 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 sram_dout0[4]
port 89 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 sram_dout0[5]
port 90 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 sram_dout0[6]
port 91 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 sram_dout0[7]
port 92 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 sram_dout0[8]
port 93 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 sram_dout0[9]
port 94 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 sram_dout1[0]
port 95 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 sram_dout1[10]
port 96 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 97 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 sram_dout1[12]
port 98 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 sram_dout1[13]
port 99 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 sram_dout1[14]
port 100 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 sram_dout1[15]
port 101 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 sram_dout1[16]
port 102 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout1[17]
port 103 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 sram_dout1[18]
port 104 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 sram_dout1[19]
port 105 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 sram_dout1[1]
port 106 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 sram_dout1[20]
port 107 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 sram_dout1[21]
port 108 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 sram_dout1[22]
port 109 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 sram_dout1[23]
port 110 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 sram_dout1[24]
port 111 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 sram_dout1[25]
port 112 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 sram_dout1[26]
port 113 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 sram_dout1[27]
port 114 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[28]
port 115 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[29]
port 116 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 sram_dout1[2]
port 117 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 sram_dout1[30]
port 118 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 sram_dout1[31]
port 119 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 sram_dout1[3]
port 120 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 sram_dout1[4]
port 121 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 sram_dout1[5]
port 122 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 sram_dout1[6]
port 123 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 sram_dout1[7]
port 124 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 sram_dout1[8]
port 125 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 sram_dout1[9]
port 126 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 sram_web0
port 127 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 sram_wmask0[0]
port 128 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 sram_wmask0[1]
port 129 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 sram_wmask0[2]
port 130 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 sram_wmask0[3]
port 131 nsew signal output
rlabel metal4 s 4208 2128 4528 39760 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 39760 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 39760 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 39760 6 vssd1
port 133 nsew ground bidirectional
rlabel metal3 s 0 688 800 808 6 wb_ack_o
port 134 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 wb_adr_i[0]
port 135 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 wb_adr_i[10]
port 136 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[11]
port 137 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[12]
port 138 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[13]
port 139 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[14]
port 140 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 wb_adr_i[15]
port 141 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wb_adr_i[16]
port 142 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 wb_adr_i[17]
port 143 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 wb_adr_i[18]
port 144 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 wb_adr_i[19]
port 145 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wb_adr_i[1]
port 146 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 wb_adr_i[20]
port 147 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wb_adr_i[21]
port 148 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 wb_adr_i[22]
port 149 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 wb_adr_i[23]
port 150 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wb_adr_i[2]
port 151 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wb_adr_i[3]
port 152 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 wb_adr_i[4]
port 153 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 wb_adr_i[5]
port 154 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wb_adr_i[6]
port 155 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wb_adr_i[7]
port 156 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wb_adr_i[8]
port 157 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 wb_adr_i[9]
port 158 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 wb_clk_i
port 159 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 wb_cyc_i
port 160 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wb_data_i[0]
port 161 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 wb_data_i[10]
port 162 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[11]
port 163 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[12]
port 164 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[13]
port 165 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[14]
port 166 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wb_data_i[15]
port 167 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 wb_data_i[16]
port 168 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wb_data_i[17]
port 169 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 wb_data_i[18]
port 170 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wb_data_i[19]
port 171 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 wb_data_i[1]
port 172 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 wb_data_i[20]
port 173 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 wb_data_i[21]
port 174 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_data_i[22]
port 175 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_data_i[23]
port 176 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 wb_data_i[24]
port 177 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 wb_data_i[25]
port 178 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 wb_data_i[26]
port 179 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 wb_data_i[27]
port 180 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 wb_data_i[28]
port 181 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 wb_data_i[29]
port 182 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wb_data_i[2]
port 183 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 wb_data_i[30]
port 184 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 wb_data_i[31]
port 185 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 wb_data_i[3]
port 186 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wb_data_i[4]
port 187 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 wb_data_i[5]
port 188 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 wb_data_i[6]
port 189 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wb_data_i[7]
port 190 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wb_data_i[8]
port 191 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wb_data_i[9]
port 192 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wb_data_o[0]
port 193 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 wb_data_o[10]
port 194 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[11]
port 195 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[12]
port 196 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[13]
port 197 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 wb_data_o[14]
port 198 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 wb_data_o[15]
port 199 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 wb_data_o[16]
port 200 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 wb_data_o[17]
port 201 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 wb_data_o[18]
port 202 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 wb_data_o[19]
port 203 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 wb_data_o[1]
port 204 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 wb_data_o[20]
port 205 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 wb_data_o[21]
port 206 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 wb_data_o[22]
port 207 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 wb_data_o[23]
port 208 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 wb_data_o[24]
port 209 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 wb_data_o[25]
port 210 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 wb_data_o[26]
port 211 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 wb_data_o[27]
port 212 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 wb_data_o[28]
port 213 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 wb_data_o[29]
port 214 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 wb_data_o[2]
port 215 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 wb_data_o[30]
port 216 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 wb_data_o[31]
port 217 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 wb_data_o[3]
port 218 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 wb_data_o[4]
port 219 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 wb_data_o[5]
port 220 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 wb_data_o[6]
port 221 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 wb_data_o[7]
port 222 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 wb_data_o[8]
port 223 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 wb_data_o[9]
port 224 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 wb_error_o
port 225 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 wb_rst_i
port 226 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wb_sel_i[0]
port 227 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_sel_i[1]
port 228 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_sel_i[2]
port 229 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 wb_sel_i[3]
port 230 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wb_stall_o
port 231 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 wb_stb_i
port 232 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 wb_we_i
port 233 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3234766
string GDS_FILE /mnt/f/WSL/ASIC/ExperiarSoC/openlane/Flash/runs/23_05_12_10_06/results/signoff/Flash.magic.gds
string GDS_START 537644
<< end >>

