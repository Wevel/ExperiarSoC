magic
tech sky130A
magscale 1 2
timestamp 1654264013
<< obsli1 >>
rect 1104 2159 88872 177361
<< obsm1 >>
rect 14 688 89962 177880
<< metal2 >>
rect 1030 179200 1086 180000
rect 3146 179200 3202 180000
rect 5262 179200 5318 180000
rect 7378 179200 7434 180000
rect 9586 179200 9642 180000
rect 11702 179200 11758 180000
rect 13818 179200 13874 180000
rect 16026 179200 16082 180000
rect 18142 179200 18198 180000
rect 20258 179200 20314 180000
rect 22374 179200 22430 180000
rect 24582 179200 24638 180000
rect 26698 179200 26754 180000
rect 28814 179200 28870 180000
rect 31022 179200 31078 180000
rect 33138 179200 33194 180000
rect 35254 179200 35310 180000
rect 37370 179200 37426 180000
rect 39578 179200 39634 180000
rect 41694 179200 41750 180000
rect 43810 179200 43866 180000
rect 46018 179200 46074 180000
rect 48134 179200 48190 180000
rect 50250 179200 50306 180000
rect 52366 179200 52422 180000
rect 54574 179200 54630 180000
rect 56690 179200 56746 180000
rect 58806 179200 58862 180000
rect 61014 179200 61070 180000
rect 63130 179200 63186 180000
rect 65246 179200 65302 180000
rect 67362 179200 67418 180000
rect 69570 179200 69626 180000
rect 71686 179200 71742 180000
rect 73802 179200 73858 180000
rect 76010 179200 76066 180000
rect 78126 179200 78182 180000
rect 80242 179200 80298 180000
rect 82358 179200 82414 180000
rect 84566 179200 84622 180000
rect 86682 179200 86738 180000
rect 88798 179200 88854 180000
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11242 0 11298 800
rect 12714 0 12770 800
rect 14186 0 14242 800
rect 15750 0 15806 800
rect 17222 0 17278 800
rect 18694 0 18750 800
rect 20166 0 20222 800
rect 21730 0 21786 800
rect 23202 0 23258 800
rect 24674 0 24730 800
rect 26238 0 26294 800
rect 27710 0 27766 800
rect 29182 0 29238 800
rect 30746 0 30802 800
rect 32218 0 32274 800
rect 33690 0 33746 800
rect 35162 0 35218 800
rect 36726 0 36782 800
rect 38198 0 38254 800
rect 39670 0 39726 800
rect 41234 0 41290 800
rect 42706 0 42762 800
rect 44178 0 44234 800
rect 45742 0 45798 800
rect 47214 0 47270 800
rect 48686 0 48742 800
rect 50158 0 50214 800
rect 51722 0 51778 800
rect 53194 0 53250 800
rect 54666 0 54722 800
rect 56230 0 56286 800
rect 57702 0 57758 800
rect 59174 0 59230 800
rect 60738 0 60794 800
rect 62210 0 62266 800
rect 63682 0 63738 800
rect 65154 0 65210 800
rect 66718 0 66774 800
rect 68190 0 68246 800
rect 69662 0 69718 800
rect 71226 0 71282 800
rect 72698 0 72754 800
rect 74170 0 74226 800
rect 75734 0 75790 800
rect 77206 0 77262 800
rect 78678 0 78734 800
rect 80150 0 80206 800
rect 81714 0 81770 800
rect 83186 0 83242 800
rect 84658 0 84714 800
rect 86222 0 86278 800
rect 87694 0 87750 800
rect 89166 0 89222 800
<< obsm2 >>
rect 18 179144 974 179625
rect 1142 179144 3090 179625
rect 3258 179144 5206 179625
rect 5374 179144 7322 179625
rect 7490 179144 9530 179625
rect 9698 179144 11646 179625
rect 11814 179144 13762 179625
rect 13930 179144 15970 179625
rect 16138 179144 18086 179625
rect 18254 179144 20202 179625
rect 20370 179144 22318 179625
rect 22486 179144 24526 179625
rect 24694 179144 26642 179625
rect 26810 179144 28758 179625
rect 28926 179144 30966 179625
rect 31134 179144 33082 179625
rect 33250 179144 35198 179625
rect 35366 179144 37314 179625
rect 37482 179144 39522 179625
rect 39690 179144 41638 179625
rect 41806 179144 43754 179625
rect 43922 179144 45962 179625
rect 46130 179144 48078 179625
rect 48246 179144 50194 179625
rect 50362 179144 52310 179625
rect 52478 179144 54518 179625
rect 54686 179144 56634 179625
rect 56802 179144 58750 179625
rect 58918 179144 60958 179625
rect 61126 179144 63074 179625
rect 63242 179144 65190 179625
rect 65358 179144 67306 179625
rect 67474 179144 69514 179625
rect 69682 179144 71630 179625
rect 71798 179144 73746 179625
rect 73914 179144 75954 179625
rect 76122 179144 78070 179625
rect 78238 179144 80186 179625
rect 80354 179144 82302 179625
rect 82470 179144 84510 179625
rect 84678 179144 86626 179625
rect 86794 179144 88742 179625
rect 88910 179144 89958 179625
rect 18 856 89958 179144
rect 18 439 698 856
rect 866 439 2170 856
rect 2338 439 3642 856
rect 3810 439 5114 856
rect 5282 439 6678 856
rect 6846 439 8150 856
rect 8318 439 9622 856
rect 9790 439 11186 856
rect 11354 439 12658 856
rect 12826 439 14130 856
rect 14298 439 15694 856
rect 15862 439 17166 856
rect 17334 439 18638 856
rect 18806 439 20110 856
rect 20278 439 21674 856
rect 21842 439 23146 856
rect 23314 439 24618 856
rect 24786 439 26182 856
rect 26350 439 27654 856
rect 27822 439 29126 856
rect 29294 439 30690 856
rect 30858 439 32162 856
rect 32330 439 33634 856
rect 33802 439 35106 856
rect 35274 439 36670 856
rect 36838 439 38142 856
rect 38310 439 39614 856
rect 39782 439 41178 856
rect 41346 439 42650 856
rect 42818 439 44122 856
rect 44290 439 45686 856
rect 45854 439 47158 856
rect 47326 439 48630 856
rect 48798 439 50102 856
rect 50270 439 51666 856
rect 51834 439 53138 856
rect 53306 439 54610 856
rect 54778 439 56174 856
rect 56342 439 57646 856
rect 57814 439 59118 856
rect 59286 439 60682 856
rect 60850 439 62154 856
rect 62322 439 63626 856
rect 63794 439 65098 856
rect 65266 439 66662 856
rect 66830 439 68134 856
rect 68302 439 69606 856
rect 69774 439 71170 856
rect 71338 439 72642 856
rect 72810 439 74114 856
rect 74282 439 75678 856
rect 75846 439 77150 856
rect 77318 439 78622 856
rect 78790 439 80094 856
rect 80262 439 81658 856
rect 81826 439 83130 856
rect 83298 439 84602 856
rect 84770 439 86166 856
rect 86334 439 87638 856
rect 87806 439 89110 856
rect 89278 439 89958 856
<< metal3 >>
rect 0 179528 800 179648
rect 89200 179528 90000 179648
rect 0 178576 800 178696
rect 89200 178712 90000 178832
rect 0 177624 800 177744
rect 89200 177760 90000 177880
rect 0 176808 800 176928
rect 89200 176944 90000 177064
rect 0 175856 800 175976
rect 89200 175992 90000 176112
rect 89200 175176 90000 175296
rect 0 174904 800 175024
rect 89200 174360 90000 174480
rect 0 173952 800 174072
rect 89200 173408 90000 173528
rect 0 173136 800 173256
rect 89200 172592 90000 172712
rect 0 172184 800 172304
rect 89200 171640 90000 171760
rect 0 171232 800 171352
rect 89200 170824 90000 170944
rect 0 170416 800 170536
rect 89200 169872 90000 169992
rect 0 169464 800 169584
rect 89200 169056 90000 169176
rect 0 168512 800 168632
rect 89200 168240 90000 168360
rect 0 167560 800 167680
rect 89200 167288 90000 167408
rect 0 166744 800 166864
rect 89200 166472 90000 166592
rect 0 165792 800 165912
rect 89200 165520 90000 165640
rect 0 164840 800 164960
rect 89200 164704 90000 164824
rect 0 164024 800 164144
rect 89200 163752 90000 163872
rect 0 163072 800 163192
rect 89200 162936 90000 163056
rect 0 162120 800 162240
rect 89200 162120 90000 162240
rect 0 161168 800 161288
rect 89200 161168 90000 161288
rect 0 160352 800 160472
rect 89200 160352 90000 160472
rect 0 159400 800 159520
rect 89200 159400 90000 159520
rect 0 158448 800 158568
rect 89200 158584 90000 158704
rect 0 157496 800 157616
rect 89200 157632 90000 157752
rect 0 156680 800 156800
rect 89200 156816 90000 156936
rect 89200 156000 90000 156120
rect 0 155728 800 155848
rect 89200 155048 90000 155168
rect 0 154776 800 154896
rect 89200 154232 90000 154352
rect 0 153960 800 154080
rect 89200 153280 90000 153400
rect 0 153008 800 153128
rect 89200 152464 90000 152584
rect 0 152056 800 152176
rect 89200 151512 90000 151632
rect 0 151104 800 151224
rect 89200 150696 90000 150816
rect 0 150288 800 150408
rect 89200 149880 90000 150000
rect 0 149336 800 149456
rect 89200 148928 90000 149048
rect 0 148384 800 148504
rect 89200 148112 90000 148232
rect 0 147568 800 147688
rect 89200 147160 90000 147280
rect 0 146616 800 146736
rect 89200 146344 90000 146464
rect 0 145664 800 145784
rect 89200 145392 90000 145512
rect 0 144712 800 144832
rect 89200 144576 90000 144696
rect 0 143896 800 144016
rect 89200 143760 90000 143880
rect 0 142944 800 143064
rect 89200 142808 90000 142928
rect 0 141992 800 142112
rect 89200 141992 90000 142112
rect 0 141176 800 141296
rect 89200 141040 90000 141160
rect 0 140224 800 140344
rect 89200 140224 90000 140344
rect 0 139272 800 139392
rect 89200 139272 90000 139392
rect 0 138320 800 138440
rect 89200 138456 90000 138576
rect 0 137504 800 137624
rect 89200 137640 90000 137760
rect 0 136552 800 136672
rect 89200 136688 90000 136808
rect 89200 135872 90000 135992
rect 0 135600 800 135720
rect 89200 134920 90000 135040
rect 0 134648 800 134768
rect 89200 134104 90000 134224
rect 0 133832 800 133952
rect 89200 133152 90000 133272
rect 0 132880 800 133000
rect 89200 132336 90000 132456
rect 0 131928 800 132048
rect 89200 131520 90000 131640
rect 0 131112 800 131232
rect 89200 130568 90000 130688
rect 0 130160 800 130280
rect 89200 129752 90000 129872
rect 0 129208 800 129328
rect 89200 128800 90000 128920
rect 0 128256 800 128376
rect 89200 127984 90000 128104
rect 0 127440 800 127560
rect 89200 127032 90000 127152
rect 0 126488 800 126608
rect 89200 126216 90000 126336
rect 0 125536 800 125656
rect 89200 125400 90000 125520
rect 0 124720 800 124840
rect 89200 124448 90000 124568
rect 0 123768 800 123888
rect 89200 123632 90000 123752
rect 0 122816 800 122936
rect 89200 122680 90000 122800
rect 0 121864 800 121984
rect 89200 121864 90000 121984
rect 0 121048 800 121168
rect 89200 120912 90000 121032
rect 0 120096 800 120216
rect 89200 120096 90000 120216
rect 0 119144 800 119264
rect 89200 119280 90000 119400
rect 0 118192 800 118312
rect 89200 118328 90000 118448
rect 0 117376 800 117496
rect 89200 117512 90000 117632
rect 0 116424 800 116544
rect 89200 116560 90000 116680
rect 89200 115744 90000 115864
rect 0 115472 800 115592
rect 0 114656 800 114776
rect 89200 114792 90000 114912
rect 89200 113976 90000 114096
rect 0 113704 800 113824
rect 89200 113160 90000 113280
rect 0 112752 800 112872
rect 89200 112208 90000 112328
rect 0 111800 800 111920
rect 89200 111392 90000 111512
rect 0 110984 800 111104
rect 89200 110440 90000 110560
rect 0 110032 800 110152
rect 89200 109624 90000 109744
rect 0 109080 800 109200
rect 89200 108672 90000 108792
rect 0 108264 800 108384
rect 89200 107856 90000 107976
rect 0 107312 800 107432
rect 89200 107040 90000 107160
rect 0 106360 800 106480
rect 89200 106088 90000 106208
rect 0 105408 800 105528
rect 89200 105272 90000 105392
rect 0 104592 800 104712
rect 89200 104320 90000 104440
rect 0 103640 800 103760
rect 89200 103504 90000 103624
rect 0 102688 800 102808
rect 89200 102552 90000 102672
rect 0 101872 800 101992
rect 89200 101736 90000 101856
rect 0 100920 800 101040
rect 89200 100920 90000 101040
rect 0 99968 800 100088
rect 89200 99968 90000 100088
rect 0 99016 800 99136
rect 89200 99152 90000 99272
rect 0 98200 800 98320
rect 89200 98200 90000 98320
rect 0 97248 800 97368
rect 89200 97384 90000 97504
rect 0 96296 800 96416
rect 89200 96432 90000 96552
rect 89200 95616 90000 95736
rect 0 95344 800 95464
rect 89200 94800 90000 94920
rect 0 94528 800 94648
rect 89200 93848 90000 93968
rect 0 93576 800 93696
rect 89200 93032 90000 93152
rect 0 92624 800 92744
rect 89200 92080 90000 92200
rect 0 91808 800 91928
rect 89200 91264 90000 91384
rect 0 90856 800 90976
rect 89200 90448 90000 90568
rect 0 89904 800 90024
rect 89200 89496 90000 89616
rect 0 88952 800 89072
rect 89200 88680 90000 88800
rect 0 88136 800 88256
rect 89200 87728 90000 87848
rect 0 87184 800 87304
rect 89200 86912 90000 87032
rect 0 86232 800 86352
rect 89200 85960 90000 86080
rect 0 85416 800 85536
rect 89200 85144 90000 85264
rect 0 84464 800 84584
rect 89200 84328 90000 84448
rect 0 83512 800 83632
rect 89200 83376 90000 83496
rect 0 82560 800 82680
rect 89200 82560 90000 82680
rect 0 81744 800 81864
rect 89200 81608 90000 81728
rect 0 80792 800 80912
rect 89200 80792 90000 80912
rect 0 79840 800 79960
rect 89200 79840 90000 79960
rect 0 78888 800 79008
rect 89200 79024 90000 79144
rect 0 78072 800 78192
rect 89200 78208 90000 78328
rect 0 77120 800 77240
rect 89200 77256 90000 77376
rect 89200 76440 90000 76560
rect 0 76168 800 76288
rect 0 75352 800 75472
rect 89200 75488 90000 75608
rect 89200 74672 90000 74792
rect 0 74400 800 74520
rect 89200 73720 90000 73840
rect 0 73448 800 73568
rect 89200 72904 90000 73024
rect 0 72496 800 72616
rect 89200 72088 90000 72208
rect 0 71680 800 71800
rect 89200 71136 90000 71256
rect 0 70728 800 70848
rect 89200 70320 90000 70440
rect 0 69776 800 69896
rect 89200 69368 90000 69488
rect 0 68960 800 69080
rect 89200 68552 90000 68672
rect 0 68008 800 68128
rect 89200 67600 90000 67720
rect 0 67056 800 67176
rect 89200 66784 90000 66904
rect 0 66104 800 66224
rect 89200 65968 90000 66088
rect 0 65288 800 65408
rect 89200 65016 90000 65136
rect 0 64336 800 64456
rect 89200 64200 90000 64320
rect 0 63384 800 63504
rect 89200 63248 90000 63368
rect 0 62568 800 62688
rect 89200 62432 90000 62552
rect 0 61616 800 61736
rect 89200 61480 90000 61600
rect 0 60664 800 60784
rect 89200 60664 90000 60784
rect 0 59712 800 59832
rect 89200 59848 90000 59968
rect 0 58896 800 59016
rect 89200 58896 90000 59016
rect 0 57944 800 58064
rect 89200 58080 90000 58200
rect 0 56992 800 57112
rect 89200 57128 90000 57248
rect 89200 56312 90000 56432
rect 0 56040 800 56160
rect 0 55224 800 55344
rect 89200 55360 90000 55480
rect 89200 54544 90000 54664
rect 0 54272 800 54392
rect 89200 53728 90000 53848
rect 0 53320 800 53440
rect 89200 52776 90000 52896
rect 0 52504 800 52624
rect 89200 51960 90000 52080
rect 0 51552 800 51672
rect 89200 51008 90000 51128
rect 0 50600 800 50720
rect 89200 50192 90000 50312
rect 0 49648 800 49768
rect 89200 49240 90000 49360
rect 0 48832 800 48952
rect 89200 48424 90000 48544
rect 0 47880 800 48000
rect 89200 47608 90000 47728
rect 0 46928 800 47048
rect 89200 46656 90000 46776
rect 0 46112 800 46232
rect 89200 45840 90000 45960
rect 0 45160 800 45280
rect 89200 44888 90000 45008
rect 0 44208 800 44328
rect 89200 44072 90000 44192
rect 0 43256 800 43376
rect 89200 43120 90000 43240
rect 0 42440 800 42560
rect 89200 42304 90000 42424
rect 0 41488 800 41608
rect 89200 41488 90000 41608
rect 0 40536 800 40656
rect 89200 40536 90000 40656
rect 0 39584 800 39704
rect 89200 39720 90000 39840
rect 0 38768 800 38888
rect 89200 38768 90000 38888
rect 0 37816 800 37936
rect 89200 37952 90000 38072
rect 0 36864 800 36984
rect 89200 37000 90000 37120
rect 0 36048 800 36168
rect 89200 36184 90000 36304
rect 89200 35368 90000 35488
rect 0 35096 800 35216
rect 89200 34416 90000 34536
rect 0 34144 800 34264
rect 89200 33600 90000 33720
rect 0 33192 800 33312
rect 89200 32648 90000 32768
rect 0 32376 800 32496
rect 89200 31832 90000 31952
rect 0 31424 800 31544
rect 89200 30880 90000 31000
rect 0 30472 800 30592
rect 89200 30064 90000 30184
rect 0 29656 800 29776
rect 89200 29248 90000 29368
rect 0 28704 800 28824
rect 89200 28296 90000 28416
rect 0 27752 800 27872
rect 89200 27480 90000 27600
rect 0 26800 800 26920
rect 89200 26528 90000 26648
rect 0 25984 800 26104
rect 89200 25712 90000 25832
rect 0 25032 800 25152
rect 89200 24760 90000 24880
rect 0 24080 800 24200
rect 89200 23944 90000 24064
rect 0 23264 800 23384
rect 89200 23128 90000 23248
rect 0 22312 800 22432
rect 89200 22176 90000 22296
rect 0 21360 800 21480
rect 89200 21360 90000 21480
rect 0 20408 800 20528
rect 89200 20408 90000 20528
rect 0 19592 800 19712
rect 89200 19592 90000 19712
rect 0 18640 800 18760
rect 89200 18640 90000 18760
rect 0 17688 800 17808
rect 89200 17824 90000 17944
rect 89200 17008 90000 17128
rect 0 16736 800 16856
rect 0 15920 800 16040
rect 89200 16056 90000 16176
rect 89200 15240 90000 15360
rect 0 14968 800 15088
rect 89200 14288 90000 14408
rect 0 14016 800 14136
rect 89200 13472 90000 13592
rect 0 13200 800 13320
rect 89200 12520 90000 12640
rect 0 12248 800 12368
rect 89200 11704 90000 11824
rect 0 11296 800 11416
rect 89200 10888 90000 11008
rect 0 10344 800 10464
rect 89200 9936 90000 10056
rect 0 9528 800 9648
rect 89200 9120 90000 9240
rect 0 8576 800 8696
rect 89200 8168 90000 8288
rect 0 7624 800 7744
rect 89200 7352 90000 7472
rect 0 6808 800 6928
rect 89200 6400 90000 6520
rect 0 5856 800 5976
rect 89200 5584 90000 5704
rect 0 4904 800 5024
rect 89200 4768 90000 4888
rect 0 3952 800 4072
rect 89200 3816 90000 3936
rect 0 3136 800 3256
rect 89200 3000 90000 3120
rect 0 2184 800 2304
rect 89200 2048 90000 2168
rect 0 1232 800 1352
rect 89200 1232 90000 1352
rect 0 416 800 536
rect 89200 416 90000 536
<< obsm3 >>
rect 880 179448 89120 179621
rect 13 178912 89963 179448
rect 13 178776 89120 178912
rect 880 178632 89120 178776
rect 880 178496 89963 178632
rect 13 177960 89963 178496
rect 13 177824 89120 177960
rect 880 177680 89120 177824
rect 880 177544 89963 177680
rect 13 177144 89963 177544
rect 13 177008 89120 177144
rect 880 176864 89120 177008
rect 880 176728 89963 176864
rect 13 176192 89963 176728
rect 13 176056 89120 176192
rect 880 175912 89120 176056
rect 880 175776 89963 175912
rect 13 175376 89963 175776
rect 13 175104 89120 175376
rect 880 175096 89120 175104
rect 880 174824 89963 175096
rect 13 174560 89963 174824
rect 13 174280 89120 174560
rect 13 174152 89963 174280
rect 880 173872 89963 174152
rect 13 173608 89963 173872
rect 13 173336 89120 173608
rect 880 173328 89120 173336
rect 880 173056 89963 173328
rect 13 172792 89963 173056
rect 13 172512 89120 172792
rect 13 172384 89963 172512
rect 880 172104 89963 172384
rect 13 171840 89963 172104
rect 13 171560 89120 171840
rect 13 171432 89963 171560
rect 880 171152 89963 171432
rect 13 171024 89963 171152
rect 13 170744 89120 171024
rect 13 170616 89963 170744
rect 880 170336 89963 170616
rect 13 170072 89963 170336
rect 13 169792 89120 170072
rect 13 169664 89963 169792
rect 880 169384 89963 169664
rect 13 169256 89963 169384
rect 13 168976 89120 169256
rect 13 168712 89963 168976
rect 880 168440 89963 168712
rect 880 168432 89120 168440
rect 13 168160 89120 168432
rect 13 167760 89963 168160
rect 880 167488 89963 167760
rect 880 167480 89120 167488
rect 13 167208 89120 167480
rect 13 166944 89963 167208
rect 880 166672 89963 166944
rect 880 166664 89120 166672
rect 13 166392 89120 166664
rect 13 165992 89963 166392
rect 880 165720 89963 165992
rect 880 165712 89120 165720
rect 13 165440 89120 165712
rect 13 165040 89963 165440
rect 880 164904 89963 165040
rect 880 164760 89120 164904
rect 13 164624 89120 164760
rect 13 164224 89963 164624
rect 880 163952 89963 164224
rect 880 163944 89120 163952
rect 13 163672 89120 163944
rect 13 163272 89963 163672
rect 880 163136 89963 163272
rect 880 162992 89120 163136
rect 13 162856 89120 162992
rect 13 162320 89963 162856
rect 880 162040 89120 162320
rect 13 161368 89963 162040
rect 880 161088 89120 161368
rect 13 160552 89963 161088
rect 880 160272 89120 160552
rect 13 159600 89963 160272
rect 880 159320 89120 159600
rect 13 158784 89963 159320
rect 13 158648 89120 158784
rect 880 158504 89120 158648
rect 880 158368 89963 158504
rect 13 157832 89963 158368
rect 13 157696 89120 157832
rect 880 157552 89120 157696
rect 880 157416 89963 157552
rect 13 157016 89963 157416
rect 13 156880 89120 157016
rect 880 156736 89120 156880
rect 880 156600 89963 156736
rect 13 156200 89963 156600
rect 13 155928 89120 156200
rect 880 155920 89120 155928
rect 880 155648 89963 155920
rect 13 155248 89963 155648
rect 13 154976 89120 155248
rect 880 154968 89120 154976
rect 880 154696 89963 154968
rect 13 154432 89963 154696
rect 13 154160 89120 154432
rect 880 154152 89120 154160
rect 880 153880 89963 154152
rect 13 153480 89963 153880
rect 13 153208 89120 153480
rect 880 153200 89120 153208
rect 880 152928 89963 153200
rect 13 152664 89963 152928
rect 13 152384 89120 152664
rect 13 152256 89963 152384
rect 880 151976 89963 152256
rect 13 151712 89963 151976
rect 13 151432 89120 151712
rect 13 151304 89963 151432
rect 880 151024 89963 151304
rect 13 150896 89963 151024
rect 13 150616 89120 150896
rect 13 150488 89963 150616
rect 880 150208 89963 150488
rect 13 150080 89963 150208
rect 13 149800 89120 150080
rect 13 149536 89963 149800
rect 880 149256 89963 149536
rect 13 149128 89963 149256
rect 13 148848 89120 149128
rect 13 148584 89963 148848
rect 880 148312 89963 148584
rect 880 148304 89120 148312
rect 13 148032 89120 148304
rect 13 147768 89963 148032
rect 880 147488 89963 147768
rect 13 147360 89963 147488
rect 13 147080 89120 147360
rect 13 146816 89963 147080
rect 880 146544 89963 146816
rect 880 146536 89120 146544
rect 13 146264 89120 146536
rect 13 145864 89963 146264
rect 880 145592 89963 145864
rect 880 145584 89120 145592
rect 13 145312 89120 145584
rect 13 144912 89963 145312
rect 880 144776 89963 144912
rect 880 144632 89120 144776
rect 13 144496 89120 144632
rect 13 144096 89963 144496
rect 880 143960 89963 144096
rect 880 143816 89120 143960
rect 13 143680 89120 143816
rect 13 143144 89963 143680
rect 880 143008 89963 143144
rect 880 142864 89120 143008
rect 13 142728 89120 142864
rect 13 142192 89963 142728
rect 880 141912 89120 142192
rect 13 141376 89963 141912
rect 880 141240 89963 141376
rect 880 141096 89120 141240
rect 13 140960 89120 141096
rect 13 140424 89963 140960
rect 880 140144 89120 140424
rect 13 139472 89963 140144
rect 880 139192 89120 139472
rect 13 138656 89963 139192
rect 13 138520 89120 138656
rect 880 138376 89120 138520
rect 880 138240 89963 138376
rect 13 137840 89963 138240
rect 13 137704 89120 137840
rect 880 137560 89120 137704
rect 880 137424 89963 137560
rect 13 136888 89963 137424
rect 13 136752 89120 136888
rect 880 136608 89120 136752
rect 880 136472 89963 136608
rect 13 136072 89963 136472
rect 13 135800 89120 136072
rect 880 135792 89120 135800
rect 880 135520 89963 135792
rect 13 135120 89963 135520
rect 13 134848 89120 135120
rect 880 134840 89120 134848
rect 880 134568 89963 134840
rect 13 134304 89963 134568
rect 13 134032 89120 134304
rect 880 134024 89120 134032
rect 880 133752 89963 134024
rect 13 133352 89963 133752
rect 13 133080 89120 133352
rect 880 133072 89120 133080
rect 880 132800 89963 133072
rect 13 132536 89963 132800
rect 13 132256 89120 132536
rect 13 132128 89963 132256
rect 880 131848 89963 132128
rect 13 131720 89963 131848
rect 13 131440 89120 131720
rect 13 131312 89963 131440
rect 880 131032 89963 131312
rect 13 130768 89963 131032
rect 13 130488 89120 130768
rect 13 130360 89963 130488
rect 880 130080 89963 130360
rect 13 129952 89963 130080
rect 13 129672 89120 129952
rect 13 129408 89963 129672
rect 880 129128 89963 129408
rect 13 129000 89963 129128
rect 13 128720 89120 129000
rect 13 128456 89963 128720
rect 880 128184 89963 128456
rect 880 128176 89120 128184
rect 13 127904 89120 128176
rect 13 127640 89963 127904
rect 880 127360 89963 127640
rect 13 127232 89963 127360
rect 13 126952 89120 127232
rect 13 126688 89963 126952
rect 880 126416 89963 126688
rect 880 126408 89120 126416
rect 13 126136 89120 126408
rect 13 125736 89963 126136
rect 880 125600 89963 125736
rect 880 125456 89120 125600
rect 13 125320 89120 125456
rect 13 124920 89963 125320
rect 880 124648 89963 124920
rect 880 124640 89120 124648
rect 13 124368 89120 124640
rect 13 123968 89963 124368
rect 880 123832 89963 123968
rect 880 123688 89120 123832
rect 13 123552 89120 123688
rect 13 123016 89963 123552
rect 880 122880 89963 123016
rect 880 122736 89120 122880
rect 13 122600 89120 122736
rect 13 122064 89963 122600
rect 880 121784 89120 122064
rect 13 121248 89963 121784
rect 880 121112 89963 121248
rect 880 120968 89120 121112
rect 13 120832 89120 120968
rect 13 120296 89963 120832
rect 880 120016 89120 120296
rect 13 119480 89963 120016
rect 13 119344 89120 119480
rect 880 119200 89120 119344
rect 880 119064 89963 119200
rect 13 118528 89963 119064
rect 13 118392 89120 118528
rect 880 118248 89120 118392
rect 880 118112 89963 118248
rect 13 117712 89963 118112
rect 13 117576 89120 117712
rect 880 117432 89120 117576
rect 880 117296 89963 117432
rect 13 116760 89963 117296
rect 13 116624 89120 116760
rect 880 116480 89120 116624
rect 880 116344 89963 116480
rect 13 115944 89963 116344
rect 13 115672 89120 115944
rect 880 115664 89120 115672
rect 880 115392 89963 115664
rect 13 114992 89963 115392
rect 13 114856 89120 114992
rect 880 114712 89120 114856
rect 880 114576 89963 114712
rect 13 114176 89963 114576
rect 13 113904 89120 114176
rect 880 113896 89120 113904
rect 880 113624 89963 113896
rect 13 113360 89963 113624
rect 13 113080 89120 113360
rect 13 112952 89963 113080
rect 880 112672 89963 112952
rect 13 112408 89963 112672
rect 13 112128 89120 112408
rect 13 112000 89963 112128
rect 880 111720 89963 112000
rect 13 111592 89963 111720
rect 13 111312 89120 111592
rect 13 111184 89963 111312
rect 880 110904 89963 111184
rect 13 110640 89963 110904
rect 13 110360 89120 110640
rect 13 110232 89963 110360
rect 880 109952 89963 110232
rect 13 109824 89963 109952
rect 13 109544 89120 109824
rect 13 109280 89963 109544
rect 880 109000 89963 109280
rect 13 108872 89963 109000
rect 13 108592 89120 108872
rect 13 108464 89963 108592
rect 880 108184 89963 108464
rect 13 108056 89963 108184
rect 13 107776 89120 108056
rect 13 107512 89963 107776
rect 880 107240 89963 107512
rect 880 107232 89120 107240
rect 13 106960 89120 107232
rect 13 106560 89963 106960
rect 880 106288 89963 106560
rect 880 106280 89120 106288
rect 13 106008 89120 106280
rect 13 105608 89963 106008
rect 880 105472 89963 105608
rect 880 105328 89120 105472
rect 13 105192 89120 105328
rect 13 104792 89963 105192
rect 880 104520 89963 104792
rect 880 104512 89120 104520
rect 13 104240 89120 104512
rect 13 103840 89963 104240
rect 880 103704 89963 103840
rect 880 103560 89120 103704
rect 13 103424 89120 103560
rect 13 102888 89963 103424
rect 880 102752 89963 102888
rect 880 102608 89120 102752
rect 13 102472 89120 102608
rect 13 102072 89963 102472
rect 880 101936 89963 102072
rect 880 101792 89120 101936
rect 13 101656 89120 101792
rect 13 101120 89963 101656
rect 880 100840 89120 101120
rect 13 100168 89963 100840
rect 880 99888 89120 100168
rect 13 99352 89963 99888
rect 13 99216 89120 99352
rect 880 99072 89120 99216
rect 880 98936 89963 99072
rect 13 98400 89963 98936
rect 880 98120 89120 98400
rect 13 97584 89963 98120
rect 13 97448 89120 97584
rect 880 97304 89120 97448
rect 880 97168 89963 97304
rect 13 96632 89963 97168
rect 13 96496 89120 96632
rect 880 96352 89120 96496
rect 880 96216 89963 96352
rect 13 95816 89963 96216
rect 13 95544 89120 95816
rect 880 95536 89120 95544
rect 880 95264 89963 95536
rect 13 95000 89963 95264
rect 13 94728 89120 95000
rect 880 94720 89120 94728
rect 880 94448 89963 94720
rect 13 94048 89963 94448
rect 13 93776 89120 94048
rect 880 93768 89120 93776
rect 880 93496 89963 93768
rect 13 93232 89963 93496
rect 13 92952 89120 93232
rect 13 92824 89963 92952
rect 880 92544 89963 92824
rect 13 92280 89963 92544
rect 13 92008 89120 92280
rect 880 92000 89120 92008
rect 880 91728 89963 92000
rect 13 91464 89963 91728
rect 13 91184 89120 91464
rect 13 91056 89963 91184
rect 880 90776 89963 91056
rect 13 90648 89963 90776
rect 13 90368 89120 90648
rect 13 90104 89963 90368
rect 880 89824 89963 90104
rect 13 89696 89963 89824
rect 13 89416 89120 89696
rect 13 89152 89963 89416
rect 880 88880 89963 89152
rect 880 88872 89120 88880
rect 13 88600 89120 88872
rect 13 88336 89963 88600
rect 880 88056 89963 88336
rect 13 87928 89963 88056
rect 13 87648 89120 87928
rect 13 87384 89963 87648
rect 880 87112 89963 87384
rect 880 87104 89120 87112
rect 13 86832 89120 87104
rect 13 86432 89963 86832
rect 880 86160 89963 86432
rect 880 86152 89120 86160
rect 13 85880 89120 86152
rect 13 85616 89963 85880
rect 880 85344 89963 85616
rect 880 85336 89120 85344
rect 13 85064 89120 85336
rect 13 84664 89963 85064
rect 880 84528 89963 84664
rect 880 84384 89120 84528
rect 13 84248 89120 84384
rect 13 83712 89963 84248
rect 880 83576 89963 83712
rect 880 83432 89120 83576
rect 13 83296 89120 83432
rect 13 82760 89963 83296
rect 880 82480 89120 82760
rect 13 81944 89963 82480
rect 880 81808 89963 81944
rect 880 81664 89120 81808
rect 13 81528 89120 81664
rect 13 80992 89963 81528
rect 880 80712 89120 80992
rect 13 80040 89963 80712
rect 880 79760 89120 80040
rect 13 79224 89963 79760
rect 13 79088 89120 79224
rect 880 78944 89120 79088
rect 880 78808 89963 78944
rect 13 78408 89963 78808
rect 13 78272 89120 78408
rect 880 78128 89120 78272
rect 880 77992 89963 78128
rect 13 77456 89963 77992
rect 13 77320 89120 77456
rect 880 77176 89120 77320
rect 880 77040 89963 77176
rect 13 76640 89963 77040
rect 13 76368 89120 76640
rect 880 76360 89120 76368
rect 880 76088 89963 76360
rect 13 75688 89963 76088
rect 13 75552 89120 75688
rect 880 75408 89120 75552
rect 880 75272 89963 75408
rect 13 74872 89963 75272
rect 13 74600 89120 74872
rect 880 74592 89120 74600
rect 880 74320 89963 74592
rect 13 73920 89963 74320
rect 13 73648 89120 73920
rect 880 73640 89120 73648
rect 880 73368 89963 73640
rect 13 73104 89963 73368
rect 13 72824 89120 73104
rect 13 72696 89963 72824
rect 880 72416 89963 72696
rect 13 72288 89963 72416
rect 13 72008 89120 72288
rect 13 71880 89963 72008
rect 880 71600 89963 71880
rect 13 71336 89963 71600
rect 13 71056 89120 71336
rect 13 70928 89963 71056
rect 880 70648 89963 70928
rect 13 70520 89963 70648
rect 13 70240 89120 70520
rect 13 69976 89963 70240
rect 880 69696 89963 69976
rect 13 69568 89963 69696
rect 13 69288 89120 69568
rect 13 69160 89963 69288
rect 880 68880 89963 69160
rect 13 68752 89963 68880
rect 13 68472 89120 68752
rect 13 68208 89963 68472
rect 880 67928 89963 68208
rect 13 67800 89963 67928
rect 13 67520 89120 67800
rect 13 67256 89963 67520
rect 880 66984 89963 67256
rect 880 66976 89120 66984
rect 13 66704 89120 66976
rect 13 66304 89963 66704
rect 880 66168 89963 66304
rect 880 66024 89120 66168
rect 13 65888 89120 66024
rect 13 65488 89963 65888
rect 880 65216 89963 65488
rect 880 65208 89120 65216
rect 13 64936 89120 65208
rect 13 64536 89963 64936
rect 880 64400 89963 64536
rect 880 64256 89120 64400
rect 13 64120 89120 64256
rect 13 63584 89963 64120
rect 880 63448 89963 63584
rect 880 63304 89120 63448
rect 13 63168 89120 63304
rect 13 62768 89963 63168
rect 880 62632 89963 62768
rect 880 62488 89120 62632
rect 13 62352 89120 62488
rect 13 61816 89963 62352
rect 880 61680 89963 61816
rect 880 61536 89120 61680
rect 13 61400 89120 61536
rect 13 60864 89963 61400
rect 880 60584 89120 60864
rect 13 60048 89963 60584
rect 13 59912 89120 60048
rect 880 59768 89120 59912
rect 880 59632 89963 59768
rect 13 59096 89963 59632
rect 880 58816 89120 59096
rect 13 58280 89963 58816
rect 13 58144 89120 58280
rect 880 58000 89120 58144
rect 880 57864 89963 58000
rect 13 57328 89963 57864
rect 13 57192 89120 57328
rect 880 57048 89120 57192
rect 880 56912 89963 57048
rect 13 56512 89963 56912
rect 13 56240 89120 56512
rect 880 56232 89120 56240
rect 880 55960 89963 56232
rect 13 55560 89963 55960
rect 13 55424 89120 55560
rect 880 55280 89120 55424
rect 880 55144 89963 55280
rect 13 54744 89963 55144
rect 13 54472 89120 54744
rect 880 54464 89120 54472
rect 880 54192 89963 54464
rect 13 53928 89963 54192
rect 13 53648 89120 53928
rect 13 53520 89963 53648
rect 880 53240 89963 53520
rect 13 52976 89963 53240
rect 13 52704 89120 52976
rect 880 52696 89120 52704
rect 880 52424 89963 52696
rect 13 52160 89963 52424
rect 13 51880 89120 52160
rect 13 51752 89963 51880
rect 880 51472 89963 51752
rect 13 51208 89963 51472
rect 13 50928 89120 51208
rect 13 50800 89963 50928
rect 880 50520 89963 50800
rect 13 50392 89963 50520
rect 13 50112 89120 50392
rect 13 49848 89963 50112
rect 880 49568 89963 49848
rect 13 49440 89963 49568
rect 13 49160 89120 49440
rect 13 49032 89963 49160
rect 880 48752 89963 49032
rect 13 48624 89963 48752
rect 13 48344 89120 48624
rect 13 48080 89963 48344
rect 880 47808 89963 48080
rect 880 47800 89120 47808
rect 13 47528 89120 47800
rect 13 47128 89963 47528
rect 880 46856 89963 47128
rect 880 46848 89120 46856
rect 13 46576 89120 46848
rect 13 46312 89963 46576
rect 880 46040 89963 46312
rect 880 46032 89120 46040
rect 13 45760 89120 46032
rect 13 45360 89963 45760
rect 880 45088 89963 45360
rect 880 45080 89120 45088
rect 13 44808 89120 45080
rect 13 44408 89963 44808
rect 880 44272 89963 44408
rect 880 44128 89120 44272
rect 13 43992 89120 44128
rect 13 43456 89963 43992
rect 880 43320 89963 43456
rect 880 43176 89120 43320
rect 13 43040 89120 43176
rect 13 42640 89963 43040
rect 880 42504 89963 42640
rect 880 42360 89120 42504
rect 13 42224 89120 42360
rect 13 41688 89963 42224
rect 880 41408 89120 41688
rect 13 40736 89963 41408
rect 880 40456 89120 40736
rect 13 39920 89963 40456
rect 13 39784 89120 39920
rect 880 39640 89120 39784
rect 880 39504 89963 39640
rect 13 38968 89963 39504
rect 880 38688 89120 38968
rect 13 38152 89963 38688
rect 13 38016 89120 38152
rect 880 37872 89120 38016
rect 880 37736 89963 37872
rect 13 37200 89963 37736
rect 13 37064 89120 37200
rect 880 36920 89120 37064
rect 880 36784 89963 36920
rect 13 36384 89963 36784
rect 13 36248 89120 36384
rect 880 36104 89120 36248
rect 880 35968 89963 36104
rect 13 35568 89963 35968
rect 13 35296 89120 35568
rect 880 35288 89120 35296
rect 880 35016 89963 35288
rect 13 34616 89963 35016
rect 13 34344 89120 34616
rect 880 34336 89120 34344
rect 880 34064 89963 34336
rect 13 33800 89963 34064
rect 13 33520 89120 33800
rect 13 33392 89963 33520
rect 880 33112 89963 33392
rect 13 32848 89963 33112
rect 13 32576 89120 32848
rect 880 32568 89120 32576
rect 880 32296 89963 32568
rect 13 32032 89963 32296
rect 13 31752 89120 32032
rect 13 31624 89963 31752
rect 880 31344 89963 31624
rect 13 31080 89963 31344
rect 13 30800 89120 31080
rect 13 30672 89963 30800
rect 880 30392 89963 30672
rect 13 30264 89963 30392
rect 13 29984 89120 30264
rect 13 29856 89963 29984
rect 880 29576 89963 29856
rect 13 29448 89963 29576
rect 13 29168 89120 29448
rect 13 28904 89963 29168
rect 880 28624 89963 28904
rect 13 28496 89963 28624
rect 13 28216 89120 28496
rect 13 27952 89963 28216
rect 880 27680 89963 27952
rect 880 27672 89120 27680
rect 13 27400 89120 27672
rect 13 27000 89963 27400
rect 880 26728 89963 27000
rect 880 26720 89120 26728
rect 13 26448 89120 26720
rect 13 26184 89963 26448
rect 880 25912 89963 26184
rect 880 25904 89120 25912
rect 13 25632 89120 25904
rect 13 25232 89963 25632
rect 880 24960 89963 25232
rect 880 24952 89120 24960
rect 13 24680 89120 24952
rect 13 24280 89963 24680
rect 880 24144 89963 24280
rect 880 24000 89120 24144
rect 13 23864 89120 24000
rect 13 23464 89963 23864
rect 880 23328 89963 23464
rect 880 23184 89120 23328
rect 13 23048 89120 23184
rect 13 22512 89963 23048
rect 880 22376 89963 22512
rect 880 22232 89120 22376
rect 13 22096 89120 22232
rect 13 21560 89963 22096
rect 880 21280 89120 21560
rect 13 20608 89963 21280
rect 880 20328 89120 20608
rect 13 19792 89963 20328
rect 880 19512 89120 19792
rect 13 18840 89963 19512
rect 880 18560 89120 18840
rect 13 18024 89963 18560
rect 13 17888 89120 18024
rect 880 17744 89120 17888
rect 880 17608 89963 17744
rect 13 17208 89963 17608
rect 13 16936 89120 17208
rect 880 16928 89120 16936
rect 880 16656 89963 16928
rect 13 16256 89963 16656
rect 13 16120 89120 16256
rect 880 15976 89120 16120
rect 880 15840 89963 15976
rect 13 15440 89963 15840
rect 13 15168 89120 15440
rect 880 15160 89120 15168
rect 880 14888 89963 15160
rect 13 14488 89963 14888
rect 13 14216 89120 14488
rect 880 14208 89120 14216
rect 880 13936 89963 14208
rect 13 13672 89963 13936
rect 13 13400 89120 13672
rect 880 13392 89120 13400
rect 880 13120 89963 13392
rect 13 12720 89963 13120
rect 13 12448 89120 12720
rect 880 12440 89120 12448
rect 880 12168 89963 12440
rect 13 11904 89963 12168
rect 13 11624 89120 11904
rect 13 11496 89963 11624
rect 880 11216 89963 11496
rect 13 11088 89963 11216
rect 13 10808 89120 11088
rect 13 10544 89963 10808
rect 880 10264 89963 10544
rect 13 10136 89963 10264
rect 13 9856 89120 10136
rect 13 9728 89963 9856
rect 880 9448 89963 9728
rect 13 9320 89963 9448
rect 13 9040 89120 9320
rect 13 8776 89963 9040
rect 880 8496 89963 8776
rect 13 8368 89963 8496
rect 13 8088 89120 8368
rect 13 7824 89963 8088
rect 880 7552 89963 7824
rect 880 7544 89120 7552
rect 13 7272 89120 7544
rect 13 7008 89963 7272
rect 880 6728 89963 7008
rect 13 6600 89963 6728
rect 13 6320 89120 6600
rect 13 6056 89963 6320
rect 880 5784 89963 6056
rect 880 5776 89120 5784
rect 13 5504 89120 5776
rect 13 5104 89963 5504
rect 880 4968 89963 5104
rect 880 4824 89120 4968
rect 13 4688 89120 4824
rect 13 4152 89963 4688
rect 880 4016 89963 4152
rect 880 3872 89120 4016
rect 13 3736 89120 3872
rect 13 3336 89963 3736
rect 880 3200 89963 3336
rect 880 3056 89120 3200
rect 13 2920 89120 3056
rect 13 2384 89963 2920
rect 880 2248 89963 2384
rect 880 2104 89120 2248
rect 13 1968 89120 2104
rect 13 1432 89963 1968
rect 880 1152 89120 1432
rect 13 616 89963 1152
rect 880 443 89120 616
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
<< obsm4 >>
rect 59 2483 4128 176765
rect 4608 2483 19488 176765
rect 19968 2483 34848 176765
rect 35328 2483 50208 176765
rect 50688 2483 65568 176765
rect 66048 2483 80928 176765
rect 81408 2483 89917 176765
<< labels >>
rlabel metal3 s 0 11296 800 11416 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 115472 800 115592 6 addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 117376 800 117496 6 addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 clk0
port 19 nsew signal output
rlabel metal3 s 0 107312 800 107432 6 clk1
port 20 nsew signal output
rlabel metal2 s 1030 179200 1086 180000 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 3146 179200 3202 180000 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 5262 179200 5318 180000 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 7378 179200 7434 180000 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 9586 179200 9642 180000 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 11702 179200 11758 180000 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 13818 179200 13874 180000 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 16026 179200 16082 180000 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 89200 2048 90000 2168 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 89200 7352 90000 7472 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 89200 37000 90000 37120 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 89200 39720 90000 39840 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 89200 42304 90000 42424 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 89200 44888 90000 45008 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 89200 47608 90000 47728 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 89200 50192 90000 50312 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 89200 52776 90000 52896 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 89200 55360 90000 55480 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 89200 58080 90000 58200 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 89200 60664 90000 60784 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 89200 10888 90000 11008 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 89200 63248 90000 63368 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 89200 65968 90000 66088 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 89200 68552 90000 68672 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 89200 71136 90000 71256 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 89200 73720 90000 73840 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 89200 76440 90000 76560 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 89200 79024 90000 79144 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 89200 81608 90000 81728 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 89200 14288 90000 14408 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 89200 17824 90000 17944 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 89200 21360 90000 21480 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 89200 23944 90000 24064 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 89200 26528 90000 26648 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 89200 29248 90000 29368 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 89200 31832 90000 31952 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 89200 34416 90000 34536 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 89200 3000 90000 3120 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 89200 8168 90000 8288 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 89200 37952 90000 38072 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 89200 40536 90000 40656 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 89200 43120 90000 43240 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 89200 45840 90000 45960 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 89200 48424 90000 48544 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 89200 51008 90000 51128 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 89200 53728 90000 53848 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 89200 56312 90000 56432 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 89200 58896 90000 59016 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 89200 61480 90000 61600 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 89200 11704 90000 11824 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 89200 64200 90000 64320 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 89200 66784 90000 66904 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 89200 69368 90000 69488 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 89200 72088 90000 72208 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 89200 74672 90000 74792 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 89200 77256 90000 77376 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 89200 79840 90000 79960 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 89200 82560 90000 82680 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 89200 84328 90000 84448 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 89200 85960 90000 86080 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 89200 15240 90000 15360 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 89200 87728 90000 87848 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 89200 89496 90000 89616 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 89200 18640 90000 18760 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 89200 22176 90000 22296 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 89200 24760 90000 24880 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 89200 27480 90000 27600 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 89200 30064 90000 30184 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 89200 32648 90000 32768 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 89200 35368 90000 35488 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 89200 9120 90000 9240 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 89200 38768 90000 38888 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 89200 41488 90000 41608 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 89200 44072 90000 44192 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 89200 46656 90000 46776 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 89200 49240 90000 49360 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 89200 51960 90000 52080 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 89200 54544 90000 54664 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 89200 57128 90000 57248 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 89200 59848 90000 59968 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 89200 62432 90000 62552 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 89200 12520 90000 12640 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 89200 65016 90000 65136 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 89200 67600 90000 67720 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 89200 70320 90000 70440 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 89200 72904 90000 73024 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 89200 75488 90000 75608 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 89200 78208 90000 78328 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 89200 80792 90000 80912 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 89200 83376 90000 83496 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 89200 85144 90000 85264 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 89200 86912 90000 87032 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 89200 16056 90000 16176 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 89200 88680 90000 88800 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 89200 90448 90000 90568 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 89200 19592 90000 19712 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 89200 23128 90000 23248 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 89200 25712 90000 25832 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 89200 28296 90000 28416 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 89200 30880 90000 31000 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 89200 33600 90000 33720 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 89200 36184 90000 36304 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 89200 3816 90000 3936 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 89200 9936 90000 10056 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 89200 13472 90000 13592 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 89200 17008 90000 17128 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 89200 20408 90000 20528 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 89200 4768 90000 4888 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 89200 5584 90000 5704 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 89200 6400 90000 6520 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 csb1[1]
port 134 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 din0[0]
port 135 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 din0[10]
port 136 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 din0[11]
port 137 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 din0[12]
port 138 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 din0[13]
port 139 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 din0[14]
port 140 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 din0[15]
port 141 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 din0[16]
port 142 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 din0[17]
port 143 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 din0[18]
port 144 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 din0[19]
port 145 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 din0[1]
port 146 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 din0[20]
port 147 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 din0[21]
port 148 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 din0[22]
port 149 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 din0[23]
port 150 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 din0[24]
port 151 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 din0[25]
port 152 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 din0[26]
port 153 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 din0[27]
port 154 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 din0[28]
port 155 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 din0[29]
port 156 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 din0[2]
port 157 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 din0[30]
port 158 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 din0[31]
port 159 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 din0[3]
port 160 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 din0[4]
port 161 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 din0[5]
port 162 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 din0[6]
port 163 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 din0[7]
port 164 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 din0[8]
port 165 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 din0[9]
port 166 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 dout0[0]
port 167 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 dout0[10]
port 168 nsew signal input
rlabel metal3 s 0 58896 800 59016 6 dout0[11]
port 169 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 dout0[12]
port 170 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 dout0[13]
port 171 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 dout0[15]
port 173 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 dout0[17]
port 175 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 dout0[18]
port 176 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 dout0[1]
port 178 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 dout0[20]
port 179 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 dout0[21]
port 180 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 dout0[22]
port 181 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 dout0[23]
port 182 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 dout0[24]
port 183 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 dout0[25]
port 184 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 dout0[26]
port 185 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 dout0[27]
port 186 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 dout0[29]
port 188 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 dout0[32]
port 192 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 dout0[33]
port 193 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 dout0[34]
port 194 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 dout0[35]
port 195 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 dout0[36]
port 196 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 dout0[37]
port 197 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 dout0[38]
port 198 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 dout0[39]
port 199 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 dout0[3]
port 200 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 dout0[40]
port 201 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 dout0[41]
port 202 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 dout0[42]
port 203 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 dout0[43]
port 204 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 dout0[44]
port 205 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 dout0[45]
port 206 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 dout0[46]
port 207 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 dout0[47]
port 208 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 dout0[48]
port 209 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 dout0[49]
port 210 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 dout0[4]
port 211 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 dout0[50]
port 212 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 dout0[51]
port 213 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 dout0[52]
port 214 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 dout0[53]
port 215 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 dout0[54]
port 216 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 dout0[55]
port 217 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 dout0[56]
port 218 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 dout0[57]
port 219 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 dout0[58]
port 220 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 dout0[59]
port 221 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 dout0[5]
port 222 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 dout0[60]
port 223 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 dout0[61]
port 224 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 dout0[62]
port 225 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 dout0[63]
port 226 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 dout0[6]
port 227 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 dout0[7]
port 228 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 dout0[8]
port 229 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 dout0[9]
port 230 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 dout1[0]
port 231 nsew signal input
rlabel metal3 s 0 127440 800 127560 6 dout1[10]
port 232 nsew signal input
rlabel metal3 s 0 128256 800 128376 6 dout1[11]
port 233 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 dout1[12]
port 234 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 dout1[13]
port 235 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 dout1[14]
port 236 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 dout1[15]
port 237 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 dout1[16]
port 238 nsew signal input
rlabel metal3 s 0 133832 800 133952 6 dout1[17]
port 239 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 dout1[18]
port 240 nsew signal input
rlabel metal3 s 0 135600 800 135720 6 dout1[19]
port 241 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 dout1[1]
port 242 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 dout1[20]
port 243 nsew signal input
rlabel metal3 s 0 137504 800 137624 6 dout1[21]
port 244 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 dout1[22]
port 245 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 dout1[23]
port 246 nsew signal input
rlabel metal3 s 0 140224 800 140344 6 dout1[24]
port 247 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 dout1[25]
port 248 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 dout1[26]
port 249 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 dout1[27]
port 250 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 dout1[28]
port 251 nsew signal input
rlabel metal3 s 0 144712 800 144832 6 dout1[29]
port 252 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 dout1[2]
port 253 nsew signal input
rlabel metal3 s 0 145664 800 145784 6 dout1[30]
port 254 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 dout1[31]
port 255 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 dout1[32]
port 256 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 dout1[33]
port 257 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 dout1[34]
port 258 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 dout1[35]
port 259 nsew signal input
rlabel metal3 s 0 151104 800 151224 6 dout1[36]
port 260 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 dout1[37]
port 261 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 dout1[38]
port 262 nsew signal input
rlabel metal3 s 0 153960 800 154080 6 dout1[39]
port 263 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 dout1[3]
port 264 nsew signal input
rlabel metal3 s 0 154776 800 154896 6 dout1[40]
port 265 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 dout1[41]
port 266 nsew signal input
rlabel metal3 s 0 156680 800 156800 6 dout1[42]
port 267 nsew signal input
rlabel metal3 s 0 157496 800 157616 6 dout1[43]
port 268 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 dout1[44]
port 269 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 dout1[45]
port 270 nsew signal input
rlabel metal3 s 0 160352 800 160472 6 dout1[46]
port 271 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 dout1[47]
port 272 nsew signal input
rlabel metal3 s 0 162120 800 162240 6 dout1[48]
port 273 nsew signal input
rlabel metal3 s 0 163072 800 163192 6 dout1[49]
port 274 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 dout1[4]
port 275 nsew signal input
rlabel metal3 s 0 164024 800 164144 6 dout1[50]
port 276 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 dout1[51]
port 277 nsew signal input
rlabel metal3 s 0 165792 800 165912 6 dout1[52]
port 278 nsew signal input
rlabel metal3 s 0 166744 800 166864 6 dout1[53]
port 279 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 dout1[54]
port 280 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 dout1[55]
port 281 nsew signal input
rlabel metal3 s 0 169464 800 169584 6 dout1[56]
port 282 nsew signal input
rlabel metal3 s 0 170416 800 170536 6 dout1[57]
port 283 nsew signal input
rlabel metal3 s 0 171232 800 171352 6 dout1[58]
port 284 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 dout1[59]
port 285 nsew signal input
rlabel metal3 s 0 122816 800 122936 6 dout1[5]
port 286 nsew signal input
rlabel metal3 s 0 173136 800 173256 6 dout1[60]
port 287 nsew signal input
rlabel metal3 s 0 173952 800 174072 6 dout1[61]
port 288 nsew signal input
rlabel metal3 s 0 174904 800 175024 6 dout1[62]
port 289 nsew signal input
rlabel metal3 s 0 175856 800 175976 6 dout1[63]
port 290 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 dout1[6]
port 291 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 dout1[7]
port 292 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 dout1[8]
port 293 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 dout1[9]
port 294 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 irq[0]
port 295 nsew signal input
rlabel metal3 s 89200 177760 90000 177880 6 irq[10]
port 296 nsew signal input
rlabel metal2 s 88798 179200 88854 180000 6 irq[11]
port 297 nsew signal input
rlabel metal3 s 89200 178712 90000 178832 6 irq[12]
port 298 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 irq[13]
port 299 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 irq[14]
port 300 nsew signal input
rlabel metal3 s 89200 179528 90000 179648 6 irq[15]
port 301 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 irq[1]
port 302 nsew signal input
rlabel metal2 s 84566 179200 84622 180000 6 irq[2]
port 303 nsew signal input
rlabel metal3 s 89200 176944 90000 177064 6 irq[3]
port 304 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 irq[4]
port 305 nsew signal input
rlabel metal2 s 86682 179200 86738 180000 6 irq[5]
port 306 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 irq[6]
port 307 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 irq[7]
port 308 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 irq[8]
port 309 nsew signal input
rlabel metal3 s 0 178576 800 178696 6 irq[9]
port 310 nsew signal input
rlabel metal3 s 0 416 800 536 6 jtag_tck
port 311 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 jtag_tdi
port 312 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 jtag_tdo
port 313 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 jtag_tms
port 314 nsew signal input
rlabel metal3 s 89200 91264 90000 91384 6 localMemory_wb_ack_o
port 315 nsew signal output
rlabel metal3 s 89200 96432 90000 96552 6 localMemory_wb_adr_i[0]
port 316 nsew signal input
rlabel metal3 s 89200 126216 90000 126336 6 localMemory_wb_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 89200 128800 90000 128920 6 localMemory_wb_adr_i[11]
port 318 nsew signal input
rlabel metal3 s 89200 131520 90000 131640 6 localMemory_wb_adr_i[12]
port 319 nsew signal input
rlabel metal3 s 89200 134104 90000 134224 6 localMemory_wb_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 89200 136688 90000 136808 6 localMemory_wb_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 89200 139272 90000 139392 6 localMemory_wb_adr_i[15]
port 322 nsew signal input
rlabel metal3 s 89200 141992 90000 142112 6 localMemory_wb_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 89200 144576 90000 144696 6 localMemory_wb_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 89200 147160 90000 147280 6 localMemory_wb_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 89200 149880 90000 150000 6 localMemory_wb_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 89200 99968 90000 100088 6 localMemory_wb_adr_i[1]
port 327 nsew signal input
rlabel metal3 s 89200 152464 90000 152584 6 localMemory_wb_adr_i[20]
port 328 nsew signal input
rlabel metal3 s 89200 155048 90000 155168 6 localMemory_wb_adr_i[21]
port 329 nsew signal input
rlabel metal3 s 89200 157632 90000 157752 6 localMemory_wb_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 89200 160352 90000 160472 6 localMemory_wb_adr_i[23]
port 331 nsew signal input
rlabel metal3 s 89200 103504 90000 103624 6 localMemory_wb_adr_i[2]
port 332 nsew signal input
rlabel metal3 s 89200 107040 90000 107160 6 localMemory_wb_adr_i[3]
port 333 nsew signal input
rlabel metal3 s 89200 110440 90000 110560 6 localMemory_wb_adr_i[4]
port 334 nsew signal input
rlabel metal3 s 89200 113160 90000 113280 6 localMemory_wb_adr_i[5]
port 335 nsew signal input
rlabel metal3 s 89200 115744 90000 115864 6 localMemory_wb_adr_i[6]
port 336 nsew signal input
rlabel metal3 s 89200 118328 90000 118448 6 localMemory_wb_adr_i[7]
port 337 nsew signal input
rlabel metal3 s 89200 120912 90000 121032 6 localMemory_wb_adr_i[8]
port 338 nsew signal input
rlabel metal3 s 89200 123632 90000 123752 6 localMemory_wb_adr_i[9]
port 339 nsew signal input
rlabel metal3 s 89200 92080 90000 92200 6 localMemory_wb_cyc_i
port 340 nsew signal input
rlabel metal3 s 89200 97384 90000 97504 6 localMemory_wb_data_i[0]
port 341 nsew signal input
rlabel metal3 s 89200 127032 90000 127152 6 localMemory_wb_data_i[10]
port 342 nsew signal input
rlabel metal3 s 89200 129752 90000 129872 6 localMemory_wb_data_i[11]
port 343 nsew signal input
rlabel metal3 s 89200 132336 90000 132456 6 localMemory_wb_data_i[12]
port 344 nsew signal input
rlabel metal3 s 89200 134920 90000 135040 6 localMemory_wb_data_i[13]
port 345 nsew signal input
rlabel metal3 s 89200 137640 90000 137760 6 localMemory_wb_data_i[14]
port 346 nsew signal input
rlabel metal3 s 89200 140224 90000 140344 6 localMemory_wb_data_i[15]
port 347 nsew signal input
rlabel metal3 s 89200 142808 90000 142928 6 localMemory_wb_data_i[16]
port 348 nsew signal input
rlabel metal3 s 89200 145392 90000 145512 6 localMemory_wb_data_i[17]
port 349 nsew signal input
rlabel metal3 s 89200 148112 90000 148232 6 localMemory_wb_data_i[18]
port 350 nsew signal input
rlabel metal3 s 89200 150696 90000 150816 6 localMemory_wb_data_i[19]
port 351 nsew signal input
rlabel metal3 s 89200 100920 90000 101040 6 localMemory_wb_data_i[1]
port 352 nsew signal input
rlabel metal3 s 89200 153280 90000 153400 6 localMemory_wb_data_i[20]
port 353 nsew signal input
rlabel metal3 s 89200 156000 90000 156120 6 localMemory_wb_data_i[21]
port 354 nsew signal input
rlabel metal3 s 89200 158584 90000 158704 6 localMemory_wb_data_i[22]
port 355 nsew signal input
rlabel metal3 s 89200 161168 90000 161288 6 localMemory_wb_data_i[23]
port 356 nsew signal input
rlabel metal3 s 89200 162936 90000 163056 6 localMemory_wb_data_i[24]
port 357 nsew signal input
rlabel metal3 s 89200 164704 90000 164824 6 localMemory_wb_data_i[25]
port 358 nsew signal input
rlabel metal3 s 89200 166472 90000 166592 6 localMemory_wb_data_i[26]
port 359 nsew signal input
rlabel metal3 s 89200 168240 90000 168360 6 localMemory_wb_data_i[27]
port 360 nsew signal input
rlabel metal3 s 89200 169872 90000 169992 6 localMemory_wb_data_i[28]
port 361 nsew signal input
rlabel metal3 s 89200 171640 90000 171760 6 localMemory_wb_data_i[29]
port 362 nsew signal input
rlabel metal3 s 89200 104320 90000 104440 6 localMemory_wb_data_i[2]
port 363 nsew signal input
rlabel metal3 s 89200 173408 90000 173528 6 localMemory_wb_data_i[30]
port 364 nsew signal input
rlabel metal3 s 89200 175176 90000 175296 6 localMemory_wb_data_i[31]
port 365 nsew signal input
rlabel metal3 s 89200 107856 90000 107976 6 localMemory_wb_data_i[3]
port 366 nsew signal input
rlabel metal3 s 89200 111392 90000 111512 6 localMemory_wb_data_i[4]
port 367 nsew signal input
rlabel metal3 s 89200 113976 90000 114096 6 localMemory_wb_data_i[5]
port 368 nsew signal input
rlabel metal3 s 89200 116560 90000 116680 6 localMemory_wb_data_i[6]
port 369 nsew signal input
rlabel metal3 s 89200 119280 90000 119400 6 localMemory_wb_data_i[7]
port 370 nsew signal input
rlabel metal3 s 89200 121864 90000 121984 6 localMemory_wb_data_i[8]
port 371 nsew signal input
rlabel metal3 s 89200 124448 90000 124568 6 localMemory_wb_data_i[9]
port 372 nsew signal input
rlabel metal3 s 89200 98200 90000 98320 6 localMemory_wb_data_o[0]
port 373 nsew signal output
rlabel metal3 s 89200 127984 90000 128104 6 localMemory_wb_data_o[10]
port 374 nsew signal output
rlabel metal3 s 89200 130568 90000 130688 6 localMemory_wb_data_o[11]
port 375 nsew signal output
rlabel metal3 s 89200 133152 90000 133272 6 localMemory_wb_data_o[12]
port 376 nsew signal output
rlabel metal3 s 89200 135872 90000 135992 6 localMemory_wb_data_o[13]
port 377 nsew signal output
rlabel metal3 s 89200 138456 90000 138576 6 localMemory_wb_data_o[14]
port 378 nsew signal output
rlabel metal3 s 89200 141040 90000 141160 6 localMemory_wb_data_o[15]
port 379 nsew signal output
rlabel metal3 s 89200 143760 90000 143880 6 localMemory_wb_data_o[16]
port 380 nsew signal output
rlabel metal3 s 89200 146344 90000 146464 6 localMemory_wb_data_o[17]
port 381 nsew signal output
rlabel metal3 s 89200 148928 90000 149048 6 localMemory_wb_data_o[18]
port 382 nsew signal output
rlabel metal3 s 89200 151512 90000 151632 6 localMemory_wb_data_o[19]
port 383 nsew signal output
rlabel metal3 s 89200 101736 90000 101856 6 localMemory_wb_data_o[1]
port 384 nsew signal output
rlabel metal3 s 89200 154232 90000 154352 6 localMemory_wb_data_o[20]
port 385 nsew signal output
rlabel metal3 s 89200 156816 90000 156936 6 localMemory_wb_data_o[21]
port 386 nsew signal output
rlabel metal3 s 89200 159400 90000 159520 6 localMemory_wb_data_o[22]
port 387 nsew signal output
rlabel metal3 s 89200 162120 90000 162240 6 localMemory_wb_data_o[23]
port 388 nsew signal output
rlabel metal3 s 89200 163752 90000 163872 6 localMemory_wb_data_o[24]
port 389 nsew signal output
rlabel metal3 s 89200 165520 90000 165640 6 localMemory_wb_data_o[25]
port 390 nsew signal output
rlabel metal3 s 89200 167288 90000 167408 6 localMemory_wb_data_o[26]
port 391 nsew signal output
rlabel metal3 s 89200 169056 90000 169176 6 localMemory_wb_data_o[27]
port 392 nsew signal output
rlabel metal3 s 89200 170824 90000 170944 6 localMemory_wb_data_o[28]
port 393 nsew signal output
rlabel metal3 s 89200 172592 90000 172712 6 localMemory_wb_data_o[29]
port 394 nsew signal output
rlabel metal3 s 89200 105272 90000 105392 6 localMemory_wb_data_o[2]
port 395 nsew signal output
rlabel metal3 s 89200 174360 90000 174480 6 localMemory_wb_data_o[30]
port 396 nsew signal output
rlabel metal3 s 89200 175992 90000 176112 6 localMemory_wb_data_o[31]
port 397 nsew signal output
rlabel metal3 s 89200 108672 90000 108792 6 localMemory_wb_data_o[3]
port 398 nsew signal output
rlabel metal3 s 89200 112208 90000 112328 6 localMemory_wb_data_o[4]
port 399 nsew signal output
rlabel metal3 s 89200 114792 90000 114912 6 localMemory_wb_data_o[5]
port 400 nsew signal output
rlabel metal3 s 89200 117512 90000 117632 6 localMemory_wb_data_o[6]
port 401 nsew signal output
rlabel metal3 s 89200 120096 90000 120216 6 localMemory_wb_data_o[7]
port 402 nsew signal output
rlabel metal3 s 89200 122680 90000 122800 6 localMemory_wb_data_o[8]
port 403 nsew signal output
rlabel metal3 s 89200 125400 90000 125520 6 localMemory_wb_data_o[9]
port 404 nsew signal output
rlabel metal3 s 89200 93032 90000 93152 6 localMemory_wb_error_o
port 405 nsew signal output
rlabel metal3 s 89200 99152 90000 99272 6 localMemory_wb_sel_i[0]
port 406 nsew signal input
rlabel metal3 s 89200 102552 90000 102672 6 localMemory_wb_sel_i[1]
port 407 nsew signal input
rlabel metal3 s 89200 106088 90000 106208 6 localMemory_wb_sel_i[2]
port 408 nsew signal input
rlabel metal3 s 89200 109624 90000 109744 6 localMemory_wb_sel_i[3]
port 409 nsew signal input
rlabel metal3 s 89200 93848 90000 93968 6 localMemory_wb_stall_o
port 410 nsew signal output
rlabel metal3 s 89200 94800 90000 94920 6 localMemory_wb_stb_i
port 411 nsew signal input
rlabel metal3 s 89200 95616 90000 95736 6 localMemory_wb_we_i
port 412 nsew signal input
rlabel metal2 s 18142 179200 18198 180000 6 manufacturerID[0]
port 413 nsew signal input
rlabel metal2 s 39578 179200 39634 180000 6 manufacturerID[10]
port 414 nsew signal input
rlabel metal2 s 20258 179200 20314 180000 6 manufacturerID[1]
port 415 nsew signal input
rlabel metal2 s 22374 179200 22430 180000 6 manufacturerID[2]
port 416 nsew signal input
rlabel metal2 s 24582 179200 24638 180000 6 manufacturerID[3]
port 417 nsew signal input
rlabel metal2 s 26698 179200 26754 180000 6 manufacturerID[4]
port 418 nsew signal input
rlabel metal2 s 28814 179200 28870 180000 6 manufacturerID[5]
port 419 nsew signal input
rlabel metal2 s 31022 179200 31078 180000 6 manufacturerID[6]
port 420 nsew signal input
rlabel metal2 s 33138 179200 33194 180000 6 manufacturerID[7]
port 421 nsew signal input
rlabel metal2 s 35254 179200 35310 180000 6 manufacturerID[8]
port 422 nsew signal input
rlabel metal2 s 37370 179200 37426 180000 6 manufacturerID[9]
port 423 nsew signal input
rlabel metal2 s 41694 179200 41750 180000 6 partID[0]
port 424 nsew signal input
rlabel metal2 s 63130 179200 63186 180000 6 partID[10]
port 425 nsew signal input
rlabel metal2 s 65246 179200 65302 180000 6 partID[11]
port 426 nsew signal input
rlabel metal2 s 67362 179200 67418 180000 6 partID[12]
port 427 nsew signal input
rlabel metal2 s 69570 179200 69626 180000 6 partID[13]
port 428 nsew signal input
rlabel metal2 s 71686 179200 71742 180000 6 partID[14]
port 429 nsew signal input
rlabel metal2 s 73802 179200 73858 180000 6 partID[15]
port 430 nsew signal input
rlabel metal2 s 43810 179200 43866 180000 6 partID[1]
port 431 nsew signal input
rlabel metal2 s 46018 179200 46074 180000 6 partID[2]
port 432 nsew signal input
rlabel metal2 s 48134 179200 48190 180000 6 partID[3]
port 433 nsew signal input
rlabel metal2 s 50250 179200 50306 180000 6 partID[4]
port 434 nsew signal input
rlabel metal2 s 52366 179200 52422 180000 6 partID[5]
port 435 nsew signal input
rlabel metal2 s 54574 179200 54630 180000 6 partID[6]
port 436 nsew signal input
rlabel metal2 s 56690 179200 56746 180000 6 partID[7]
port 437 nsew signal input
rlabel metal2 s 58806 179200 58862 180000 6 partID[8]
port 438 nsew signal input
rlabel metal2 s 61014 179200 61070 180000 6 partID[9]
port 439 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 probe_env[0]
port 440 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 probe_env[1]
port 441 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 probe_errorCode[0]
port 442 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 probe_errorCode[1]
port 443 nsew signal output
rlabel metal2 s 754 0 810 800 6 probe_isBranch
port 444 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 probe_isCompressed
port 445 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 probe_isLoad
port 446 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 probe_isStore
port 447 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 probe_jtagInstruction[0]
port 448 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 probe_jtagInstruction[1]
port 449 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 probe_jtagInstruction[2]
port 450 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 probe_jtagInstruction[3]
port 451 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 probe_jtagInstruction[4]
port 452 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 probe_opcode[0]
port 453 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 probe_opcode[1]
port 454 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 probe_opcode[2]
port 455 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 probe_opcode[3]
port 456 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 probe_opcode[4]
port 457 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 probe_opcode[5]
port 458 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 probe_opcode[6]
port 459 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 probe_programCounter[0]
port 460 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 probe_programCounter[10]
port 461 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 probe_programCounter[11]
port 462 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 probe_programCounter[12]
port 463 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 probe_programCounter[13]
port 464 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 probe_programCounter[14]
port 465 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 probe_programCounter[15]
port 466 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 probe_programCounter[16]
port 467 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 probe_programCounter[17]
port 468 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 probe_programCounter[18]
port 469 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 probe_programCounter[19]
port 470 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 probe_programCounter[1]
port 471 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 probe_programCounter[20]
port 472 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 probe_programCounter[21]
port 473 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 probe_programCounter[22]
port 474 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 probe_programCounter[23]
port 475 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 probe_programCounter[24]
port 476 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 probe_programCounter[25]
port 477 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 probe_programCounter[26]
port 478 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 probe_programCounter[27]
port 479 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 probe_programCounter[28]
port 480 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 probe_programCounter[29]
port 481 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 probe_programCounter[2]
port 482 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 probe_programCounter[30]
port 483 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 probe_programCounter[31]
port 484 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 probe_programCounter[3]
port 485 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 probe_programCounter[4]
port 486 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 probe_programCounter[5]
port 487 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 probe_programCounter[6]
port 488 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 probe_programCounter[7]
port 489 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 probe_programCounter[8]
port 490 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 probe_programCounter[9]
port 491 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 probe_state[0]
port 492 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 probe_state[1]
port 493 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 probe_takeBranch
port 494 nsew signal output
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 495 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 495 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 495 nsew power input
rlabel metal2 s 76010 179200 76066 180000 6 versionID[0]
port 496 nsew signal input
rlabel metal2 s 78126 179200 78182 180000 6 versionID[1]
port 497 nsew signal input
rlabel metal2 s 80242 179200 80298 180000 6 versionID[2]
port 498 nsew signal input
rlabel metal2 s 82358 179200 82414 180000 6 versionID[3]
port 499 nsew signal input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 500 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 500 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 500 nsew ground input
rlabel metal3 s 89200 416 90000 536 6 wb_clk_i
port 501 nsew signal input
rlabel metal3 s 89200 1232 90000 1352 6 wb_rst_i
port 502 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 web0
port 503 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 wmask0[0]
port 504 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 wmask0[1]
port 505 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 wmask0[2]
port 506 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 wmask0[3]
port 507 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 90000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 54922762
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/finishing/ExperiarCore.magic.gds
string GDS_START 1531032
<< end >>

