* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt CaravelHost caravel_irq[0] caravel_irq[1] caravel_irq[2] caravel_irq[3] caravel_uart_rx
+ caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0] caravel_wb_adr_o[10] caravel_wb_adr_o[11]
+ caravel_wb_adr_o[12] caravel_wb_adr_o[13] caravel_wb_adr_o[14] caravel_wb_adr_o[15]
+ caravel_wb_adr_o[16] caravel_wb_adr_o[17] caravel_wb_adr_o[18] caravel_wb_adr_o[19]
+ caravel_wb_adr_o[1] caravel_wb_adr_o[20] caravel_wb_adr_o[21] caravel_wb_adr_o[22]
+ caravel_wb_adr_o[23] caravel_wb_adr_o[24] caravel_wb_adr_o[25] caravel_wb_adr_o[26]
+ caravel_wb_adr_o[27] caravel_wb_adr_o[2] caravel_wb_adr_o[3] caravel_wb_adr_o[4]
+ caravel_wb_adr_o[5] caravel_wb_adr_o[6] caravel_wb_adr_o[7] caravel_wb_adr_o[8]
+ caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0] caravel_wb_data_i[10]
+ caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13] caravel_wb_data_i[14]
+ caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17] caravel_wb_data_i[18]
+ caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20] caravel_wb_data_i[21]
+ caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24] caravel_wb_data_i[25]
+ caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28] caravel_wb_data_i[29]
+ caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31] caravel_wb_data_i[3]
+ caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6] caravel_wb_data_i[7]
+ caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0] caravel_wb_data_o[10]
+ caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13] caravel_wb_data_o[14]
+ caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17] caravel_wb_data_o[18]
+ caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20] caravel_wb_data_o[21]
+ caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24] caravel_wb_data_o[25]
+ caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28] caravel_wb_data_o[29]
+ caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31] caravel_wb_data_o[3]
+ caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6] caravel_wb_data_o[7]
+ caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i caravel_wb_sel_o[0]
+ caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3] caravel_wb_stall_i caravel_wb_stb_o
+ caravel_wb_we_o core0Index[0] core0Index[1] core0Index[2] core0Index[3] core0Index[4]
+ core0Index[5] core0Index[6] core0Index[7] core1Index[0] core1Index[1] core1Index[2]
+ core1Index[3] core1Index[4] core1Index[5] core1Index[6] core1Index[7] manufacturerID[0]
+ manufacturerID[10] manufacturerID[1] manufacturerID[2] manufacturerID[3] manufacturerID[4]
+ manufacturerID[5] manufacturerID[6] manufacturerID[7] manufacturerID[8] manufacturerID[9]
+ partID[0] partID[10] partID[11] partID[12] partID[13] partID[14] partID[15] partID[1]
+ partID[2] partID[3] partID[4] partID[5] partID[6] partID[7] partID[8] partID[9]
+ vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12]
+ wbs_data_i[13] wbs_data_i[14] wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18]
+ wbs_data_i[19] wbs_data_i[1] wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23]
+ wbs_data_i[24] wbs_data_i[25] wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29]
+ wbs_data_i[2] wbs_data_i[30] wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5]
+ wbs_data_i[6] wbs_data_i[7] wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10]
+ wbs_data_o[11] wbs_data_o[12] wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16]
+ wbs_data_o[17] wbs_data_o[18] wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21]
+ wbs_data_o[22] wbs_data_o[23] wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27]
+ wbs_data_o[28] wbs_data_o[29] wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3]
+ wbs_data_o[4] wbs_data_o[5] wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7963_ _8483_/CLK _7963_/D vssd1 vssd1 vccd1 vccd1 _7963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7894_ _7894_/CLK _7894_/D vssd1 vssd1 vccd1 vccd1 _7894_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3626_ clkbuf_0__3626_/X vssd1 vssd1 vccd1 vccd1 _7434__9/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3988_ _3988_/A vssd1 vssd1 vccd1 vccd1 _8398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6776_ _8498_/Q _7473_/B vssd1 vssd1 vccd1 vccd1 _6777_/B sky130_fd_sc_hd__xor2_1
X_5727_ _5727_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5743_/S sky130_fd_sc_hd__nor2_2
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8446_ _8446_/CLK _8446_/D vssd1 vssd1 vccd1 vccd1 _8446_/Q sky130_fd_sc_hd__dfxtp_2
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _7903_/D sky130_fd_sc_hd__clkbuf_1
X_5589_ _5565_/X _7933_/Q _5593_/S vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__mux2_1
X_8377_ _8377_/CLK _8377_/D vssd1 vssd1 vccd1 vccd1 _8377_/Q sky130_fd_sc_hd__dfxtp_1
X_4609_ _4903_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _4610_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7328_ _8316_/Q _7337_/B vssd1 vssd1 vccd1 vccd1 _7328_/X sky130_fd_sc_hd__or2_1
XFILLER_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7065__542 _7068__545/A vssd1 vssd1 vccd1 vccd1 _8223_/CLK sky130_fd_sc_hd__inv_2
X_6848__389 _6849__390/A vssd1 vssd1 vccd1 vccd1 _8057_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7102__71 _7104__73/A vssd1 vssd1 vccd1 vccd1 _8252_/CLK sky130_fd_sc_hd__inv_2
X_6705__349 _6706__350/A vssd1 vssd1 vccd1 vccd1 _8013_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4960_/A vssd1 vssd1 vccd1 vccd1 _8111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4891_ _4789_/X _7856_/Q _4790_/X _8089_/Q _4663_/A vssd1 vssd1 vccd1 vccd1 _4891_/X
+ sky130_fd_sc_hd__o221a_1
X_3911_ _3911_/A vssd1 vssd1 vccd1 vccd1 _8460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _6973__468/A sky130_fd_sc_hd__clkbuf_4
X_3842_ _3842_/A _3842_/B _3842_/C _3842_/D vssd1 vssd1 vccd1 vccd1 _3843_/C sky130_fd_sc_hd__or4_1
X_6630_ _5915_/A _7962_/Q _6634_/S vssd1 vssd1 vccd1 vccd1 _6631_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5512_ _7987_/Q _4356_/A _5512_/S vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__mux2_1
X_8300_ _8315_/CLK _8300_/D vssd1 vssd1 vccd1 vccd1 _8300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6675__325/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8231_ _8231_/CLK _8231_/D vssd1 vssd1 vccd1 vccd1 _8231_/Q sky130_fd_sc_hd__dfxtp_1
X_5443_ _5443_/A vssd1 vssd1 vccd1 vccd1 _8021_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3241_ _6604_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3241_/X sky130_fd_sc_hd__clkbuf_16
X_5374_ _5373_/X _8052_/Q _5374_/S vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__mux2_1
X_8162_ _8162_/CLK _8162_/D vssd1 vssd1 vccd1 vccd1 _8162_/Q sky130_fd_sc_hd__dfxtp_1
X_4325_ _4340_/S vssd1 vssd1 vccd1 vccd1 _4334_/S sky130_fd_sc_hd__buf_2
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8093_ _8093_/CLK _8093_/D vssd1 vssd1 vccd1 vccd1 _8093_/Q sky130_fd_sc_hd__dfxtp_1
X_4256_ _4256_/A vssd1 vssd1 vccd1 vccd1 _8285_/D sky130_fd_sc_hd__clkbuf_1
X_7044_ _7044_/A vssd1 vssd1 vccd1 vccd1 _7044_/X sky130_fd_sc_hd__buf_1
X_7644__50 _7644__50/A vssd1 vssd1 vccd1 vccd1 _8473_/CLK sky130_fd_sc_hd__inv_2
X_4187_ _4187_/A vssd1 vssd1 vccd1 vccd1 _8338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7946_ _7946_/CLK _7946_/D vssd1 vssd1 vccd1 vccd1 _7946_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7877_ _7877_/CLK _7877_/D vssd1 vssd1 vccd1 vccd1 _7877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6759_ _8421_/Q vssd1 vssd1 vccd1 vccd1 _6789_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8429_ _8430_/CLK _8429_/D vssd1 vssd1 vccd1 vccd1 _8429_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3439_ _7108_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3439_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3756_ clkbuf_0__3756_/X vssd1 vssd1 vccd1 vccd1 _7629__37/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7384__144 _7384__144/A vssd1 vssd1 vccd1 vccd1 _8355_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__3281_ clkbuf_0__3281_/X vssd1 vssd1 vccd1 vccd1 _6718__354/A sky130_fd_sc_hd__clkbuf_16
X_7618__28 _7619__29/A vssd1 vssd1 vccd1 vccd1 _8451_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _6892_/A vssd1 vssd1 vccd1 vccd1 _7598_/A sky130_fd_sc_hd__clkbuf_2
X_4110_ _8122_/Q vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__inv_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _8382_/Q _4018_/X _4043_/S vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _5992_/A vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__clkbuf_1
X_7800_ _7800_/CLK _7800_/D vssd1 vssd1 vccd1 vccd1 _7800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _7731_/CLK _7731_/D vssd1 vssd1 vccd1 vccd1 _7731_/Q sky130_fd_sc_hd__dfxtp_1
X_4943_ _4943_/A vssd1 vssd1 vccd1 vccd1 _8118_/D sky130_fd_sc_hd__clkbuf_1
X_7662_ _7662_/A vssd1 vssd1 vccd1 vccd1 _7662_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4874_ _7776_/Q _4814_/X _4794_/A _4873_/X vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__o22a_1
X_6613_ _6613_/A vssd1 vssd1 vccd1 vccd1 _7954_/D sky130_fd_sc_hd__clkbuf_1
X_3825_ _8071_/Q vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7593_ _8440_/Q _7595_/B vssd1 vssd1 vccd1 vccd1 _7593_/X sky130_fd_sc_hd__or2_1
X_6475_ _6294_/A _6474_/Y _6289_/A vssd1 vssd1 vccd1 vccd1 _6477_/B sky130_fd_sc_hd__o21ai_1
XFILLER_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8214_ _8214_/CLK _8214_/D vssd1 vssd1 vccd1 vccd1 _8214_/Q sky130_fd_sc_hd__dfxtp_1
X_5426_ _3889_/X _8028_/Q _5428_/S vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3224_ _6522_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3224_/X sky130_fd_sc_hd__clkbuf_16
X_5357_ _5568_/A vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3610_ clkbuf_0__3610_/X vssd1 vssd1 vccd1 vccd1 _7351__117/A sky130_fd_sc_hd__clkbuf_4
X_8145_ _8145_/CLK _8145_/D vssd1 vssd1 vccd1 vccd1 _8145_/Q sky130_fd_sc_hd__dfxtp_1
X_4308_ _8262_/Q _4177_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__mux2_1
X_5288_ _8365_/Q _5178_/X _5179_/X _8357_/Q _5037_/A vssd1 vssd1 vccd1 vccd1 _5288_/X
+ sky130_fd_sc_hd__o221a_1
XINSDIODE2_4 _7775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8076_ _8076_/CLK _8076_/D vssd1 vssd1 vccd1 vccd1 _8076_/Q sky130_fd_sc_hd__dfxtp_1
X_7257__111 _7259__113/A vssd1 vssd1 vccd1 vccd1 _8294_/CLK sky130_fd_sc_hd__inv_2
X_4239_ _8292_/Q _4238_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7929_ _7929_/CLK _7929_/D vssd1 vssd1 vccd1 vccd1 _7929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _8150_/Q _4431_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5211_ _5261_/S vssd1 vssd1 vccd1 vccd1 _5235_/S sky130_fd_sc_hd__buf_2
X_6191_ _6184_/X _7966_/Q _6186_/X _6188_/X _7755_/Q vssd1 vssd1 vccd1 vccd1 _7755_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5142_ _5062_/X _5141_/X _5278_/A vssd1 vssd1 vccd1 vccd1 _5142_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5073_ _5073_/A vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__buf_2
X_4024_ _4024_/A vssd1 vssd1 vccd1 vccd1 _8389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5975_ _5975_/A vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7714_ _7200_/A _7707_/C _7713_/X _6421_/X vssd1 vssd1 vccd1 vccd1 _8496_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4926_ _4932_/A _4926_/B vssd1 vssd1 vccd1 vccd1 _4926_/Y sky130_fd_sc_hd__nand2_1
X_4857_ _4757_/X _4855_/X _4856_/X vssd1 vssd1 vccd1 vccd1 _4857_/X sky130_fd_sc_hd__o21a_1
X_7645_ _7649_/A _7645_/B vssd1 vssd1 vccd1 vccd1 _8474_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7576_ _7576_/A vssd1 vssd1 vccd1 vccd1 _8433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4788_ _8154_/Q _4770_/X _4787_/X _8116_/Q vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__a22o_1
X_7011__499 _7012__500/A vssd1 vssd1 vccd1 vccd1 _8180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3239_ clkbuf_0__3239_/X vssd1 vssd1 vccd1 vccd1 _6595__303/A sky130_fd_sc_hd__clkbuf_4
X_6458_ _7846_/Q _7961_/Q _6466_/S vssd1 vssd1 vccd1 vccd1 _6459_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5409_ _5409_/A vssd1 vssd1 vccd1 vccd1 _8037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6389_ _8486_/Q vssd1 vssd1 vccd1 vccd1 _7683_/A sky130_fd_sc_hd__buf_2
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8128_ _8128_/CLK _8128_/D vssd1 vssd1 vccd1 vccd1 _8128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8059_ _8059_/CLK _8059_/D vssd1 vssd1 vccd1 vccd1 _8059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7081__54 _7082__55/A vssd1 vssd1 vccd1 vccd1 _8235_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6554__271 _6554__271/A vssd1 vssd1 vccd1 vccd1 _7911_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7136__99 _7136__99/A vssd1 vssd1 vccd1 vccd1 _8280_/CLK sky130_fd_sc_hd__inv_2
X_6927__434 _6928__435/A vssd1 vssd1 vccd1 vccd1 _8112_/CLK sky130_fd_sc_hd__inv_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5760_ _5760_/A vssd1 vssd1 vccd1 vccd1 _7857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5727_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5707_/S sky130_fd_sc_hd__nor2_2
X_4711_ _4663_/X _4710_/X _4644_/X vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7430_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7430_/X sky130_fd_sc_hd__buf_1
X_4642_ _4642_/A vssd1 vssd1 vccd1 vccd1 _4653_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7361_ _7392_/A vssd1 vssd1 vccd1 vccd1 _7361_/X sky130_fd_sc_hd__buf_1
X_4573_ _4573_/A vssd1 vssd1 vccd1 vccd1 _8158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7292_ _7292_/A _7292_/B vssd1 vssd1 vccd1 vccd1 _7292_/Y sky130_fd_sc_hd__nand2_1
X_6312_ _7654_/A _6312_/B vssd1 vssd1 vccd1 vccd1 _6352_/A sky130_fd_sc_hd__nor2_2
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6243_ _7600_/A _6242_/X _6482_/A vssd1 vssd1 vccd1 vccd1 _7321_/A sky130_fd_sc_hd__a21o_4
XFILLER_115_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7397__154 _7398__155/A vssd1 vssd1 vccd1 vccd1 _8365_/CLK sky130_fd_sc_hd__inv_2
X_6174_ _6167_/X _7955_/Q _6170_/X _6172_/X _7744_/Q vssd1 vssd1 vccd1 vccd1 _7744_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5125_ _8463_/Q _8024_/Q _7989_/Q _8455_/Q _5063_/X _5111_/X vssd1 vssd1 vccd1 vccd1
+ _5125_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3240_ clkbuf_0__3240_/X vssd1 vssd1 vccd1 vccd1 _6600__307/A sky130_fd_sc_hd__clkbuf_4
X_4007_ _8393_/Q _4006_/X _4011_/S vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5958_ _5958_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__and2_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _5727_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5777_/S sky130_fd_sc_hd__or2_2
Xclkbuf_0__3756_ _7627_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3756_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5889_ _7707_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__or2_1
X_6874__396 _6878__400/A vssd1 vssd1 vccd1 vccd1 _8072_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7559_ _7582_/A _7559_/B vssd1 vssd1 vccd1 vccd1 _7560_/A sky130_fd_sc_hd__and2_1
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3438_ clkbuf_0__3438_/X vssd1 vssd1 vccd1 vccd1 _7120_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clkbuf_opt_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029__513 _7029__513/A vssd1 vssd1 vccd1 vccd1 _8194_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6861_ _8438_/Q _6863_/B vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__and2_1
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5812_ _5812_/A vssd1 vssd1 vccd1 vccd1 _7785_/D sky130_fd_sc_hd__clkbuf_1
X_6792_ _6792_/A _7468_/B _7468_/C vssd1 vssd1 vccd1 vccd1 _6792_/X sky130_fd_sc_hd__and3_1
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5743_ _7864_/Q _5580_/A _5743_/S vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3610_ _7349_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3610_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8533__232 vssd1 vssd1 vccd1 vccd1 _8533__232/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
X_8462_ _8462_/CLK _8462_/D vssd1 vssd1 vccd1 vccd1 _8462_/Q sky130_fd_sc_hd__dfxtp_1
X_5674_ _5689_/S vssd1 vssd1 vccd1 vccd1 _5683_/S sky130_fd_sc_hd__buf_2
X_8393_ _8393_/CLK _8393_/D vssd1 vssd1 vccd1 vccd1 _8393_/Q sky130_fd_sc_hd__dfxtp_1
X_4625_ _4798_/A vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__clkbuf_2
X_4556_ _4556_/A vssd1 vssd1 vccd1 vccd1 _8165_/D sky130_fd_sc_hd__clkbuf_1
X_7344_ _8086_/Q _7324_/A _7326_/A _7343_/X _7331_/A vssd1 vssd1 vccd1 vccd1 _8323_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_116_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_5_0_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_4487_ _4487_/A vssd1 vssd1 vccd1 vccd1 _8194_/D sky130_fd_sc_hd__clkbuf_1
X_7275_ _7282_/A _7275_/B vssd1 vssd1 vccd1 vccd1 _8299_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6226_ _7774_/Q _6225_/X _6480_/A vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__o21a_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6482_/A sky130_fd_sc_hd__buf_2
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5108_ _5108_/A vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__buf_2
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6088_ _7827_/Q input13/X _6107_/A vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__mux2_1
X_5039_ _5196_/S vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__buf_2
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3223_ clkbuf_0__3223_/X vssd1 vssd1 vccd1 vccd1 _6518__242/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8517__216 vssd1 vssd1 vccd1 vccd1 _8517__216/HI core0Index[3] sky130_fd_sc_hd__conb_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7348__115 _7348__115/A vssd1 vssd1 vccd1 vccd1 _8326_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6261__197 _6263__199/A vssd1 vssd1 vccd1 vccd1 _7789_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4410_ _8066_/Q vssd1 vssd1 vccd1 vccd1 _4410_/X sky130_fd_sc_hd__clkbuf_2
X_5390_ _5369_/X _8045_/Q _5392_/S vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _4341_/A vssd1 vssd1 vccd1 vccd1 _8247_/D sky130_fd_sc_hd__clkbuf_1
X_4272_ _4272_/A vssd1 vssd1 vccd1 vccd1 _8278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6011_ _7808_/Q input3/X _6123_/B vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6567__281 _6569__283/A vssd1 vssd1 vccd1 vccd1 _7921_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7962_ _7964_/CLK _7962_/D vssd1 vssd1 vccd1 vccd1 _7962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7251__106 _7252__107/A vssd1 vssd1 vccd1 vccd1 _8289_/CLK sky130_fd_sc_hd__inv_2
X_7893_ _7893_/CLK _7893_/D vssd1 vssd1 vccd1 vccd1 _7893_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3625_ clkbuf_0__3625_/X vssd1 vssd1 vccd1 vccd1 _7426__2/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6844_ _6844_/A vssd1 vssd1 vccd1 vccd1 _6844_/X sky130_fd_sc_hd__buf_1
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ _3940_/X _8398_/Q _3989_/S vssd1 vssd1 vccd1 vccd1 _3988_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6775_ _7476_/B _7476_/C _6774_/A vssd1 vssd1 vccd1 vccd1 _6775_/Y sky130_fd_sc_hd__a21oi_1
X_5726_ _5726_/A vssd1 vssd1 vccd1 vccd1 _7872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8445_ _8497_/CLK _8445_/D vssd1 vssd1 vccd1 vccd1 _8445_/Q sky130_fd_sc_hd__dfxtp_2
X_5657_ _5557_/X _7903_/Q _5665_/S vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__mux2_1
X_5588_ _5588_/A vssd1 vssd1 vccd1 vccd1 _7934_/D sky130_fd_sc_hd__clkbuf_1
X_8376_ _8376_/CLK _8376_/D vssd1 vssd1 vccd1 vccd1 _8376_/Q sky130_fd_sc_hd__dfxtp_1
X_4608_ _4608_/A _4608_/B vssd1 vssd1 vccd1 vccd1 _6938_/B sky130_fd_sc_hd__nor2_2
XFILLER_117_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4539_ _8172_/Q _4439_/X _4543_/S vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7327_ _7343_/B vssd1 vssd1 vccd1 vccd1 _7337_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6209_ _7597_/A _7765_/Q _6217_/S vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__mux2_1
X_7189_ _8303_/Q _7211_/A _7211_/B _7217_/A vssd1 vssd1 vccd1 vccd1 _7191_/A sky130_fd_sc_hd__nand4_1
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4890_ _4801_/X _7976_/Q _7880_/Q _4769_/X _4757_/A vssd1 vssd1 vccd1 vccd1 _4890_/X
+ sky130_fd_sc_hd__a221o_1
X_3910_ _8460_/Q _3886_/X _3914_/S vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _6012_/A vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__clkinv_4
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6560_ _6584_/A vssd1 vssd1 vccd1 vccd1 _6560_/X sky130_fd_sc_hd__buf_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5511_ _5511_/A vssd1 vssd1 vccd1 vccd1 _7988_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6667__318/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6491_ _6491_/A vssd1 vssd1 vccd1 vccd1 _6491_/X sky130_fd_sc_hd__buf_1
X_8230_ _8230_/CLK _8230_/D vssd1 vssd1 vccd1 vccd1 _8230_/Q sky130_fd_sc_hd__dfxtp_1
X_5442_ _8021_/Q _4448_/X _5446_/S vssd1 vssd1 vccd1 vccd1 _5443_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3240_ _6598_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3240_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5373_ _5580_/A vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8161_ _8161_/CLK _8161_/D vssd1 vssd1 vccd1 vccd1 _8161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4324_ _5466_/A _4343_/B vssd1 vssd1 vccd1 vccd1 _4340_/S sky130_fd_sc_hd__nor2_4
X_8092_ _8092_/CLK _8092_/D vssd1 vssd1 vccd1 vccd1 _8092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4255_ _8285_/Q _4182_/X _4261_/S vssd1 vssd1 vccd1 vccd1 _4256_/A sky130_fd_sc_hd__mux2_1
X_4186_ _8338_/Q _4185_/X _4192_/S vssd1 vssd1 vccd1 vccd1 _4187_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7945_ _7945_/CLK _7945_/D vssd1 vssd1 vccd1 vccd1 _7945_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7876_ _7876_/CLK _7876_/D vssd1 vssd1 vccd1 vccd1 _7876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6279__211 _6283__215/A vssd1 vssd1 vccd1 vccd1 _7803_/CLK sky130_fd_sc_hd__inv_2
X_6914__425 _6914__425/A vssd1 vssd1 vccd1 vccd1 _8103_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6758_ _7698_/A _7492_/B vssd1 vssd1 vccd1 vccd1 _6794_/A sky130_fd_sc_hd__nand2_1
X_6689_ _6701_/A vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__buf_1
X_5709_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5725_/S sky130_fd_sc_hd__or2_2
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8428_ _8430_/CLK _8428_/D vssd1 vssd1 vccd1 vccd1 _8428_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3438_ _7107_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3438_/X sky130_fd_sc_hd__clkbuf_16
X_8359_ _8359_/CLK _8359_/D vssd1 vssd1 vccd1 vccd1 _8359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3755_ clkbuf_0__3755_/X vssd1 vssd1 vccd1 vccd1 _7626__35/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921__429 _6922__430/A vssd1 vssd1 vccd1 vccd1 _8107_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7418__171 _7419__172/A vssd1 vssd1 vccd1 vccd1 _8382_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6518__242 _6518__242/A vssd1 vssd1 vccd1 vccd1 _7882_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4040_ _4040_/A vssd1 vssd1 vccd1 vccd1 _8383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5991_ _7965_/Q _5993_/B vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__and2_2
X_7730_ _7730_/CLK _7730_/D vssd1 vssd1 vccd1 vccd1 _7730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4942_ _8118_/Q _4232_/X _4946_/S vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__mux2_1
X_7661_ _5920_/A _7657_/X _7660_/Y vssd1 vssd1 vccd1 vccd1 _7661_/X sky130_fd_sc_hd__a21o_1
X_4873_ _4787_/A _7904_/Q _7896_/Q _4753_/A vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__a22o_1
X_6612_ _7693_/A _7954_/Q _6616_/S vssd1 vssd1 vccd1 vccd1 _6613_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7592_ _8440_/Q _7578_/A _7591_/X _7582_/X vssd1 vssd1 vccd1 vccd1 _8439_/D sky130_fd_sc_hd__o211a_1
X_3824_ _5018_/C _5018_/D _5018_/B vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6474_ _6228_/C _7675_/B _6412_/B vssd1 vssd1 vccd1 vccd1 _6474_/Y sky130_fd_sc_hd__a21oi_1
X_8213_ _8213_/CLK _8213_/D vssd1 vssd1 vccd1 vccd1 _8213_/Q sky130_fd_sc_hd__dfxtp_1
X_5425_ _5425_/A vssd1 vssd1 vccd1 vccd1 _8029_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3223_ _6516_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3223_/X sky130_fd_sc_hd__clkbuf_16
X_5356_ _8064_/Q vssd1 vssd1 vccd1 vccd1 _5568_/A sky130_fd_sc_hd__buf_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8144_ _8144_/CLK _8144_/D vssd1 vssd1 vccd1 vccd1 _8144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _4322_/S vssd1 vssd1 vccd1 vccd1 _4316_/S sky130_fd_sc_hd__buf_2
X_5287_ _8333_/Q _8341_/Q _5301_/S vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_5 _7775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8075_ _8075_/CLK _8075_/D vssd1 vssd1 vccd1 vccd1 _8075_/Q sky130_fd_sc_hd__dfxtp_1
X_7026_ _7026_/A vssd1 vssd1 vccd1 vccd1 _7026_/X sky130_fd_sc_hd__buf_1
X_4238_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__clkbuf_2
X_6727__361 _6728__362/A vssd1 vssd1 vccd1 vccd1 _8028_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4169_ _8344_/Q _4010_/X _4169_/S vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7928_ _7928_/CLK _7928_/D vssd1 vssd1 vccd1 vccd1 _7928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7859_ _7859_/CLK _7859_/D vssd1 vssd1 vccd1 vccd1 _7859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7023__508 _7024__509/A vssd1 vssd1 vccd1 vccd1 _8189_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7623__32 _7624__33/A vssd1 vssd1 vccd1 vccd1 _8455_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6490__220 _6490__220/A vssd1 vssd1 vccd1 vccd1 _7860_/CLK sky130_fd_sc_hd__inv_2
X_5210_ _5307_/S vssd1 vssd1 vccd1 vccd1 _5261_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6190_ _6184_/X _7965_/Q _6186_/X _6188_/X _7754_/Q vssd1 vssd1 vccd1 vccd1 _7754_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5141_ _8393_/Q _8385_/Q _7788_/Q _8401_/Q _5063_/X _5064_/X vssd1 vssd1 vccd1 vccd1
+ _5141_/X sky130_fd_sc_hd__mux4_1
X_5072_ _5152_/A _5072_/B vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__and2_1
X_4023_ _8389_/Q _4022_/X _4023_/S vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _5974_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__and2_1
X_7713_ _7607_/A _7707_/B _7704_/Y vssd1 vssd1 vccd1 vccd1 _7713_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _4925_/A vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4856_ _8184_/Q _4789_/X _4790_/X _8160_/Q _4715_/A vssd1 vssd1 vccd1 vccd1 _4856_/X
+ sky130_fd_sc_hd__o221a_1
X_7575_ _7575_/A _7575_/B _7575_/C vssd1 vssd1 vccd1 vccd1 _7576_/A sky130_fd_sc_hd__and3_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4787_ _4787_/A vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3238_ clkbuf_0__3238_/X vssd1 vssd1 vccd1 vccd1 _6598_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6457_ _6468_/A vssd1 vssd1 vccd1 vccd1 _6466_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5408_ _5369_/X _8037_/Q _5410_/S vssd1 vssd1 vccd1 vccd1 _5409_/A sky130_fd_sc_hd__mux2_1
X_6388_ _7820_/Q _6383_/X _6371_/X _6387_/X _6378_/X vssd1 vssd1 vccd1 vccd1 _7820_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5339_ _5044_/X _5331_/X _5338_/Y _5249_/X vssd1 vssd1 vccd1 vccd1 _8069_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8127_ _8127_/CLK _8127_/D vssd1 vssd1 vccd1 vccd1 _8127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8058_ _8058_/CLK _8058_/D vssd1 vssd1 vccd1 vccd1 _8058_/Q sky130_fd_sc_hd__dfxtp_1
X_6660__312 _6663__315/A vssd1 vssd1 vccd1 vccd1 _7976_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8550__249 vssd1 vssd1 vccd1 vccd1 _8550__249/HI versionID[3] sky130_fd_sc_hd__conb_1
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7439__13 _7439__13/A vssd1 vssd1 vccd1 vccd1 _8399_/CLK sky130_fd_sc_hd__inv_2
X_6966__462 _6968__464/A vssd1 vssd1 vccd1 vccd1 _8143_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6561__276 _6563__278/A vssd1 vssd1 vccd1 vccd1 _7916_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5690_ _5690_/A vssd1 vssd1 vccd1 vccd1 _7888_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _8094_/Q _7981_/Q _7885_/Q _7861_/Q _4630_/A _4633_/A vssd1 vssd1 vccd1 vccd1
+ _4710_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4641_ _8096_/Q _7983_/Q _7887_/Q _7863_/Q _4638_/X _4640_/X vssd1 vssd1 vccd1 vccd1
+ _4641_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4572_ _4404_/X _8158_/Q _4580_/S vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7291_ _7297_/A _7291_/B vssd1 vssd1 vccd1 vccd1 _8305_/D sky130_fd_sc_hd__nor2_1
X_6311_ _6311_/A vssd1 vssd1 vccd1 vccd1 _6311_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6242_ _6242_/A vssd1 vssd1 vccd1 vccd1 _6242_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173_ _6167_/X _7954_/Q _6170_/X _6172_/X _7743_/Q vssd1 vssd1 vccd1 vccd1 _7743_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_97_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5124_ _7797_/Q _8005_/Q _8284_/Q _8032_/Q _5241_/S _5052_/X vssd1 vssd1 vccd1 vccd1
+ _5124_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5055_ _5084_/B _5066_/B vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__or2_2
X_4006_ _4353_/A vssd1 vssd1 vccd1 vccd1 _4006_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5957_ _5957_/A vssd1 vssd1 vccd1 vccd1 _5957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3755_ _7621_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3755_/X sky130_fd_sc_hd__clkbuf_16
X_4908_ _4999_/A _4999_/B _4999_/C vssd1 vssd1 vccd1 vccd1 _5833_/B sky130_fd_sc_hd__nand3b_4
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _5888_/A vssd1 vssd1 vccd1 vccd1 _5888_/X sky130_fd_sc_hd__clkbuf_1
X_7627_ _7639_/A vssd1 vssd1 vccd1 vccd1 _7627_/X sky130_fd_sc_hd__buf_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839_ _4926_/B _4819_/X _4825_/X _4838_/X vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__a31o_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7558_ _8430_/Q _7510_/B _7556_/X _7557_/Y vssd1 vssd1 vccd1 vccd1 _7559_/B sky130_fd_sc_hd__a22o_1
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7489_ _8413_/Q vssd1 vssd1 vccd1 vccd1 _7508_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3437_ clkbuf_0__3437_/X vssd1 vssd1 vccd1 vccd1 _7106__75/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6667__318 _6667__318/A vssd1 vssd1 vccd1 vccd1 _7982_/CLK sky130_fd_sc_hd__inv_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _6860_/A vssd1 vssd1 vccd1 vccd1 _8063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5811_ _3889_/X _7785_/Q _5813_/S vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__mux2_1
X_6791_ _7468_/B _7468_/C _6792_/A vssd1 vssd1 vccd1 vccd1 _6791_/Y sky130_fd_sc_hd__a21oi_1
X_5742_ _5742_/A vssd1 vssd1 vccd1 vccd1 _7865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5673_ _5745_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5689_/S sky130_fd_sc_hd__nor2_2
X_8461_ _8461_/CLK _8461_/D vssd1 vssd1 vccd1 vccd1 _8461_/Q sky130_fd_sc_hd__dfxtp_1
X_8392_ _8392_/CLK _8392_/D vssd1 vssd1 vccd1 vccd1 _8392_/Q sky130_fd_sc_hd__dfxtp_1
X_4624_ _4766_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__or2_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6273__206 _6275__208/A vssd1 vssd1 vccd1 vccd1 _7798_/CLK sky130_fd_sc_hd__inv_2
X_4555_ _4410_/X _8165_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__mux2_1
X_7343_ _8323_/Q _7343_/B vssd1 vssd1 vccd1 vccd1 _7343_/X sky130_fd_sc_hd__or2_1
XFILLER_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4486_ _8194_/Q _4238_/X _4486_/S vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__mux2_1
X_7274_ _8299_/Q _7264_/X _7272_/X _7273_/Y vssd1 vssd1 vccd1 vccd1 _7275_/B sky130_fd_sc_hd__o2bb2a_1
X_6225_ _6008_/A _6423_/A _6016_/A _7773_/Q vssd1 vssd1 vccd1 vccd1 _6225_/X sky130_fd_sc_hd__a31o_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6146_/X _7767_/Q _6149_/X _6153_/X _7735_/Q vssd1 vssd1 vccd1 vccd1 _7735_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5105_/X _5106_/X _5186_/S vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _6072_/X _6084_/X _6086_/X _6075_/X vssd1 vssd1 vccd1 vccd1 _6087_/X sky130_fd_sc_hd__o211a_1
X_5038_ _5038_/A vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3222_ clkbuf_0__3222_/X vssd1 vssd1 vccd1 vccd1 _6514__239/A sky130_fd_sc_hd__clkbuf_4
X_7412__166 _7414__168/A vssd1 vssd1 vccd1 vccd1 _8377_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6989_ _6989_/A vssd1 vssd1 vccd1 vccd1 _6989_/X sky130_fd_sc_hd__buf_1
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6512__237 _6514__239/A vssd1 vssd1 vccd1 vccd1 _7877_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _8247_/Q _4200_/X _4340_/S vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__mux2_1
X_4271_ _8278_/Q _4177_/X _4279_/S vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7140__101 _7141__102/A vssd1 vssd1 vccd1 vccd1 _8282_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6061_/A vssd1 vssd1 vccd1 vccd1 _6123_/B sky130_fd_sc_hd__buf_4
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7961_ _8483_/CLK _7961_/D vssd1 vssd1 vccd1 vccd1 _7961_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7892_ _7892_/CLK _7892_/D vssd1 vssd1 vccd1 vccd1 _7892_/Q sky130_fd_sc_hd__dfxtp_1
X_6721__356 _6723__358/A vssd1 vssd1 vccd1 vccd1 _8023_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3624_ clkbuf_0__3624_/X vssd1 vssd1 vccd1 vccd1 _7448_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3986_ _3986_/A vssd1 vssd1 vccd1 vccd1 _8399_/D sky130_fd_sc_hd__clkbuf_1
X_6774_ _6774_/A _7476_/B _7476_/C vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__and3_1
X_5725_ _4156_/X _7872_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _5671_/S vssd1 vssd1 vccd1 vccd1 _5665_/S sky130_fd_sc_hd__buf_2
X_8444_ _8497_/CLK _8444_/D vssd1 vssd1 vccd1 vccd1 _8444_/Q sky130_fd_sc_hd__dfxtp_1
X_4607_ _4607_/A _4607_/B _4607_/C _4113_/B vssd1 vssd1 vccd1 vccd1 _4608_/B sky130_fd_sc_hd__or4b_2
X_5587_ _5562_/X _7934_/Q _5593_/S vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__mux2_1
X_8375_ _8375_/CLK _8375_/D vssd1 vssd1 vccd1 vccd1 _8375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4538_ _4538_/A vssd1 vssd1 vccd1 vccd1 _8173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7326_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7326_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ _4359_/X _8201_/Q _4473_/S vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__mux2_1
X_6208_ _6223_/S vssd1 vssd1 vccd1 vccd1 _6217_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7188_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _7471_/A sky130_fd_sc_hd__inv_2
XFILLER_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7354__120 _7354__120/A vssd1 vssd1 vccd1 vccd1 _8331_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7072__548 _7074__550/A vssd1 vssd1 vccd1 vccd1 _8229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _5328_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5510_ _7988_/Q _4353_/A _5512_/S vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5441_ _5441_/A vssd1 vssd1 vccd1 vccd1 _8022_/D sky130_fd_sc_hd__clkbuf_1
X_5372_ _8060_/Q vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__clkbuf_4
X_8160_ _8160_/CLK _8160_/D vssd1 vssd1 vccd1 vccd1 _8160_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _4323_/A vssd1 vssd1 vccd1 vccd1 _8255_/D sky130_fd_sc_hd__clkbuf_1
X_8091_ _8091_/CLK _8091_/D vssd1 vssd1 vccd1 vccd1 _8091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _4254_/A vssd1 vssd1 vccd1 vccd1 _8286_/D sky130_fd_sc_hd__clkbuf_1
X_4185_ _8447_/Q vssd1 vssd1 vccd1 vccd1 _4185_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7944_ _7944_/CLK _7944_/D vssd1 vssd1 vccd1 vccd1 _7944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _7875_/CLK _7875_/D vssd1 vssd1 vccd1 vccd1 _7875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6757_ _6757_/A _6757_/B vssd1 vssd1 vccd1 vccd1 _7492_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5708_ _5708_/A vssd1 vssd1 vccd1 vccd1 _7880_/D sky130_fd_sc_hd__clkbuf_1
X_3969_ _3969_/A vssd1 vssd1 vccd1 vccd1 _8405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5639_ _5557_/X _7911_/Q _5647_/S vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__mux2_1
X_8427_ _8430_/CLK _8427_/D vssd1 vssd1 vccd1 vccd1 _8427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3437_ _7101_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3437_/X sky130_fd_sc_hd__clkbuf_16
X_8358_ _8358_/CLK _8358_/D vssd1 vssd1 vccd1 vccd1 _8358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7309_ _7309_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _8312_/D sky130_fd_sc_hd__nor2_1
XFILLER_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8289_ _8289_/CLK _8289_/D vssd1 vssd1 vccd1 vccd1 _8289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5990_ _5990_/A vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4941_ _4941_/A vssd1 vssd1 vccd1 vccd1 _8119_/D sky130_fd_sc_hd__clkbuf_1
X_4872_ _4760_/X _7912_/Q _4814_/X _7920_/Q _4696_/S vssd1 vssd1 vccd1 vccd1 _4872_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0__f__3615_ clkbuf_0__3615_/X vssd1 vssd1 vccd1 vccd1 _7376__137/A sky130_fd_sc_hd__clkbuf_16
X_7660_ _8018_/Q _7704_/B vssd1 vssd1 vccd1 vccd1 _7660_/Y sky130_fd_sc_hd__nand2_2
X_3823_ _8074_/Q _8069_/Q vssd1 vssd1 vccd1 vccd1 _5018_/B sky130_fd_sc_hd__xnor2_1
X_6611_ _6611_/A vssd1 vssd1 vccd1 vccd1 _7953_/D sky130_fd_sc_hd__clkbuf_1
X_7591_ _8439_/Q _7595_/B vssd1 vssd1 vccd1 vccd1 _7591_/X sky130_fd_sc_hd__or2_1
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8141_/CLK sky130_fd_sc_hd__clkbuf_16
X_6473_ _6473_/A vssd1 vssd1 vccd1 vccd1 _7675_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8212_ _8212_/CLK _8212_/D vssd1 vssd1 vccd1 vccd1 _8212_/Q sky130_fd_sc_hd__dfxtp_1
X_5424_ _3886_/X _8029_/Q _5428_/S vssd1 vssd1 vccd1 vccd1 _5425_/A sky130_fd_sc_hd__mux2_1
Xoutput200 _6122_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
Xclkbuf_0__3222_ _6510_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3222_/X sky130_fd_sc_hd__clkbuf_16
X_8143_ _8143_/CLK _8143_/D vssd1 vssd1 vccd1 vccd1 _8143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5355_ _5355_/A vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_6 _4188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5286_ _8397_/Q _5163_/X _5295_/A _5284_/X _5285_/X vssd1 vssd1 vccd1 vccd1 _5286_/X
+ sky130_fd_sc_hd__o221a_1
X_4306_ _5779_/A _4343_/B vssd1 vssd1 vccd1 vccd1 _4322_/S sky130_fd_sc_hd__nor2_4
X_8074_ _8074_/CLK _8074_/D vssd1 vssd1 vccd1 vccd1 _8074_/Q sky130_fd_sc_hd__dfxtp_1
X_4237_ _4237_/A vssd1 vssd1 vccd1 vccd1 _8293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7093__64 _7094__65/A vssd1 vssd1 vccd1 vccd1 _8245_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4168_/A vssd1 vssd1 vccd1 vccd1 _8345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4099_ _8357_/Q _4022_/X _4099_/S vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7927_ _7927_/CLK _7927_/D vssd1 vssd1 vccd1 vccd1 _7927_/Q sky130_fd_sc_hd__dfxtp_1
X_7858_ _7858_/CLK _7858_/D vssd1 vssd1 vccd1 vccd1 _7858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6809_ _8425_/Q _6796_/A _6786_/B _6749_/A _8426_/Q vssd1 vssd1 vccd1 vccd1 _6810_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7789_ _7789_/CLK _7789_/D vssd1 vssd1 vccd1 vccd1 _7789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _8361_/Q _8345_/Q _8337_/Q _8369_/Q _5060_/X _5044_/X vssd1 vssd1 vccd1 vccd1
+ _5140_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5071_ _8473_/Q _8214_/Q _8206_/Q _8238_/Q _5060_/A _5070_/X vssd1 vssd1 vccd1 vccd1
+ _5072_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4022_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5973_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5982_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7712_ _7197_/A _7707_/C _7711_/X _6421_/X vssd1 vssd1 vccd1 vccd1 _8495_/D sky130_fd_sc_hd__o211a_1
X_4924_ _4924_/A vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7367__130 _7367__130/A vssd1 vssd1 vccd1 vccd1 _8341_/CLK sky130_fd_sc_hd__inv_2
X_4855_ _8152_/Q _4770_/X _4787_/X _8114_/Q vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4786_ _4777_/X _4779_/X _4785_/X _4673_/X vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__a211o_1
X_7574_ _8433_/Q _7556_/A vssd1 vssd1 vccd1 vccd1 _7575_/C sky130_fd_sc_hd__or2b_1
XFILLER_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3237_ clkbuf_0__3237_/X vssd1 vssd1 vccd1 vccd1 _6676_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6456_ _6456_/A vssd1 vssd1 vccd1 vccd1 _7845_/D sky130_fd_sc_hd__clkbuf_1
X_5407_ _5407_/A vssd1 vssd1 vccd1 vccd1 _8038_/D sky130_fd_sc_hd__clkbuf_1
X_6387_ _8487_/Q _6390_/B _6387_/C vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__and3_1
X_5338_ _5338_/A _5338_/B vssd1 vssd1 vccd1 vccd1 _5338_/Y sky130_fd_sc_hd__nand2_1
X_8126_ _8126_/CLK _8126_/D vssd1 vssd1 vccd1 vccd1 _8126_/Q sky130_fd_sc_hd__dfxtp_4
X_8057_ _8057_/CLK _8057_/D vssd1 vssd1 vccd1 vccd1 _8057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5269_ _7785_/Q _8382_/Q _5269_/S vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _4640_/A vssd1 vssd1 vccd1 vccd1 _4640_/X sky130_fd_sc_hd__buf_2
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6310_ _6310_/A _6310_/B vssd1 vssd1 vccd1 vccd1 _6311_/A sky130_fd_sc_hd__nor2_1
X_4571_ _4586_/S vssd1 vssd1 vccd1 vccd1 _4580_/S sky130_fd_sc_hd__buf_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7290_ _7184_/A _7280_/X _7286_/X _7289_/Y vssd1 vssd1 vccd1 vccd1 _7291_/B sky130_fd_sc_hd__o2bb2a_1
X_6241_ _8288_/Q _8287_/Q vssd1 vssd1 vccd1 vccd1 _7270_/A sky130_fd_sc_hd__nor2_2
X_6172_ _6172_/A vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__clkbuf_2
X_5123_ _5123_/A vssd1 vssd1 vccd1 vccd1 _5241_/S sky130_fd_sc_hd__buf_6
XFILLER_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5054_ _5054_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__nor2_1
X_4005_ _8446_/Q vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__buf_2
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5956_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__and2_1
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5887_ _7611_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__or2_1
X_4907_ _8130_/Q vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4838_ _4721_/X _4828_/X _4831_/X _4837_/X _4622_/A vssd1 vssd1 vccd1 vccd1 _4838_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4769_ _4769_/A vssd1 vssd1 vccd1 vccd1 _4769_/X sky130_fd_sc_hd__clkbuf_2
X_7557_ _7557_/A _7557_/B vssd1 vssd1 vccd1 vccd1 _7557_/Y sky130_fd_sc_hd__nor2_1
X_7488_ _8414_/Q vssd1 vssd1 vccd1 vccd1 _7504_/A sky130_fd_sc_hd__clkbuf_2
X_6439_ _6439_/A vssd1 vssd1 vccd1 vccd1 _7837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8109_ _8109_/CLK _8109_/D vssd1 vssd1 vccd1 vccd1 _8109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3436_ clkbuf_0__3436_/X vssd1 vssd1 vccd1 vccd1 _7098__68/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6940__444 _6941__445/A vssd1 vssd1 vccd1 vccd1 _8123_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_23_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8490_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7036__519 _7037__520/A vssd1 vssd1 vccd1 vccd1 _8200_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5810_ _5810_/A vssd1 vssd1 vccd1 vccd1 _7786_/D sky130_fd_sc_hd__clkbuf_1
X_6790_ _6789_/B _6789_/C _6789_/A vssd1 vssd1 vccd1 vccd1 _7468_/C sky130_fd_sc_hd__a21o_1
X_5741_ _7865_/Q _5577_/A _5743_/S vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8460_ _8460_/CLK _8460_/D vssd1 vssd1 vccd1 vccd1 _8460_/Q sky130_fd_sc_hd__dfxtp_1
X_5672_ _5672_/A vssd1 vssd1 vccd1 vccd1 _7896_/D sky130_fd_sc_hd__clkbuf_1
X_7411_ _7411_/A vssd1 vssd1 vccd1 vccd1 _7411_/X sky130_fd_sc_hd__buf_1
X_4623_ _4623_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__and2_1
X_8391_ _8391_/CLK _8391_/D vssd1 vssd1 vccd1 vccd1 _8391_/Q sky130_fd_sc_hd__dfxtp_1
X_4554_ _4554_/A vssd1 vssd1 vccd1 vccd1 _8166_/D sky130_fd_sc_hd__clkbuf_1
X_7342_ _8085_/Q _7324_/A _7326_/A _7341_/X _7331_/A vssd1 vssd1 vccd1 vccd1 _8322_/D
+ sky130_fd_sc_hd__o311a_1
X_7273_ _7273_/A _7273_/B vssd1 vssd1 vccd1 vccd1 _7273_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4485_ _4485_/A vssd1 vssd1 vccd1 vccd1 _8195_/D sky130_fd_sc_hd__clkbuf_1
X_6224_ _6224_/A vssd1 vssd1 vccd1 vccd1 _7772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6146_/X _7766_/Q _6149_/X _6153_/X _7734_/Q vssd1 vssd1 vccd1 vccd1 _7734_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5106_ _8261_/Q _8253_/Q _8245_/Q _8269_/Q _5078_/X _5070_/X vssd1 vssd1 vccd1 vccd1
+ _5106_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _7751_/Q _6111_/A vssd1 vssd1 vccd1 vccd1 _6086_/X sky130_fd_sc_hd__or2_1
X_5037_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3221_ clkbuf_0__3221_/X vssd1 vssd1 vccd1 vccd1 _6508__234/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _5939_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__or2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7609_ _7609_/A _7615_/B _7613_/C vssd1 vssd1 vccd1 vccd1 _7610_/A sky130_fd_sc_hd__and3_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput100 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _7699_/A sky130_fd_sc_hd__buf_4
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3419_ clkbuf_0__3419_/X vssd1 vssd1 vccd1 vccd1 _7038_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6673__323 _6675__325/A vssd1 vssd1 vccd1 vccd1 _7987_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _4285_/S vssd1 vssd1 vccd1 vccd1 _4279_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _8483_/CLK _7960_/D vssd1 vssd1 vccd1 vccd1 _7960_/Q sky130_fd_sc_hd__dfxtp_4
X_7891_ _7891_/CLK _7891_/D vssd1 vssd1 vccd1 vccd1 _7891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6979__473 _6979__473/A vssd1 vssd1 vccd1 vccd1 _8154_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3623_ clkbuf_0__3623_/X vssd1 vssd1 vccd1 vccd1 _7422__175/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _3937_/X _8399_/Q _3989_/S vssd1 vssd1 vccd1 vccd1 _3986_/A sky130_fd_sc_hd__mux2_1
X_6773_ _8416_/Q _7473_/B _6782_/B vssd1 vssd1 vccd1 vccd1 _7476_/C sky130_fd_sc_hd__a21o_1
X_5724_ _5724_/A vssd1 vssd1 vccd1 vccd1 _7873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5655_ _5655_/A _5815_/B vssd1 vssd1 vccd1 vccd1 _5671_/S sky130_fd_sc_hd__or2_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8443_ _8497_/CLK _8443_/D vssd1 vssd1 vccd1 vccd1 _8443_/Q sky130_fd_sc_hd__dfxtp_1
X_6574__287 _6574__287/A vssd1 vssd1 vccd1 vccd1 _7927_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8374_ _8374_/CLK _8374_/D vssd1 vssd1 vccd1 vccd1 _8374_/Q sky130_fd_sc_hd__dfxtp_1
X_4606_ _8141_/Q vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__clkbuf_2
X_5586_ _5586_/A vssd1 vssd1 vccd1 vccd1 _7935_/D sky130_fd_sc_hd__clkbuf_1
X_7325_ _7325_/A vssd1 vssd1 vccd1 vccd1 _7326_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4537_ _8173_/Q _4436_/X _4543_/S vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4468_ _4468_/A vssd1 vssd1 vccd1 vccd1 _8202_/D sky130_fd_sc_hd__clkbuf_1
X_7256_ _7349_/A vssd1 vssd1 vccd1 vccd1 _7256_/X sky130_fd_sc_hd__buf_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6207_ _6207_/A _6642_/B vssd1 vssd1 vccd1 vccd1 _6223_/S sky130_fd_sc_hd__nand2_2
X_7187_ _7289_/A _7289_/B _7698_/A vssd1 vssd1 vccd1 vccd1 _7187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4399_ _4399_/A vssd1 vssd1 vccd1 vccd1 _8225_/D sky130_fd_sc_hd__clkbuf_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6069_ _7822_/Q input8/X _6077_/S vssd1 vssd1 vccd1 vccd1 _6069_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8523__222 vssd1 vssd1 vccd1 vccd1 _8523__222/HI core1Index[2] sky130_fd_sc_hd__conb_1
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6824__370 _6824__370/A vssd1 vssd1 vccd1 vccd1 _8038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5440_ _8022_/Q _4445_/X _5440_/S vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371_ _5371_/A vssd1 vssd1 vccd1 vccd1 _8053_/D sky130_fd_sc_hd__clkbuf_1
X_4322_ _8255_/Q _4200_/X _4322_/S vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__mux2_1
X_8090_ _8090_/CLK _8090_/D vssd1 vssd1 vccd1 vccd1 _8090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _8286_/Q _4177_/X _4261_/S vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4184_ _4184_/A vssd1 vssd1 vccd1 vccd1 _8339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7943_ _7943_/CLK _7943_/D vssd1 vssd1 vccd1 vccd1 _7943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7874_ _7874_/CLK _7874_/D vssd1 vssd1 vccd1 vccd1 _7874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6825_ _6825_/A vssd1 vssd1 vccd1 vccd1 _6825_/X sky130_fd_sc_hd__buf_1
X_3968_ _8405_/Q _3892_/X _3968_/S vssd1 vssd1 vccd1 vccd1 _3969_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6756_ _6808_/B _6808_/C _8423_/Q vssd1 vssd1 vccd1 vccd1 _6757_/B sky130_fd_sc_hd__a21o_1
X_6953__454 _6954__455/A vssd1 vssd1 vccd1 vccd1 _8133_/CLK sky130_fd_sc_hd__inv_2
X_5707_ _7880_/Q _4996_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5708_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3899_ _3914_/S vssd1 vssd1 vccd1 vccd1 _3908_/S sky130_fd_sc_hd__buf_2
X_5638_ _5653_/S vssd1 vssd1 vccd1 vccd1 _5647_/S sky130_fd_sc_hd__buf_2
X_7049__529 _7050__530/A vssd1 vssd1 vccd1 vccd1 _8210_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3399_ clkbuf_0__3399_/X vssd1 vssd1 vccd1 vccd1 _7013_/A sky130_fd_sc_hd__clkbuf_4
X_8426_ _8430_/CLK _8426_/D vssd1 vssd1 vccd1 vccd1 _8426_/Q sky130_fd_sc_hd__dfxtp_1
X_5569_ _5568_/X _7940_/Q _5572_/S vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3436_ _7095_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3436_/X sky130_fd_sc_hd__clkbuf_16
X_8357_ _8357_/CLK _8357_/D vssd1 vssd1 vccd1 vccd1 _8357_/Q sky130_fd_sc_hd__dfxtp_1
X_7308_ _8312_/Q _7295_/A _7272_/A _7155_/B vssd1 vssd1 vccd1 vccd1 _7309_/B sky130_fd_sc_hd__o2bb2a_1
X_8288_ _8315_/CLK _8288_/D vssd1 vssd1 vccd1 vccd1 _8288_/Q sky130_fd_sc_hd__dfxtp_1
X_7239_ _7241_/A _7241_/B _7478_/A vssd1 vssd1 vccd1 vccd1 _7239_/X sky130_fd_sc_hd__a21bo_1
X_7635__42 _7635__42/A vssd1 vssd1 vccd1 vccd1 _8465_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6525__248 _6527__250/A vssd1 vssd1 vccd1 vccd1 _7888_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _8119_/Q _4229_/X _4946_/S vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__mux2_1
X_4871_ _4749_/X _7800_/Q _7725_/Q _4795_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4871_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6610_ _7696_/A _7953_/Q _6616_/S vssd1 vssd1 vccd1 vccd1 _6611_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7590_ _8439_/Q _7578_/X _7589_/X _7582_/X vssd1 vssd1 vccd1 vccd1 _8438_/D sky130_fd_sc_hd__o211a_1
X_3822_ _8073_/Q _8068_/Q vssd1 vssd1 vccd1 vccd1 _5018_/D sky130_fd_sc_hd__or2b_1
X_6541_ _6547_/A vssd1 vssd1 vccd1 vccd1 _6541_/X sky130_fd_sc_hd__buf_1
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6472_ _6472_/A vssd1 vssd1 vccd1 vccd1 _7852_/D sky130_fd_sc_hd__clkbuf_1
X_8211_ _8211_/CLK _8211_/D vssd1 vssd1 vccd1 vccd1 _8211_/Q sky130_fd_sc_hd__dfxtp_1
X_5423_ _5423_/A vssd1 vssd1 vccd1 vccd1 _8030_/D sky130_fd_sc_hd__clkbuf_1
Xoutput201 _6124_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
X_5354_ _5353_/X _8057_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3221_ _6504_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3221_/X sky130_fd_sc_hd__clkbuf_16
X_8142_ _8481_/CLK _8142_/D vssd1 vssd1 vccd1 vccd1 _8142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6686__333 _6688__335/A vssd1 vssd1 vccd1 vccd1 _7997_/CLK sky130_fd_sc_hd__inv_2
X_4305_ _4305_/A vssd1 vssd1 vccd1 vccd1 _8263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5285_ _8389_/Q _5285_/B vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__or2_1
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_7 _4359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8073_ _8073_/CLK _8073_/D vssd1 vssd1 vccd1 vccd1 _8073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4236_ _8293_/Q _4235_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__mux2_1
X_7078__51 _7079__52/A vssd1 vssd1 vccd1 vccd1 _8232_/CLK sky130_fd_sc_hd__inv_2
X_4167_ _8345_/Q _4006_/X _4169_/S vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _8358_/D sky130_fd_sc_hd__clkbuf_1
X_7926_ _7926_/CLK _7926_/D vssd1 vssd1 vccd1 vccd1 _7926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7857_ _7857_/CLK _7857_/D vssd1 vssd1 vccd1 vccd1 _7857_/Q sky130_fd_sc_hd__dfxtp_1
X_6808_ _6808_/A _6808_/B _6808_/C vssd1 vssd1 vccd1 vccd1 _6810_/A sky130_fd_sc_hd__nand3_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7788_ _7788_/CLK _7788_/D vssd1 vssd1 vccd1 vccd1 _7788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6739_ _8422_/Q _8421_/Q _8420_/Q _8419_/Q vssd1 vssd1 vccd1 vccd1 _6749_/A sky130_fd_sc_hd__and4_1
XFILLER_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6734__367 _6734__367/A vssd1 vssd1 vccd1 vccd1 _8034_/CLK sky130_fd_sc_hd__inv_2
X_8409_ _8409_/CLK _8409_/D vssd1 vssd1 vccd1 vccd1 _8409_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3419_ _7013_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3419_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6531__252 _6531__252/A vssd1 vssd1 vccd1 vccd1 _7892_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _5164_/A vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__buf_2
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4021_ _8442_/Q vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__buf_2
XFILLER_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5972_ _5972_/A vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7711_ _7609_/A _7707_/B _7704_/Y vssd1 vssd1 vccd1 vccd1 _7711_/X sky130_fd_sc_hd__a21o_1
X_4923_ _4923_/A _4923_/B vssd1 vssd1 vccd1 vccd1 _8127_/D sky130_fd_sc_hd__nor2_1
X_7429__5 _7429__5/A vssd1 vssd1 vccd1 vccd1 _8391_/CLK sky130_fd_sc_hd__inv_2
X_4854_ _4849_/X _4850_/X _4853_/X _4673_/X vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__a211o_1
XFILLER_60_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4785_ _8194_/Q _4765_/X _4661_/A _4784_/X vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__o211a_1
X_6837__380 _6837__380/A vssd1 vssd1 vccd1 vccd1 _8048_/CLK sky130_fd_sc_hd__inv_2
X_7573_ _6820_/C _7564_/Y _7572_/X _7556_/X vssd1 vssd1 vccd1 vccd1 _7575_/B sky130_fd_sc_hd__a211o_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3236_ clkbuf_0__3236_/X vssd1 vssd1 vccd1 vccd1 _6589__300/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6455_ _7845_/Q _7960_/Q _6455_/S vssd1 vssd1 vccd1 vccd1 _6456_/A sky130_fd_sc_hd__mux2_1
X_5406_ _5365_/X _8038_/Q _5410_/S vssd1 vssd1 vccd1 vccd1 _5407_/A sky130_fd_sc_hd__mux2_1
X_6386_ _7819_/Q _6383_/X _6371_/X _6385_/X _6378_/X vssd1 vssd1 vccd1 vccd1 _7819_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5337_ _5214_/X _5331_/X _5336_/Y _5249_/X vssd1 vssd1 vccd1 vccd1 _8070_/D sky130_fd_sc_hd__o211a_1
X_8125_ _8125_/CLK _8125_/D vssd1 vssd1 vccd1 vccd1 _8125_/Q sky130_fd_sc_hd__dfxtp_1
X_8056_ _8056_/CLK _8056_/D vssd1 vssd1 vccd1 vccd1 _8056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _5220_/X _5266_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _5268_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_85_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4219_ _8326_/Q _4153_/X _4221_/S vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__mux2_1
X_7007_ _7007_/A vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__buf_1
X_5199_ _8282_/Q _8003_/Q _5307_/S vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7909_ _7909_/CLK _7909_/D vssd1 vssd1 vccd1 vccd1 _7909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6973__468 _6973__468/A vssd1 vssd1 vccd1 vccd1 _8149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _5655_/A _4936_/A vssd1 vssd1 vccd1 vccd1 _4586_/S sky130_fd_sc_hd__or2_2
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6240_ _8315_/Q _6236_/X _6238_/X _7320_/C vssd1 vssd1 vccd1 vccd1 _6240_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6171_ _6167_/X _7953_/Q _6170_/X _6163_/X _7742_/Q vssd1 vssd1 vccd1 vccd1 _7742_/D
+ sky130_fd_sc_hd__o32a_1
X_5122_ _5038_/X _5119_/X _5121_/X vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__a21o_1
X_7445__18 _7445__18/A vssd1 vssd1 vccd1 vccd1 _8404_/CLK sky130_fd_sc_hd__inv_2
X_7431__6 _7432__7/A vssd1 vssd1 vccd1 vccd1 _8392_/CLK sky130_fd_sc_hd__inv_2
X_5053_ _8465_/Q _8026_/Q _7991_/Q _8457_/Q _5294_/S _5052_/X vssd1 vssd1 vccd1 vccd1
+ _5053_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4004_ _4004_/A vssd1 vssd1 vccd1 vccd1 _8394_/D sky130_fd_sc_hd__clkbuf_1
X_8503__253 vssd1 vssd1 vccd1 vccd1 partID[4] _8503__253/LO sky130_fd_sc_hd__conb_1
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5955_ _5955_/A vssd1 vssd1 vccd1 vccd1 _5955_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5886_ _5943_/B vssd1 vssd1 vccd1 vccd1 _5895_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4906_ _5709_/B vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__buf_2
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4837_ _4832_/X _4833_/X _4836_/X _4773_/A vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6538__258 _6539__259/A vssd1 vssd1 vccd1 vccd1 _7898_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4768_ _7947_/Q _4653_/B _4767_/X vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__a21o_1
X_7556_ _7556_/A vssd1 vssd1 vccd1 vccd1 _7556_/X sky130_fd_sc_hd__clkbuf_2
X_4699_ _4735_/A _4698_/X _4665_/A vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__a21o_1
X_7487_ _7487_/A _7487_/B _7487_/C _7487_/D vssd1 vssd1 vccd1 vccd1 _7490_/A sky130_fd_sc_hd__or4_2
XFILLER_107_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3219_ clkbuf_0__3219_/X vssd1 vssd1 vccd1 vccd1 _6522_/A sky130_fd_sc_hd__clkbuf_4
X_6438_ _7837_/Q _5963_/A _6444_/S vssd1 vssd1 vccd1 vccd1 _6439_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8108_ _8108_/CLK _8108_/D vssd1 vssd1 vccd1 vccd1 _8108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6369_ _6369_/A _6369_/B vssd1 vssd1 vccd1 vccd1 _6370_/A sky130_fd_sc_hd__or2_1
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8039_ _8039_/CLK _8039_/D vssd1 vssd1 vccd1 vccd1 _8039_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3435_ clkbuf_0__3435_/X vssd1 vssd1 vccd1 vccd1 _7092__63/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _7866_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5580_/X _7896_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5672_/A sky130_fd_sc_hd__mux2_1
X_8390_ _8390_/CLK _8390_/D vssd1 vssd1 vccd1 vccd1 _8390_/Q sky130_fd_sc_hd__dfxtp_1
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _4622_/X sky130_fd_sc_hd__clkbuf_2
X_4553_ _4404_/X _8166_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__mux2_1
X_7341_ _8322_/Q _7343_/B vssd1 vssd1 vccd1 vccd1 _7341_/X sky130_fd_sc_hd__or2_1
X_4484_ _8195_/Q _4235_/X _4486_/S vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__mux2_1
X_7272_ _7272_/A vssd1 vssd1 vccd1 vccd1 _7272_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6223_ _7615_/A _7772_/Q _6223_/S vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6154_ _6146_/X _7765_/Q _6149_/X _6153_/X _7733_/Q vssd1 vssd1 vccd1 vccd1 _7733_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _8379_/Q _8277_/Q _8014_/Q _8229_/Q _5111_/A _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5105_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6085_/A vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__buf_2
X_8540__239 vssd1 vssd1 vccd1 vccd1 _8540__239/HI partID[1] sky130_fd_sc_hd__conb_1
X_5036_ _5073_/A vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__buf_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3220_ clkbuf_0__3220_/X vssd1 vssd1 vccd1 vccd1 _6500__227/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5938_ _5938_/A vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _6006_/B vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7608_ _7608_/A vssd1 vssd1 vccd1 vccd1 _8445_/D sky130_fd_sc_hd__clkbuf_1
X_7539_ _7546_/A _7539_/B vssd1 vssd1 vccd1 vccd1 _8422_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _7696_/A sky130_fd_sc_hd__buf_4
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3418_ clkbuf_0__3418_/X vssd1 vssd1 vccd1 vccd1 _7009__497/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7000__490 _7000__490/A vssd1 vssd1 vccd1 vccd1 _8171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7042__524 _7043__525/A vssd1 vssd1 vccd1 vccd1 _8205_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6680__328 _6681__329/A vssd1 vssd1 vccd1 vccd1 _7992_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7890_ _7890_/CLK _7890_/D vssd1 vssd1 vccd1 vccd1 _7890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3622_ clkbuf_0__3622_/X vssd1 vssd1 vccd1 vccd1 _7414__168/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3984_ _3984_/A vssd1 vssd1 vccd1 vccd1 _8400_/D sky130_fd_sc_hd__clkbuf_1
X_6772_ _6782_/B _6782_/C _7473_/B vssd1 vssd1 vccd1 vccd1 _7476_/B sky130_fd_sc_hd__nand3_2
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5723_ _4153_/X _7873_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5654_ _5654_/A vssd1 vssd1 vccd1 vccd1 _7904_/D sky130_fd_sc_hd__clkbuf_1
X_8442_ _8442_/CLK _8442_/D vssd1 vssd1 vccd1 vccd1 _8442_/Q sky130_fd_sc_hd__dfxtp_2
X_8373_ _8373_/CLK _8373_/D vssd1 vssd1 vccd1 vccd1 _8373_/Q sky130_fd_sc_hd__dfxtp_1
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _8143_/D sky130_fd_sc_hd__clkbuf_1
X_5585_ _5557_/X _7935_/Q _5593_/S vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__mux2_1
X_7324_ _7324_/A vssd1 vssd1 vccd1 vccd1 _7648_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4536_ _4536_/A vssd1 vssd1 vccd1 vccd1 _8174_/D sky130_fd_sc_hd__clkbuf_1
X_6986__478 _6988__480/A vssd1 vssd1 vccd1 vccd1 _8159_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4467_ _4356_/X _8202_/Q _4467_/S vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__mux2_1
X_4398_ _4359_/X _8225_/Q _4402_/S vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__mux2_1
X_6206_ _6206_/A _6231_/B vssd1 vssd1 vccd1 vccd1 _6642_/B sky130_fd_sc_hd__nor2_4
X_7186_ _8491_/Q _7289_/A _7289_/B vssd1 vssd1 vccd1 vccd1 _7186_/X sky130_fd_sc_hd__and3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6068_ _6053_/X _6065_/X _6067_/X _6056_/X vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__o211a_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5019_ _5019_/A _5019_/B _5018_/X vssd1 vssd1 vccd1 vccd1 _6895_/C sky130_fd_sc_hd__or3b_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_4_0_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5370_ _5369_/X _8053_/Q _5374_/S vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4321_ _4321_/A vssd1 vssd1 vccd1 vccd1 _8256_/D sky130_fd_sc_hd__clkbuf_1
X_4252_ _4267_/S vssd1 vssd1 vccd1 vccd1 _4261_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4183_ _8339_/Q _4182_/X _4192_/S vssd1 vssd1 vccd1 vccd1 _4184_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7942_ _7942_/CLK _7942_/D vssd1 vssd1 vccd1 vccd1 _7942_/Q sky130_fd_sc_hd__dfxtp_1
X_6580__292 _6580__292/A vssd1 vssd1 vccd1 vccd1 _7932_/CLK sky130_fd_sc_hd__inv_2
X_7873_ _7873_/CLK _7873_/D vssd1 vssd1 vccd1 vccd1 _7873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3967_ _3967_/A vssd1 vssd1 vccd1 vccd1 _8406_/D sky130_fd_sc_hd__clkbuf_1
X_6755_ _8423_/Q _6808_/B _6808_/C vssd1 vssd1 vccd1 vccd1 _6757_/A sky130_fd_sc_hd__nand3_1
X_5706_ _5706_/A vssd1 vssd1 vccd1 vccd1 _7881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3898_ _4083_/A _5502_/A vssd1 vssd1 vccd1 vccd1 _3914_/S sky130_fd_sc_hd__nor2_2
X_8425_ _8425_/CLK _8425_/D vssd1 vssd1 vccd1 vccd1 _8425_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3398_ clkbuf_0__3398_/X vssd1 vssd1 vccd1 vccd1 _6914__425/A sky130_fd_sc_hd__clkbuf_4
X_5637_ _5727_/A _5815_/B vssd1 vssd1 vccd1 vccd1 _5653_/S sky130_fd_sc_hd__or2_2
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3435_ _7089_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3435_/X sky130_fd_sc_hd__clkbuf_16
X_5568_ _5568_/A vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8356_ _8356_/CLK _8356_/D vssd1 vssd1 vccd1 vccd1 _8356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4519_ _4347_/X _8181_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7307_ _7309_/A _7307_/B vssd1 vssd1 vccd1 vccd1 _8311_/D sky130_fd_sc_hd__nor2_1
X_8287_ _8315_/CLK _8287_/D vssd1 vssd1 vccd1 vccd1 _8287_/Q sky130_fd_sc_hd__dfxtp_2
X_8546__245 vssd1 vssd1 vccd1 vccd1 _8546__245/HI partID[13] sky130_fd_sc_hd__conb_1
X_5499_ _5499_/A vssd1 vssd1 vccd1 vccd1 _7993_/D sky130_fd_sc_hd__clkbuf_1
X_7238_ _7305_/A _7305_/B _7680_/A vssd1 vssd1 vccd1 vccd1 _7238_/Y sky130_fd_sc_hd__a21oi_1
X_7169_ _7176_/A vssd1 vssd1 vccd1 vccd1 _7193_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6599__306 _6600__307/A vssd1 vssd1 vccd1 vccd1 _7946_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4870_ _4425_/X _4610_/A _4869_/X _4841_/X vssd1 vssd1 vccd1 vccd1 _8134_/D sky130_fd_sc_hd__o211a_1
X_3821_ _8068_/Q _3920_/B vssd1 vssd1 vccd1 vccd1 _5018_/C sky130_fd_sc_hd__or2b_1
XFILLER_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6471_ _7852_/Q _7967_/Q _6714_/S vssd1 vssd1 vccd1 vccd1 _6472_/A sky130_fd_sc_hd__mux2_1
X_8210_ _8210_/CLK _8210_/D vssd1 vssd1 vccd1 vccd1 _8210_/Q sky130_fd_sc_hd__dfxtp_1
X_5422_ _3883_/X _8030_/Q _5422_/S vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5353_ _5565_/A vssd1 vssd1 vccd1 vccd1 _5353_/X sky130_fd_sc_hd__buf_2
Xclkbuf_0__3220_ _6498_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3220_/X sky130_fd_sc_hd__clkbuf_16
Xoutput202 _6030_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
X_8141_ _8141_/CLK _8141_/D vssd1 vssd1 vccd1 vccd1 _8141_/Q sky130_fd_sc_hd__dfxtp_1
X_4304_ _3943_/X _8263_/Q _4304_/S vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__mux2_1
X_5284_ _7784_/Q _8381_/Q _5294_/S vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__mux2_1
X_8072_ _8072_/CLK _8072_/D vssd1 vssd1 vccd1 vccd1 _8072_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_8 _4445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4235_ _8064_/Q vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__buf_2
XFILLER_114_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _4166_/A vssd1 vssd1 vccd1 vccd1 _8346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _8358_/Q _4018_/X _4099_/S vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7925_ _7925_/CLK _7925_/D vssd1 vssd1 vccd1 vccd1 _7925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7055__534 _7056__535/A vssd1 vssd1 vccd1 vccd1 _8215_/CLK sky130_fd_sc_hd__inv_2
X_7856_ _7856_/CLK _7856_/D vssd1 vssd1 vccd1 vccd1 _7856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6807_ _7457_/A _7457_/B _6395_/A vssd1 vssd1 vccd1 vccd1 _7499_/B sky130_fd_sc_hd__a21bo_1
X_7787_ _7787_/CLK _7787_/D vssd1 vssd1 vccd1 vccd1 _7787_/Q sky130_fd_sc_hd__dfxtp_1
X_4999_ _4999_/A _4999_/B _4999_/C vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__nand3_4
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6738_ _6751_/A vssd1 vssd1 vccd1 vccd1 _6789_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8408_ _8408_/CLK _8408_/D vssd1 vssd1 vccd1 vccd1 _8408_/Q sky130_fd_sc_hd__dfxtp_1
X_8339_ _8339_/CLK _8339_/D vssd1 vssd1 vccd1 vccd1 _8339_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3418_ _7007_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3418_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6587__298 _6588__299/A vssd1 vssd1 vccd1 vccd1 _7938_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8496_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4020_ _4020_/A vssd1 vssd1 vccd1 vccd1 _8390_/D sky130_fd_sc_hd__clkbuf_1
X_6904__416 _6906__418/A vssd1 vssd1 vccd1 vccd1 _8094_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5971_ _5971_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__and2_1
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7710_ _7478_/A _7707_/C _7709_/X _6421_/X vssd1 vssd1 vccd1 vccd1 _8494_/D sky130_fd_sc_hd__o211a_1
X_4922_ _4903_/B _4911_/C _4900_/X vssd1 vssd1 vccd1 vccd1 _4923_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _8192_/Q _4762_/X _4661_/A _4852_/X vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__o211a_1
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4784_ _7891_/Q _4767_/X _4782_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__o22a_1
X_7572_ _6819_/A _7572_/B _7572_/C vssd1 vssd1 vccd1 vccd1 _7572_/X sky130_fd_sc_hd__and3b_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3235_ clkbuf_0__3235_/X vssd1 vssd1 vccd1 vccd1 _6583__295/A sky130_fd_sc_hd__clkbuf_4
X_6454_ _6454_/A vssd1 vssd1 vccd1 vccd1 _7844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5405_ _5405_/A vssd1 vssd1 vccd1 vccd1 _8039_/D sky130_fd_sc_hd__clkbuf_1
X_6385_ _7689_/A _6390_/B _6387_/C vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__and3_1
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5336_ _5338_/A _5336_/B vssd1 vssd1 vccd1 vccd1 _5336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8124_ _8124_/CLK _8124_/D vssd1 vssd1 vccd1 vccd1 _8124_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8055_ _8055_/CLK _8055_/D vssd1 vssd1 vccd1 vccd1 _8055_/Q sky130_fd_sc_hd__dfxtp_1
X_5267_ _8366_/Q _5214_/A _5189_/X _8358_/Q _5074_/X vssd1 vssd1 vccd1 vccd1 _5267_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ _4218_/A vssd1 vssd1 vccd1 vccd1 _8327_/D sky130_fd_sc_hd__clkbuf_1
X_5198_ _8461_/Q _5292_/B _5108_/A _5197_/X vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__o211a_1
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _4149_/A vssd1 vssd1 vccd1 vccd1 _8352_/D sky130_fd_sc_hd__clkbuf_1
X_7908_ _7908_/CLK _7908_/D vssd1 vssd1 vccd1 vccd1 _7908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7839_ _8478_/CLK _7839_/D vssd1 vssd1 vccd1 vccd1 _7839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6257__194 _6258__195/A vssd1 vssd1 vccd1 vccd1 _7786_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6170_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5121_ _5062_/X _5120_/X _5278_/A vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__a21o_1
X_5052_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5052_/X sky130_fd_sc_hd__buf_2
XFILLER_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4003_ _8394_/Q _4002_/X _4011_/S vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5954_ _5954_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__and2_1
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__clkbuf_1
X_4905_ _6854_/A _4921_/A vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__nand2_2
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4836_ _8046_/Q _4765_/A _4659_/A _4835_/X vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7555_ _7504_/A _7577_/B _7508_/B vssd1 vssd1 vccd1 vccd1 _7556_/A sky130_fd_sc_hd__a21o_1
XFILLER_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4767_ _4767_/A vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4698_ _7782_/Q _7902_/Q _7910_/Q _7950_/Q _4650_/A _4640_/A vssd1 vssd1 vccd1 vccd1
+ _4698_/X sky130_fd_sc_hd__mux4_1
X_7486_ _7486_/A _7486_/B _7486_/C _7486_/D vssd1 vssd1 vccd1 vccd1 _7487_/D sky130_fd_sc_hd__or4_1
Xclkbuf_1_1_0__3218_ clkbuf_0__3218_/X vssd1 vssd1 vccd1 vccd1 _6494__223/A sky130_fd_sc_hd__clkbuf_4
X_6437_ _6437_/A vssd1 vssd1 vccd1 vccd1 _7836_/D sky130_fd_sc_hd__clkbuf_1
X_6368_ _7816_/Q _7654_/B _6365_/X _6367_/X vssd1 vssd1 vccd1 vccd1 _6369_/B sky130_fd_sc_hd__o22a_1
XFILLER_96_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8107_ _8107_/CLK _8107_/D vssd1 vssd1 vccd1 vccd1 _8107_/Q sky130_fd_sc_hd__dfxtp_1
X_5319_ _5319_/A _5322_/B vssd1 vssd1 vccd1 vccd1 _5319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6299_ _6355_/A vssd1 vssd1 vccd1 vccd1 _6299_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8038_ _8038_/CLK _8038_/D vssd1 vssd1 vccd1 vccd1 _8038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3434_ clkbuf_0__3434_/X vssd1 vssd1 vccd1 vccd1 _7088__60/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6699__344 _6700__345/A vssd1 vssd1 vccd1 vccd1 _8008_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7450__22 _7450__22/A vssd1 vssd1 vccd1 vccd1 _8408_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5670_ _5670_/A vssd1 vssd1 vccd1 vccd1 _7897_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4621_ _8126_/Q _4674_/B vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__xor2_2
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4552_ _4567_/S vssd1 vssd1 vccd1 vccd1 _4561_/S sky130_fd_sc_hd__buf_2
X_7340_ _8084_/Q _7324_/A _7326_/A _7339_/X _7331_/X vssd1 vssd1 vccd1 vccd1 _8321_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_116_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4483_ _4483_/A vssd1 vssd1 vccd1 vccd1 _8196_/D sky130_fd_sc_hd__clkbuf_1
X_7271_ _7286_/A vssd1 vssd1 vccd1 vccd1 _7272_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6222_ _6222_/A vssd1 vssd1 vccd1 vccd1 _7771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6172_/A vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__clkbuf_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5104_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__buf_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _7826_/Q input12/X _6107_/A vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5035_ _5054_/B _5046_/B vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__nor2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6544__263 _6544__263/A vssd1 vssd1 vccd1 vccd1 _7903_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5937_ _5937_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__or2_1
XFILLER_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5868_ _5868_/A vssd1 vssd1 vccd1 vccd1 _6006_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7607_ _7607_/A _7615_/B _7613_/C vssd1 vssd1 vccd1 vccd1 _7608_/A sky130_fd_sc_hd__and3_1
X_4819_ _4813_/X _4815_/X _4818_/X _4928_/B vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__a211o_1
X_5799_ _3812_/X _7791_/Q _5807_/S vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7538_ _8422_/Q _7530_/X _7527_/X _6763_/Y vssd1 vssd1 vccd1 vccd1 _7539_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7469_ _7468_/B _7468_/C _7468_/A vssd1 vssd1 vccd1 vccd1 _7472_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__buf_6
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3417_ clkbuf_0__3417_/X vssd1 vssd1 vccd1 vccd1 _7006__495/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3279_ clkbuf_0__3279_/X vssd1 vssd1 vccd1 vccd1 _6703__347/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7387__146 _7389__148/A vssd1 vssd1 vccd1 vccd1 _8357_/CLK sky130_fd_sc_hd__inv_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6487__217 _6488__218/A vssd1 vssd1 vccd1 vccd1 _7857_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3621_ clkbuf_0__3621_/X vssd1 vssd1 vccd1 vccd1 _7410__165/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771_ _8415_/Q vssd1 vssd1 vccd1 vccd1 _7473_/B sky130_fd_sc_hd__buf_2
X_3983_ _3934_/X _8400_/Q _3983_/S vssd1 vssd1 vccd1 vccd1 _3984_/A sky130_fd_sc_hd__mux2_1
X_5722_ _5722_/A vssd1 vssd1 vccd1 vccd1 _7874_/D sky130_fd_sc_hd__clkbuf_1
X_5653_ _5580_/X _7904_/Q _5653_/S vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__mux2_1
X_8441_ _8441_/CLK _8441_/D vssd1 vssd1 vccd1 vccd1 _8441_/Q sky130_fd_sc_hd__dfxtp_1
X_5584_ _5599_/S vssd1 vssd1 vccd1 vccd1 _5593_/S sky130_fd_sc_hd__clkbuf_4
X_8372_ _8372_/CLK _8372_/D vssd1 vssd1 vccd1 vccd1 _8372_/Q sky130_fd_sc_hd__dfxtp_1
X_4604_ _8143_/Q _4454_/X _4604_/S vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__mux2_1
X_4535_ _8174_/Q _4431_/X _4543_/S vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__mux2_1
X_7323_ _7323_/A vssd1 vssd1 vccd1 vccd1 _7324_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4466_ _4466_/A vssd1 vssd1 vccd1 vccd1 _8203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4397_ _4397_/A vssd1 vssd1 vccd1 vccd1 _8226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7185_ _7193_/B _7217_/B _7184_/A vssd1 vssd1 vccd1 vccd1 _7289_/B sky130_fd_sc_hd__a21o_1
X_6205_ _7975_/Q _6146_/X _6161_/A _6172_/A _7764_/Q vssd1 vssd1 vccd1 vccd1 _7764_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _7746_/Q _6082_/B vssd1 vssd1 vccd1 vccd1 _6067_/X sky130_fd_sc_hd__or2_1
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7019__505 _7019__505/A vssd1 vssd1 vccd1 vccd1 _8186_/CLK sky130_fd_sc_hd__inv_2
X_5018_ _5018_/A _5018_/B _5018_/C _5018_/D vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__and4_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601__308 _6603__310/A vssd1 vssd1 vccd1 vccd1 _7948_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4320_ _8256_/Q _4197_/X _4322_/S vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _5502_/B _5779_/B vssd1 vssd1 vccd1 vccd1 _4267_/S sky130_fd_sc_hd__nor2_2
X_4182_ _8448_/Q vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _7941_/CLK _7941_/D vssd1 vssd1 vccd1 vccd1 _7941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7872_ _7872_/CLK _7872_/D vssd1 vssd1 vccd1 vccd1 _7872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3966_ _8406_/Q _3889_/X _3968_/S vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6754_ _7459_/A _6754_/B vssd1 vssd1 vccd1 vccd1 _7497_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6992__483 _6994__485/A vssd1 vssd1 vccd1 vccd1 _8164_/CLK sky130_fd_sc_hd__inv_2
X_5705_ _7881_/Q _4993_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5636_ _5636_/A vssd1 vssd1 vccd1 vccd1 _7912_/D sky130_fd_sc_hd__clkbuf_1
X_3897_ _5321_/A _3897_/B vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__or2_2
X_8424_ _8425_/CLK _8424_/D vssd1 vssd1 vccd1 vccd1 _8424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3397_ clkbuf_0__3397_/X vssd1 vssd1 vccd1 vccd1 _6908__420/A sky130_fd_sc_hd__clkbuf_4
X_5567_ _5567_/A vssd1 vssd1 vccd1 vccd1 _7941_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3434_ _7083_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3434_/X sky130_fd_sc_hd__clkbuf_16
X_8355_ _8355_/CLK _8355_/D vssd1 vssd1 vccd1 vccd1 _8355_/Q sky130_fd_sc_hd__dfxtp_1
X_4518_ _4518_/A vssd1 vssd1 vccd1 vccd1 _8182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8286_ _8286_/CLK _8286_/D vssd1 vssd1 vccd1 vccd1 _8286_/Q sky130_fd_sc_hd__dfxtp_1
X_5498_ _5369_/X _7993_/Q _5500_/S vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__mux2_1
X_7306_ _8311_/Q _7295_/X _7272_/A _7305_/Y vssd1 vssd1 vccd1 vccd1 _7307_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4449_ _8209_/Q _4448_/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__mux2_1
X_7237_ _7680_/A _7305_/A _7305_/B vssd1 vssd1 vccd1 vccd1 _7237_/X sky130_fd_sc_hd__and3_1
XFILLER_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7168_ _8301_/Q vssd1 vssd1 vccd1 vccd1 _7211_/B sky130_fd_sc_hd__clkbuf_2
X_6251__189 _6252__190/A vssd1 vssd1 vccd1 vccd1 _7781_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6119_ _6119_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6119_/X sky130_fd_sc_hd__and2_1
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7641__47 _7643__49/A vssd1 vssd1 vccd1 vccd1 _8470_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3820_ _3920_/B vssd1 vssd1 vccd1 vccd1 _5328_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6470_ _6470_/A vssd1 vssd1 vccd1 vccd1 _7851_/D sky130_fd_sc_hd__clkbuf_1
X_5421_ _5421_/A vssd1 vssd1 vccd1 vccd1 _8031_/D sky130_fd_sc_hd__clkbuf_1
X_5352_ _8065_/Q vssd1 vssd1 vccd1 vccd1 _5565_/A sky130_fd_sc_hd__buf_2
Xoutput203 _6033_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
X_8140_ _8140_/CLK _8140_/D vssd1 vssd1 vccd1 vccd1 _8140_/Q sky130_fd_sc_hd__dfxtp_1
X_4303_ _4303_/A vssd1 vssd1 vccd1 vccd1 _8264_/D sky130_fd_sc_hd__clkbuf_1
X_8071_ _8071_/CLK _8071_/D vssd1 vssd1 vccd1 vccd1 _8071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5283_ _3940_/X _5022_/A _5281_/X _5282_/X vssd1 vssd1 vccd1 vccd1 _8080_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _8294_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_9 _6105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4165_ _8346_/Q _4002_/X _4169_/S vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4096_/A vssd1 vssd1 vccd1 vccd1 _8359_/D sky130_fd_sc_hd__clkbuf_1
X_7924_ _7924_/CLK _7924_/D vssd1 vssd1 vccd1 vccd1 _7924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7855_ _8498_/CLK _7855_/D vssd1 vssd1 vccd1 vccd1 _7855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6806_ _6395_/A _7457_/A _7457_/B vssd1 vssd1 vccd1 vccd1 _7499_/A sky130_fd_sc_hd__nand3b_1
X_4998_ _4998_/A vssd1 vssd1 vccd1 vccd1 _8097_/D sky130_fd_sc_hd__clkbuf_1
X_6693__339 _6694__340/A vssd1 vssd1 vccd1 vccd1 _8003_/CLK sky130_fd_sc_hd__inv_2
X_7786_ _7786_/CLK _7786_/D vssd1 vssd1 vccd1 vccd1 _7786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8513__212 vssd1 vssd1 vccd1 vccd1 _8513__212/HI caravel_irq[3] sky130_fd_sc_hd__conb_1
X_6737_ _8418_/Q _8417_/Q _8416_/Q _8415_/Q vssd1 vssd1 vccd1 vccd1 _6751_/A sky130_fd_sc_hd__and4_1
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3949_ _3949_/A _5328_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _5321_/B sky130_fd_sc_hd__and3_1
X_5619_ _5745_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5635_/S sky130_fd_sc_hd__nor2_2
X_8407_ _8407_/CLK _8407_/D vssd1 vssd1 vccd1 vccd1 _8407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8338_ _8338_/CLK _8338_/D vssd1 vssd1 vccd1 vccd1 _8338_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3417_ _7001_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3417_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8269_ _8269_/CLK _8269_/D vssd1 vssd1 vccd1 vccd1 _8269_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3279_ _6701_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3279_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7084__56 _7085__57/A vssd1 vssd1 vccd1 vccd1 _8237_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6999__489 _6999__489/A vssd1 vssd1 vccd1 vccd1 _8170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6269__203 _6271__205/A vssd1 vssd1 vccd1 vccd1 _7795_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5970_ _5970_/A vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4921_ _4921_/A _4921_/B vssd1 vssd1 vccd1 vccd1 _8128_/D sky130_fd_sc_hd__nor2_1
X_4852_ _7889_/Q _4767_/A _4851_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4783_ _4793_/A vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__clkbuf_2
X_7571_ _8432_/Q _7563_/A _8433_/Q vssd1 vssd1 vccd1 vccd1 _7572_/B sky130_fd_sc_hd__a21o_1
X_6522_ _6522_/A vssd1 vssd1 vccd1 vccd1 _6522_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3234_ clkbuf_0__3234_/X vssd1 vssd1 vccd1 vccd1 _6574__287/A sky130_fd_sc_hd__clkbuf_4
X_7408__163 _7409__164/A vssd1 vssd1 vccd1 vccd1 _8374_/CLK sky130_fd_sc_hd__inv_2
X_6453_ _7844_/Q _7959_/Q _6455_/S vssd1 vssd1 vccd1 vccd1 _6454_/A sky130_fd_sc_hd__mux2_1
X_5404_ _5361_/X _8039_/Q _5404_/S vssd1 vssd1 vccd1 vccd1 _5405_/A sky130_fd_sc_hd__mux2_1
X_6384_ _8488_/Q vssd1 vssd1 vccd1 vccd1 _7689_/A sky130_fd_sc_hd__buf_2
X_8123_ _8123_/CLK _8123_/D vssd1 vssd1 vccd1 vccd1 _8123_/Q sky130_fd_sc_hd__dfxtp_4
X_5335_ _5054_/A _5331_/X _5334_/Y _5249_/X vssd1 vssd1 vccd1 vccd1 _8071_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8054_ _8054_/CLK _8054_/D vssd1 vssd1 vccd1 vccd1 _8054_/Q sky130_fd_sc_hd__dfxtp_1
X_5266_ _8334_/Q _8342_/Q _5269_/S vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _8327_/Q _4150_/X _4221_/S vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__mux2_1
X_5197_ _8453_/Q _5046_/B _5196_/X _5207_/A vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6508__234 _6508__234/A vssd1 vssd1 vccd1 vccd1 _7874_/CLK sky130_fd_sc_hd__inv_2
X_4148_ _8352_/Q _4147_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4079_ _3940_/X _8366_/Q _4081_/S vssd1 vssd1 vccd1 vccd1 _4080_/A sky130_fd_sc_hd__mux2_1
X_7907_ _7907_/CLK _7907_/D vssd1 vssd1 vccd1 vccd1 _7907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7838_ _8497_/CLK _7838_/D vssd1 vssd1 vccd1 vccd1 _7838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7769_ _8308_/CLK _7769_/D vssd1 vssd1 vccd1 vccd1 _7769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6717__353 _6718__354/A vssd1 vssd1 vccd1 vccd1 _8020_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6910__421 _6911__422/A vssd1 vssd1 vccd1 vccd1 _8099_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _8394_/Q _8386_/Q _7789_/Q _8402_/Q _5063_/X _5064_/X vssd1 vssd1 vccd1 vccd1
+ _5120_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5051_ _5164_/A vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__buf_2
XFILLER_97_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4350_/A vssd1 vssd1 vccd1 vccd1 _4002_/X sky130_fd_sc_hd__buf_2
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5953_ _5953_/A vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _7609_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__or2_1
X_4904_ _4904_/A _4923_/A vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__and2_1
X_4835_ _8107_/Q _4767_/A _4834_/X _4793_/A vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _4766_/A vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__clkbuf_2
X_7554_ _7554_/A _7554_/B vssd1 vssd1 vccd1 vccd1 _8429_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4697_ _7926_/Q _7806_/Q _7731_/Q _7918_/Q _4670_/X _4638_/X vssd1 vssd1 vccd1 vccd1
+ _4697_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1_0__3217_ clkbuf_0__3217_/X vssd1 vssd1 vccd1 vccd1 _6490__220/A sky130_fd_sc_hd__clkbuf_4
X_7485_ _7483_/Y _7484_/X _6395_/A _6746_/A vssd1 vssd1 vccd1 vccd1 _7486_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6436_ _7836_/Q _5960_/A _6444_/S vssd1 vssd1 vccd1 vccd1 _6437_/A sky130_fd_sc_hd__mux2_1
X_6367_ _7698_/A _8017_/Q _6292_/B _6352_/A _6343_/A vssd1 vssd1 vccd1 vccd1 _6367_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8106_ _8106_/CLK _8106_/D vssd1 vssd1 vccd1 vccd1 _8106_/Q sky130_fd_sc_hd__dfxtp_1
X_5318_ _3897_/B _5322_/B _5317_/X _5282_/X vssd1 vssd1 vccd1 vccd1 _8077_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6298_ _7654_/A _6312_/B vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__or2_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8037_ _8037_/CLK _8037_/D vssd1 vssd1 vccd1 vccd1 _8037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8497_/CLK sky130_fd_sc_hd__clkbuf_16
X_5249_ _6892_/A vssd1 vssd1 vccd1 vccd1 _5249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3433_ clkbuf_0__3433_/X vssd1 vssd1 vccd1 vccd1 _7079__52/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7068__545 _7068__545/A vssd1 vssd1 vccd1 vccd1 _8226_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7012__500 _7012__500/A vssd1 vssd1 vccd1 vccd1 _8181_/CLK sky130_fd_sc_hd__inv_2
X_4620_ _4653_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4674_/B sky130_fd_sc_hd__and2_2
XFILLER_116_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4551_ _5815_/A _4936_/A vssd1 vssd1 vccd1 vccd1 _4567_/S sky130_fd_sc_hd__or2_2
X_4482_ _8196_/Q _4232_/X _4486_/S vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7270_ _7270_/A _7270_/B vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__or2_1
XFILLER_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6221_ _7707_/A _7771_/Q _6223_/S vssd1 vssd1 vccd1 vccd1 _6222_/A sky130_fd_sc_hd__mux2_1
X_6152_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__buf_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5103_ _5099_/X _5100_/X _5102_/X vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__a21o_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6072_/X _6081_/X _6082_/X _6075_/X vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__o211a_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5034_ _5164_/A _5196_/S _8070_/Q vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__a21oi_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5936_ _5936_/A vssd1 vssd1 vccd1 vccd1 _5936_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5867_ _5867_/A vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7606_ _7703_/A vssd1 vssd1 vccd1 vccd1 _7615_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4818_ _7778_/Q _4765_/X _4816_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _4818_/X sky130_fd_sc_hd__o211a_1
X_5798_ _5813_/S vssd1 vssd1 vccd1 vccd1 _5807_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4749_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__clkbuf_2
X_7537_ _7546_/A _7537_/B vssd1 vssd1 vccd1 vccd1 _8421_/D sky130_fd_sc_hd__nor2_1
X_7468_ _7468_/A _7468_/B _7468_/C vssd1 vssd1 vccd1 vccd1 _7472_/A sky130_fd_sc_hd__and3_1
X_6419_ _6419_/A _7503_/A _7649_/B _7604_/B vssd1 vssd1 vccd1 vccd1 _6419_/X sky130_fd_sc_hd__or4b_2
X_7399_ _7417_/A vssd1 vssd1 vccd1 vccd1 _7399_/X sky130_fd_sc_hd__buf_1
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _6606_/A sky130_fd_sc_hd__buf_6
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3416_ clkbuf_0__3416_/X vssd1 vssd1 vccd1 vccd1 _6999__489/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3278_ clkbuf_0__3278_/X vssd1 vssd1 vccd1 vccd1 _6700__345/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7105__74 _7106__75/A vssd1 vssd1 vccd1 vccd1 _8255_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3620_ clkbuf_0__3620_/X vssd1 vssd1 vccd1 vccd1 _7401__157/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3982_ _3982_/A vssd1 vssd1 vccd1 vccd1 _8401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6770_ _8416_/Q vssd1 vssd1 vccd1 vccd1 _6782_/C sky130_fd_sc_hd__clkbuf_2
X_5721_ _4150_/X _7874_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5652_ _5652_/A vssd1 vssd1 vccd1 vccd1 _7905_/D sky130_fd_sc_hd__clkbuf_1
X_8440_ _8441_/CLK _8440_/D vssd1 vssd1 vccd1 vccd1 _8440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5583_ _5673_/B _5709_/B vssd1 vssd1 vccd1 vccd1 _5599_/S sky130_fd_sc_hd__or2_4
X_4603_ _4603_/A vssd1 vssd1 vccd1 vccd1 _8144_/D sky130_fd_sc_hd__clkbuf_1
X_8371_ _8371_/CLK _8371_/D vssd1 vssd1 vccd1 vccd1 _8371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4534_ _4549_/S vssd1 vssd1 vccd1 vccd1 _4543_/S sky130_fd_sc_hd__buf_2
X_7322_ _8315_/Q _7331_/A _7318_/X _7321_/Y vssd1 vssd1 vccd1 vccd1 _8315_/D sky130_fd_sc_hd__a31o_1
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _4353_/X _8203_/Q _4467_/S vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__mux2_1
X_4396_ _4356_/X _8226_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__mux2_1
X_7184_ _7184_/A _7217_/A _7217_/B vssd1 vssd1 vccd1 vccd1 _7289_/A sky130_fd_sc_hd__nand3_1
X_6204_ _7974_/Q _6146_/X _6161_/A _6172_/A _7763_/Q vssd1 vssd1 vccd1 vccd1 _7763_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6066_ _6085_/A vssd1 vssd1 vccd1 vccd1 _6082_/B sky130_fd_sc_hd__clkbuf_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _8089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3063_ clkbuf_0__3063_/X vssd1 vssd1 vccd1 vccd1 _6283__215/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5919_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5928_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6493__222 _6494__223/A vssd1 vssd1 vccd1 vccd1 _7862_/CLK sky130_fd_sc_hd__inv_2
X_8530__229 vssd1 vssd1 vccd1 vccd1 _8530__229/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
X_6870__393 _6872__395/A vssd1 vssd1 vccd1 vccd1 _8069_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4250_/A _4287_/B _5321_/A vssd1 vssd1 vccd1 vccd1 _5779_/B sky130_fd_sc_hd__nand3_4
X_7402__158 _7404__160/A vssd1 vssd1 vccd1 vccd1 _8369_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4181_ _4181_/A vssd1 vssd1 vccd1 vccd1 _8340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7940_ _7940_/CLK _7940_/D vssd1 vssd1 vccd1 vccd1 _7940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7871_ _7871_/CLK _7871_/D vssd1 vssd1 vccd1 vccd1 _7871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6502__229 _6503__230/A vssd1 vssd1 vccd1 vccd1 _7869_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3965_ _3965_/A vssd1 vssd1 vccd1 vccd1 _8407_/D sky130_fd_sc_hd__clkbuf_1
X_6753_ _7484_/B _7484_/C vssd1 vssd1 vccd1 vccd1 _6754_/B sky130_fd_sc_hd__nand2_1
X_5704_ _5704_/A vssd1 vssd1 vccd1 vccd1 _7882_/D sky130_fd_sc_hd__clkbuf_1
X_3896_ _4287_/A _8076_/Q vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__nand2_1
X_5635_ _7912_/Q _4996_/X _5635_/S vssd1 vssd1 vccd1 vccd1 _5636_/A sky130_fd_sc_hd__mux2_1
X_8423_ _8425_/CLK _8423_/D vssd1 vssd1 vccd1 vccd1 _8423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3396_ clkbuf_0__3396_/X vssd1 vssd1 vccd1 vccd1 _6902__415/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3433_ _7077_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3433_/X sky130_fd_sc_hd__clkbuf_16
X_5566_ _5565_/X _7941_/Q _5572_/S vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__mux2_1
X_8354_ _8354_/CLK _8354_/D vssd1 vssd1 vccd1 vccd1 _8354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4517_ _4342_/X _8182_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__mux2_1
X_8285_ _8285_/CLK _8285_/D vssd1 vssd1 vccd1 vccd1 _8285_/Q sky130_fd_sc_hd__dfxtp_1
X_5497_ _5497_/A vssd1 vssd1 vccd1 vccd1 _7994_/D sky130_fd_sc_hd__clkbuf_1
X_7305_ _7305_/A _7305_/B vssd1 vssd1 vccd1 vccd1 _7305_/Y sky130_fd_sc_hd__nand2_1
X_7025__510 _7025__510/A vssd1 vssd1 vccd1 vccd1 _8191_/CLK sky130_fd_sc_hd__inv_2
X_4448_ _8444_/Q vssd1 vssd1 vccd1 vccd1 _4448_/X sky130_fd_sc_hd__buf_4
X_7236_ _7234_/X _7236_/B _7236_/C _7236_/D vssd1 vssd1 vccd1 vccd1 _7246_/C sky130_fd_sc_hd__and4b_1
X_4379_ _4379_/A vssd1 vssd1 vccd1 vccd1 _8234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7167_ _8302_/Q vssd1 vssd1 vccd1 vccd1 _7211_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _7761_/Q _6111_/X _6112_/X _6117_/X _6109_/X vssd1 vssd1 vccd1 vccd1 _6118_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _6034_/X _6046_/X _6048_/X _6037_/X vssd1 vssd1 vccd1 vccd1 _6049_/X sky130_fd_sc_hd__o211a_1
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6557__274 _6558__275/A vssd1 vssd1 vccd1 vccd1 _7914_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5420_ _3880_/X _8031_/Q _5422_/S vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__mux2_1
X_5351_ _5351_/A vssd1 vssd1 vccd1 vccd1 _8058_/D sky130_fd_sc_hd__clkbuf_1
Xoutput204 _6038_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4302_ _3940_/X _8264_/Q _4304_/S vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__mux2_1
X_8070_ _8070_/CLK _8070_/D vssd1 vssd1 vccd1 vccd1 _8070_/Q sky130_fd_sc_hd__dfxtp_2
X_5282_ _7598_/A vssd1 vssd1 vccd1 vccd1 _5282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _8294_/Q _4232_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4164_ _4164_/A vssd1 vssd1 vccd1 vccd1 _8347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _8359_/Q _4014_/X _4099_/S vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7923_ _7923_/CLK _7923_/D vssd1 vssd1 vccd1 vccd1 _7923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7854_ _8017_/CLK _7854_/D vssd1 vssd1 vccd1 vccd1 _7854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7785_ _7785_/CLK _7785_/D vssd1 vssd1 vccd1 vccd1 _7785_/Q sky130_fd_sc_hd__dfxtp_1
X_6805_ _8428_/Q _6745_/B _8429_/Q vssd1 vssd1 vccd1 vccd1 _7457_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6877__399 _6878__400/A vssd1 vssd1 vccd1 vccd1 _8075_/CLK sky130_fd_sc_hd__inv_2
X_4997_ _8097_/Q _4996_/X _4997_/S vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__mux2_1
X_6736_ _8426_/Q _8425_/Q _8424_/Q _8423_/Q vssd1 vssd1 vccd1 vccd1 _6808_/A sky130_fd_sc_hd__and4_1
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ _3948_/A vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__clkbuf_2
X_3879_ _3879_/A vssd1 vssd1 vccd1 vccd1 _8471_/D sky130_fd_sc_hd__clkbuf_1
X_5618_ _5618_/A vssd1 vssd1 vccd1 vccd1 _7920_/D sky130_fd_sc_hd__clkbuf_1
X_6598_ _6598_/A vssd1 vssd1 vccd1 vccd1 _6598_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3379_ clkbuf_0__3379_/X vssd1 vssd1 vccd1 vccd1 _6851__391/A sky130_fd_sc_hd__clkbuf_4
X_8406_ _8406_/CLK _8406_/D vssd1 vssd1 vccd1 vccd1 _8406_/Q sky130_fd_sc_hd__dfxtp_1
X_5549_ _7947_/Q _4987_/X _5549_/S vssd1 vssd1 vccd1 vccd1 _5550_/A sky130_fd_sc_hd__mux2_1
X_8337_ _8337_/CLK _8337_/D vssd1 vssd1 vccd1 vccd1 _8337_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3416_ _6995_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3416_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8268_ _8268_/CLK _8268_/D vssd1 vssd1 vccd1 vccd1 _8268_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3278_ _6695_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3278_/X sky130_fd_sc_hd__clkbuf_16
X_8199_ _8199_/CLK _8199_/D vssd1 vssd1 vccd1 vccd1 _8199_/Q sky130_fd_sc_hd__dfxtp_1
X_7219_ _7195_/A _7195_/B _7459_/A vssd1 vssd1 vccd1 vccd1 _7219_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936__441 _6937__442/A vssd1 vssd1 vccd1 vccd1 _8119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_opt_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8309_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4920_ _4904_/A _4923_/A _4900_/X vssd1 vssd1 vccd1 vccd1 _4921_/B sky130_fd_sc_hd__o21ai_1
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4851_ _4801_/A _7993_/Q _7929_/Q _4787_/A vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__a22o_1
X_8536__235 vssd1 vssd1 vccd1 vccd1 _8536__235/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _4801_/A _7995_/Q _7931_/Q _4787_/A vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__a22o_1
X_7570_ _8432_/Q _7562_/Y _7569_/X _7514_/X vssd1 vssd1 vccd1 vccd1 _8432_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3233_ clkbuf_0__3233_/X vssd1 vssd1 vccd1 vccd1 _6571__285/A sky130_fd_sc_hd__clkbuf_4
X_6452_ _6452_/A vssd1 vssd1 vccd1 vccd1 _7843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _5403_/A vssd1 vssd1 vccd1 vccd1 _8040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6383_ _6401_/A vssd1 vssd1 vccd1 vccd1 _6383_/X sky130_fd_sc_hd__clkbuf_2
X_8122_ _8122_/CLK _8122_/D vssd1 vssd1 vccd1 vccd1 _8122_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5334_ _5338_/A _5334_/B vssd1 vssd1 vccd1 vccd1 _5334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8053_ _8053_/CLK _8053_/D vssd1 vssd1 vccd1 vccd1 _8053_/Q sky130_fd_sc_hd__dfxtp_1
X_5265_ _5083_/X _5254_/Y _5257_/Y _5264_/X vssd1 vssd1 vccd1 vccd1 _5280_/A sky130_fd_sc_hd__a31o_1
Xclkbuf_0__3063_ _6278_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3063_/X sky130_fd_sc_hd__clkbuf_16
X_5196_ _7987_/Q _8022_/Q _5196_/S vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__mux2_1
X_4216_ _4216_/A vssd1 vssd1 vccd1 vccd1 _8328_/D sky130_fd_sc_hd__clkbuf_1
X_4147_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _4147_/X sky130_fd_sc_hd__buf_2
XFILLER_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4078_ _4078_/A vssd1 vssd1 vccd1 vccd1 _8367_/D sky130_fd_sc_hd__clkbuf_1
X_7906_ _7906_/CLK _7906_/D vssd1 vssd1 vccd1 vccd1 _7906_/Q sky130_fd_sc_hd__dfxtp_1
X_7837_ _8497_/CLK _7837_/D vssd1 vssd1 vccd1 vccd1 _7837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7768_ _8308_/CLK _7768_/D vssd1 vssd1 vccd1 vccd1 _7768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7699_ _7699_/A _7699_/B vssd1 vssd1 vccd1 vccd1 _7699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6669__320 _6669__320/A vssd1 vssd1 vccd1 vccd1 _7984_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5190_/S vssd1 vssd1 vccd1 vccd1 _5294_/S sky130_fd_sc_hd__buf_4
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4001_ _8447_/Q vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7254__109 _7255__110/A vssd1 vssd1 vccd1 vccd1 _8292_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5952_ _5952_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__and2_1
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _4903_/A _4903_/B _7645_/B vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__and3_1
X_5883_ _5883_/A vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4834_ _4780_/A _8038_/Q _7866_/Q _4781_/A vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4765_ _4765_/A vssd1 vssd1 vccd1 vccd1 _4765_/X sky130_fd_sc_hd__buf_2
X_7553_ _8429_/Q _7510_/B _7544_/X _7458_/B vssd1 vssd1 vccd1 vccd1 _7554_/B sky130_fd_sc_hd__o2bb2a_1
X_6504_ _6510_/A vssd1 vssd1 vccd1 vccd1 _6504_/X sky130_fd_sc_hd__buf_1
X_4696_ _4692_/X _4693_/X _4696_/S vssd1 vssd1 vccd1 vccd1 _4696_/X sky130_fd_sc_hd__mux2_1
X_7484_ _8486_/Q _7484_/B _7484_/C vssd1 vssd1 vccd1 vccd1 _7484_/X sky130_fd_sc_hd__and3_1
XFILLER_106_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6435_ _6468_/A vssd1 vssd1 vccd1 vccd1 _6444_/S sky130_fd_sc_hd__clkbuf_2
X_6366_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _7698_/A sky130_fd_sc_hd__clkbuf_4
X_8105_ _8105_/CLK _8105_/D vssd1 vssd1 vccd1 vccd1 _8105_/Q sky130_fd_sc_hd__dfxtp_1
X_5317_ _4287_/B _5316_/A _5328_/B _4250_/A vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__a31o_1
X_6137__178 _6138__179/A vssd1 vssd1 vccd1 vccd1 _7727_/CLK sky130_fd_sc_hd__inv_2
X_8036_ _8036_/CLK _8036_/D vssd1 vssd1 vccd1 vccd1 _8036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6297_ _7659_/B _6297_/B vssd1 vssd1 vccd1 vccd1 _6312_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5248_ _8081_/Q _5024_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5248_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_0_0__3432_ clkbuf_0__3432_/X vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__clkbuf_4
X_5179_ _5215_/A vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__buf_2
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7117__83 _7118__84/A vssd1 vssd1 vccd1 vccd1 _8264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7435__10 _7434__9/A vssd1 vssd1 vccd1 vccd1 _8396_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7357__122 _7360__125/A vssd1 vssd1 vccd1 vccd1 _8333_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4550_ _4550_/A vssd1 vssd1 vccd1 vccd1 _8167_/D sky130_fd_sc_hd__clkbuf_1
X_4481_ _4481_/A vssd1 vssd1 vccd1 vccd1 _8197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _6220_/A vssd1 vssd1 vccd1 vccd1 _7770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6151_ _6157_/A _6231_/B vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__or2_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5102_ _5062_/X _5101_/X _5056_/X vssd1 vssd1 vccd1 vccd1 _5102_/X sky130_fd_sc_hd__a21o_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _7750_/Q _6082_/B vssd1 vssd1 vccd1 vccd1 _6082_/X sky130_fd_sc_hd__or2_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5033_ _8068_/Q vssd1 vssd1 vccd1 vccd1 _5196_/S sky130_fd_sc_hd__buf_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5935_ _5935_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__or2_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5866_ _6606_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__and2_1
XFILLER_34_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4817_ _4796_/A _7906_/Q _7898_/Q _4753_/A _4757_/A vssd1 vssd1 vccd1 vccd1 _4817_/X
+ sky130_fd_sc_hd__a221o_1
X_7605_ _7605_/A vssd1 vssd1 vccd1 vccd1 _8444_/D sky130_fd_sc_hd__clkbuf_1
X_5797_ _5797_/A _5797_/B vssd1 vssd1 vccd1 vccd1 _5813_/S sky130_fd_sc_hd__or2_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _4769_/A vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7536_ _7468_/B _7468_/C _7516_/X _7522_/X _6789_/A vssd1 vssd1 vccd1 vccd1 _7537_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7467_ _6802_/A _6757_/A _6757_/B _7465_/X _7466_/Y vssd1 vssd1 vccd1 vccd1 _7486_/A
+ sky130_fd_sc_hd__a311o_1
X_4679_ _4612_/X _8140_/Q _4924_/A _4676_/X _4678_/X vssd1 vssd1 vccd1 vccd1 _4679_/X
+ sky130_fd_sc_hd__a221o_1
X_6418_ _7654_/B _6418_/B vssd1 vssd1 vccd1 vccd1 _7604_/B sky130_fd_sc_hd__nor2_2
X_6551__269 _6552__270/A vssd1 vssd1 vccd1 vccd1 _7909_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6349_ _6289_/A _6346_/X _6348_/X _6369_/A vssd1 vssd1 vccd1 vccd1 _6349_/X sky130_fd_sc_hd__a31o_1
Xinput104 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _6624_/A sky130_fd_sc_hd__buf_6
XFILLER_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8019_ _8019_/CLK _8019_/D vssd1 vssd1 vccd1 vccd1 _8019_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3415_ clkbuf_0__3415_/X vssd1 vssd1 vccd1 vccd1 _6991__482/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__3430_ clkbuf_0__3430_/X vssd1 vssd1 vccd1 vccd1 _7073__549/A sky130_fd_sc_hd__clkbuf_16
XFILLER_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7074__550 _7074__550/A vssd1 vssd1 vccd1 vccd1 _8231_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3277_ clkbuf_0__3277_/X vssd1 vssd1 vccd1 vccd1 _6692__338/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3628_ clkbuf_0__3628_/X vssd1 vssd1 vccd1 vccd1 _7445__18/A sky130_fd_sc_hd__clkbuf_16
XFILLER_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3981_ _3931_/X _8401_/Q _3983_/S vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5720_ _5720_/A vssd1 vssd1 vccd1 vccd1 _7875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5651_ _5577_/X _7905_/Q _5653_/S vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5582_ _5582_/A vssd1 vssd1 vccd1 vccd1 _7936_/D sky130_fd_sc_hd__clkbuf_1
X_4602_ _8144_/Q _4451_/X _4604_/S vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__mux2_1
X_8370_ _8370_/CLK _8370_/D vssd1 vssd1 vccd1 vccd1 _8370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4533_ _5779_/A _4588_/A vssd1 vssd1 vccd1 vccd1 _4549_/S sky130_fd_sc_hd__nor2_2
X_7321_ _7321_/A _7321_/B _7321_/C vssd1 vssd1 vccd1 vccd1 _7321_/Y sky130_fd_sc_hd__nor3_1
X_4464_ _4464_/A vssd1 vssd1 vccd1 vccd1 _8204_/D sky130_fd_sc_hd__clkbuf_1
X_6203_ _7973_/Q _6197_/X _6161_/A _6198_/X _7762_/Q vssd1 vssd1 vccd1 vccd1 _7762_/D
+ sky130_fd_sc_hd__o32a_1
X_6882__402 _6882__402/A vssd1 vssd1 vccd1 vccd1 _8078_/CLK sky130_fd_sc_hd__inv_2
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _8227_/D sky130_fd_sc_hd__clkbuf_1
X_7183_ _7183_/A _7183_/B _7236_/B vssd1 vssd1 vccd1 vccd1 _7222_/C sky130_fd_sc_hd__and3_1
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6134_ _6259_/A vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__buf_1
XFILLER_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7111__78 _7113__80/A vssd1 vssd1 vccd1 vccd1 _8259_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6065_ _7821_/Q input7/X _6077_/S vssd1 vssd1 vccd1 vccd1 _6065_/X sky130_fd_sc_hd__mux2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _4428_/X _8089_/Q _5016_/S vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5918_ _5918_/A vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3062_ clkbuf_0__3062_/X vssd1 vssd1 vccd1 vccd1 _6275__208/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5849_ _4156_/X _7725_/Q _5849_/S vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__mux2_1
X_6930__436 _6932__438/A vssd1 vssd1 vccd1 vccd1 _8114_/CLK sky130_fd_sc_hd__inv_2
X_7519_ _7597_/A _6242_/X _6482_/A vssd1 vssd1 vccd1 vccd1 _7535_/A sky130_fd_sc_hd__a21o_1
X_8499_ _8499_/CLK _8499_/D vssd1 vssd1 vccd1 vccd1 _8499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4180_ _8340_/Q _4177_/X _4192_/S vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7870_ _7870_/CLK _7870_/D vssd1 vssd1 vccd1 vccd1 _7870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6821_ _6821_/A vssd1 vssd1 vccd1 vccd1 _8035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _8407_/Q _3886_/X _3968_/S vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__mux2_1
X_6752_ _6808_/A _6786_/B _6749_/A _8427_/Q vssd1 vssd1 vccd1 vccd1 _7484_/C sky130_fd_sc_hd__a31o_1
X_6683_ _6683_/A vssd1 vssd1 vccd1 vccd1 _6683_/X sky130_fd_sc_hd__buf_1
X_5703_ _7882_/Q _4990_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__mux2_1
X_3895_ _3972_/B vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__buf_2
X_5634_ _5634_/A vssd1 vssd1 vccd1 vccd1 _7913_/D sky130_fd_sc_hd__clkbuf_1
X_8422_ _8425_/CLK _8422_/D vssd1 vssd1 vccd1 vccd1 _8422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3432_ _7076_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3432_/X sky130_fd_sc_hd__clkbuf_16
X_8353_ _8353_/CLK _8353_/D vssd1 vssd1 vccd1 vccd1 _8353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5565_ _5565_/A vssd1 vssd1 vccd1 vccd1 _5565_/X sky130_fd_sc_hd__clkbuf_2
X_7304_ _7309_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _8310_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4516_ _4531_/S vssd1 vssd1 vccd1 vccd1 _4525_/S sky130_fd_sc_hd__buf_2
X_8284_ _8284_/CLK _8284_/D vssd1 vssd1 vccd1 vccd1 _8284_/Q sky130_fd_sc_hd__dfxtp_1
X_5496_ _5365_/X _7994_/Q _5500_/S vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__mux2_1
X_4447_ _4447_/A vssd1 vssd1 vccd1 vccd1 _8210_/D sky130_fd_sc_hd__clkbuf_1
X_7235_ _8487_/Q _7195_/Y _7186_/X _7187_/Y _7216_/X vssd1 vssd1 vccd1 vccd1 _7236_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7166_ _7217_/A _7217_/B vssd1 vssd1 vccd1 vccd1 _7232_/B sky130_fd_sc_hd__nand2_1
X_4378_ _4356_/X _8234_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__mux2_1
X_7096__66 _7098__68/A vssd1 vssd1 vccd1 vccd1 _8247_/CLK sky130_fd_sc_hd__inv_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6117_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6117_/X sky130_fd_sc_hd__and2_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6663__315 _6663__315/A vssd1 vssd1 vccd1 vccd1 _7979_/CLK sky130_fd_sc_hd__inv_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6048_ _7741_/Q _6063_/B vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__or2_1
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _7999_/CLK _7999_/D vssd1 vssd1 vccd1 vccd1 _7999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6889__408 _6891__410/A vssd1 vssd1 vccd1 vccd1 _8084_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6969__465 _6969__465/A vssd1 vssd1 vccd1 vccd1 _8146_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7626__35 _7626__35/A vssd1 vssd1 vccd1 vccd1 _8458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6564__279 _6565__280/A vssd1 vssd1 vccd1 vccd1 _7919_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5350_ _5349_/X _8058_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__mux2_1
X_7434__9 _7434__9/A vssd1 vssd1 vccd1 vccd1 _8395_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput205 _6041_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4301_ _4301_/A vssd1 vssd1 vccd1 vccd1 _8265_/D sky130_fd_sc_hd__clkbuf_1
X_5281_ _8080_/Q _5025_/A _5246_/A _5280_/Y _5088_/A vssd1 vssd1 vccd1 vccd1 _5281_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7020_ _7026_/A vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__buf_1
X_4232_ _8065_/Q vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__buf_2
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4163_ _8347_/Q _3998_/X _4169_/S vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__mux2_1
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _8360_/D sky130_fd_sc_hd__clkbuf_1
X_7922_ _7922_/CLK _7922_/D vssd1 vssd1 vccd1 vccd1 _7922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7853_ _8017_/CLK _7853_/D vssd1 vssd1 vccd1 vccd1 _7853_/Q sky130_fd_sc_hd__dfxtp_1
X_7784_ _7784_/CLK _7784_/D vssd1 vssd1 vccd1 vccd1 _7784_/Q sky130_fd_sc_hd__dfxtp_1
X_4996_ _8060_/Q vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6804_ _7683_/A _7498_/B _7497_/A _6794_/X _6803_/X vssd1 vssd1 vccd1 vccd1 _6816_/B
+ sky130_fd_sc_hd__o2111a_1
X_3947_ _4250_/A _5319_/A _3972_/B vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__or3b_4
XFILLER_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6735_ _7597_/A _6242_/X _6157_/A vssd1 vssd1 vccd1 vccd1 _7575_/A sky130_fd_sc_hd__a21oi_4
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3878_ _8471_/Q _3877_/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5617_ _5580_/X _7920_/Q _5617_/S vssd1 vssd1 vccd1 vccd1 _5618_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3378_ clkbuf_0__3378_/X vssd1 vssd1 vccd1 vccd1 _6849__390/A sky130_fd_sc_hd__clkbuf_4
X_8405_ _8405_/CLK _8405_/D vssd1 vssd1 vccd1 vccd1 _8405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5548_ _5548_/A vssd1 vssd1 vccd1 vccd1 _7948_/D sky130_fd_sc_hd__clkbuf_1
X_8336_ _8336_/CLK _8336_/D vssd1 vssd1 vccd1 vccd1 _8336_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3415_ _6989_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3415_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_3_0_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8267_ _8267_/CLK _8267_/D vssd1 vssd1 vccd1 vccd1 _8267_/Q sky130_fd_sc_hd__dfxtp_1
X_5479_ _5479_/A vssd1 vssd1 vccd1 vccd1 _8002_/D sky130_fd_sc_hd__clkbuf_1
X_7218_ _7292_/A _7292_/B _6802_/A vssd1 vssd1 vccd1 vccd1 _7218_/X sky130_fd_sc_hd__a21o_1
X_8198_ _8198_/CLK _8198_/D vssd1 vssd1 vccd1 vccd1 _8198_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3277_ _6689_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3277_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7149_ _8304_/Q _8303_/Q _8302_/Q _8301_/Q vssd1 vssd1 vccd1 vccd1 _7173_/A sky130_fd_sc_hd__and4_1
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7351__117 _7351__117/A vssd1 vssd1 vccd1 vccd1 _8328_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943__446 _6944__447/A vssd1 vssd1 vccd1 vccd1 _8125_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _8290_/Q _4778_/X _8098_/Q _4762_/X _4696_/S vssd1 vssd1 vccd1 vccd1 _4850_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4781_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3232_ clkbuf_0__3232_/X vssd1 vssd1 vccd1 vccd1 _6563__278/A sky130_fd_sc_hd__clkbuf_4
X_6276__209 _6277__210/A vssd1 vssd1 vccd1 vccd1 _7801_/CLK sky130_fd_sc_hd__inv_2
X_6451_ _7843_/Q _5976_/A _6455_/S vssd1 vssd1 vccd1 vccd1 _6452_/A sky130_fd_sc_hd__mux2_1
X_5402_ _5357_/X _8040_/Q _5404_/S vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__mux2_1
X_6382_ _7818_/Q _6343_/X _6371_/X _6381_/X _6378_/X vssd1 vssd1 vccd1 vccd1 _7818_/D
+ sky130_fd_sc_hd__a221o_1
X_5333_ _8072_/Q _5331_/X _5332_/Y _5249_/X vssd1 vssd1 vccd1 vccd1 _8072_/D sky130_fd_sc_hd__o211a_1
X_8121_ _8478_/CLK _8121_/D vssd1 vssd1 vccd1 vccd1 _8121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8052_ _8052_/CLK _8052_/D vssd1 vssd1 vccd1 vccd1 _8052_/Q sky130_fd_sc_hd__dfxtp_1
X_5264_ _5056_/X _5260_/Y _5263_/Y _5031_/A vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__a31o_1
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3062_ _6272_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3062_/X sky130_fd_sc_hd__clkbuf_16
X_5195_ _5174_/X _5193_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__o21a_1
X_4215_ _8328_/Q _4147_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__mux2_1
X_4146_ _4146_/A vssd1 vssd1 vccd1 vccd1 _8353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _3937_/X _8367_/Q _4081_/S vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__mux2_1
X_7905_ _7905_/CLK _7905_/D vssd1 vssd1 vccd1 vccd1 _7905_/Q sky130_fd_sc_hd__dfxtp_1
X_7415__169 _7416__170/A vssd1 vssd1 vccd1 vccd1 _8380_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7836_ _8497_/CLK _7836_/D vssd1 vssd1 vccd1 vccd1 _7836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4979_ _8103_/Q _4978_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4980_/A sky130_fd_sc_hd__mux2_1
X_7767_ _8308_/CLK _7767_/D vssd1 vssd1 vccd1 vccd1 _7767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7698_ _7698_/A _7698_/B vssd1 vssd1 vccd1 vccd1 _7698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6649_ _6649_/A vssd1 vssd1 vccd1 vccd1 _7970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8319_ _8442_/CLK _8319_/D vssd1 vssd1 vccd1 vccd1 _8319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7143__104 _7144__105/A vssd1 vssd1 vccd1 vccd1 _8285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _8395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6724__359 _6725__360/A vssd1 vssd1 vccd1 vccd1 _8026_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5951_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4902_ _8132_/Q _4903_/A _4900_/X _4901_/Y vssd1 vssd1 vccd1 vccd1 _8132_/D sky130_fd_sc_hd__o211a_1
X_5882_ _7607_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__or2_1
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7621_ _7633_/A vssd1 vssd1 vccd1 vccd1 _7621_/X sky130_fd_sc_hd__buf_1
X_4833_ _4789_/X _7858_/Q _4803_/X _8091_/Q _4663_/A vssd1 vssd1 vccd1 vccd1 _4833_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4764_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__clkbuf_2
X_7552_ _7554_/A _7552_/B vssd1 vssd1 vccd1 vccd1 _8428_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7483_ _7484_/B _7484_/C _8486_/Q vssd1 vssd1 vccd1 vccd1 _7483_/Y sky130_fd_sc_hd__a21oi_1
X_4695_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4696_/S sky130_fd_sc_hd__buf_2
X_6434_ _6434_/A vssd1 vssd1 vccd1 vccd1 _7835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6365_ _6353_/X _6364_/X _6355_/X vssd1 vssd1 vccd1 vccd1 _6365_/X sky130_fd_sc_hd__o21a_1
X_8104_ _8104_/CLK _8104_/D vssd1 vssd1 vccd1 vccd1 _8104_/Q sky130_fd_sc_hd__dfxtp_1
X_6296_ _6296_/A _7658_/A vssd1 vssd1 vccd1 vccd1 _6297_/B sky130_fd_sc_hd__nor2_1
X_5316_ _5316_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5247_ _5231_/X _5245_/X _5338_/A vssd1 vssd1 vccd1 vccd1 _5247_/Y sky130_fd_sc_hd__o21ai_1
X_8035_ _8439_/CLK _8035_/D vssd1 vssd1 vccd1 vccd1 _8035_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3431_ clkbuf_0__3431_/X vssd1 vssd1 vccd1 vccd1 _7392_/A sky130_fd_sc_hd__clkbuf_4
X_5178_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__buf_2
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4129_ _4129_/A _4129_/B _4129_/C _4608_/A vssd1 vssd1 vccd1 vccd1 _7645_/B sky130_fd_sc_hd__or4b_2
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7819_ _8489_/CLK _7819_/D vssd1 vssd1 vccd1 vccd1 _7819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6827__372 _6827__372/A vssd1 vssd1 vccd1 vccd1 _8040_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3629_ clkbuf_0__3629_/X vssd1 vssd1 vccd1 vccd1 _7450__22/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7364__127 _7366__129/A vssd1 vssd1 vccd1 vccd1 _8338_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _8197_/Q _4229_/X _4486_/S vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6150_ _7774_/Q _7773_/Q vssd1 vssd1 vccd1 vccd1 _6231_/B sky130_fd_sc_hd__or2b_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _8464_/Q _8025_/Q _7990_/Q _8456_/Q _5063_/X _5064_/X vssd1 vssd1 vccd1 vccd1
+ _5101_/X sky130_fd_sc_hd__mux4_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7825_/Q input11/X _6107_/A vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__mux2_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _8069_/Q vssd1 vssd1 vccd1 vccd1 _5164_/A sky130_fd_sc_hd__buf_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8060_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6983_ _6989_/A vssd1 vssd1 vccd1 vccd1 _6983_/X sky130_fd_sc_hd__buf_1
X_5934_ _5934_/A vssd1 vssd1 vccd1 vccd1 _5934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6956__456 _6957__457/A vssd1 vssd1 vccd1 vccd1 _8135_/CLK sky130_fd_sc_hd__inv_2
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__clkbuf_1
X_4816_ _7946_/Q _4653_/B _4767_/X vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__a21o_1
X_7604_ _7604_/A _7604_/B _7604_/C vssd1 vssd1 vccd1 vccd1 _7605_/A sky130_fd_sc_hd__and3_1
X_6143__183 _6143__183/A vssd1 vssd1 vccd1 vccd1 _7732_/CLK sky130_fd_sc_hd__inv_2
X_5796_ _5796_/A vssd1 vssd1 vccd1 vccd1 _7792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4747_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__clkbuf_2
X_7535_ _7535_/A vssd1 vssd1 vccd1 vccd1 _7546_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7466_ _7465_/B _7465_/C _7492_/A vssd1 vssd1 vccd1 vccd1 _7466_/Y sky130_fd_sc_hd__a21oi_1
X_4678_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4678_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6417_ _8482_/Q vssd1 vssd1 vccd1 vccd1 _7503_/A sky130_fd_sc_hd__inv_2
X_6348_ _8478_/Q _6311_/A _6347_/X _6355_/B _6352_/A vssd1 vssd1 vccd1 vccd1 _6348_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput105 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _6642_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8018_ _8481_/CLK _8018_/D vssd1 vssd1 vccd1 vccd1 _8018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3414_ clkbuf_0__3414_/X vssd1 vssd1 vccd1 vccd1 _6988__480/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3276_ clkbuf_0__3276_/X vssd1 vssd1 vccd1 vccd1 _6685__332/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _8402_/D sky130_fd_sc_hd__clkbuf_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5650_ _5650_/A vssd1 vssd1 vccd1 vccd1 _7906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4601_ _4601_/A vssd1 vssd1 vccd1 vccd1 _8145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5581_ _5580_/X _7936_/Q _5581_/S vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A vssd1 vssd1 vccd1 vccd1 _8175_/D sky130_fd_sc_hd__clkbuf_1
X_7320_ _8315_/Q _7320_/B _7320_/C _7320_/D vssd1 vssd1 vccd1 vccd1 _7321_/C sky130_fd_sc_hd__or4_1
XFILLER_116_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4463_ _4350_/X _8204_/Q _4467_/S vssd1 vssd1 vccd1 vccd1 _4464_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _7972_/Q _6197_/X _6195_/X _6198_/X _7761_/Q vssd1 vssd1 vccd1 vccd1 _7761_/D
+ sky130_fd_sc_hd__o32a_1
X_4394_ _4353_/X _8227_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__mux2_1
X_7182_ _8488_/Q _7182_/B vssd1 vssd1 vccd1 vccd1 _7236_/B sky130_fd_sc_hd__xor2_1
X_6133_ _6559_/A vssd1 vssd1 vccd1 vccd1 _6133_/X sky130_fd_sc_hd__buf_1
XFILLER_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6064_ _6053_/X _6062_/X _6063_/X _6056_/X vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__o211a_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _8090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3061_ clkbuf_0__3061_/X vssd1 vssd1 vccd1 vccd1 _6268__202/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__or2_4
X_6897_ _6909_/A vssd1 vssd1 vccd1 vccd1 _6897_/X sky130_fd_sc_hd__buf_1
X_5848_ _5848_/A vssd1 vssd1 vccd1 vccd1 _7726_/D sky130_fd_sc_hd__clkbuf_1
X_5779_ _5779_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5795_/S sky130_fd_sc_hd__nor2_2
XFILLER_21_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _7517_/A _7516_/X _7517_/Y _7514_/X vssd1 vssd1 vccd1 vccd1 _8415_/D sky130_fd_sc_hd__o211a_1
XFILLER_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8498_ _8498_/CLK _8498_/D vssd1 vssd1 vccd1 vccd1 _8498_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6527__250 _6527__250/A vssd1 vssd1 vccd1 vccd1 _7890_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6820_ _7575_/A _7584_/B _6820_/C vssd1 vssd1 vccd1 vccd1 _6821_/A sky130_fd_sc_hd__and3_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _3963_/A vssd1 vssd1 vccd1 vccd1 _8408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6751_ _6751_/A vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__buf_2
X_5702_ _5702_/A vssd1 vssd1 vccd1 vccd1 _7883_/D sky130_fd_sc_hd__clkbuf_1
X_3894_ _3894_/A vssd1 vssd1 vccd1 vccd1 _8466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6131_/A sky130_fd_sc_hd__clkbuf_4
X_5633_ _7913_/Q _4993_/X _5635_/S vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__mux2_1
X_8421_ _8425_/CLK _8421_/D vssd1 vssd1 vccd1 vccd1 _8421_/Q sky130_fd_sc_hd__dfxtp_1
X_5564_ _5564_/A vssd1 vssd1 vccd1 vccd1 _7942_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3431_ _7075_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3431_/X sky130_fd_sc_hd__clkbuf_16
X_8352_ _8352_/CLK _8352_/D vssd1 vssd1 vccd1 vccd1 _8352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4515_ _4515_/A _4588_/A vssd1 vssd1 vccd1 vccd1 _4531_/S sky130_fd_sc_hd__or2_4
X_7303_ _8310_/Q _7295_/X _7272_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7304_/B sky130_fd_sc_hd__o2bb2a_1
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _7995_/D sky130_fd_sc_hd__clkbuf_1
X_8283_ _8283_/CLK _8283_/D vssd1 vssd1 vccd1 vccd1 _8283_/Q sky130_fd_sc_hd__dfxtp_1
X_4446_ _8210_/Q _4445_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__mux2_1
X_7234_ _7692_/A _7178_/B _7231_/Y _7232_/X _7233_/Y vssd1 vssd1 vccd1 vccd1 _7234_/X
+ sky130_fd_sc_hd__a2111o_1
X_4377_ _4377_/A vssd1 vssd1 vccd1 vccd1 _8235_/D sky130_fd_sc_hd__clkbuf_1
X_7165_ _7173_/A vssd1 vssd1 vccd1 vccd1 _7217_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _7760_/Q _6111_/X _6112_/X _6115_/X _6109_/X vssd1 vssd1 vccd1 vccd1 _6116_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6047_ _6085_/A vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _7998_/CLK _7998_/D vssd1 vssd1 vccd1 vccd1 _7998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6949_ _6976_/A vssd1 vssd1 vccd1 vccd1 _6949_/X sky130_fd_sc_hd__buf_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3629_ _7448_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3629_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput206 _6045_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
X_5280_ _5280_/A _5280_/B vssd1 vssd1 vccd1 vccd1 _5280_/Y sky130_fd_sc_hd__nand2_1
X_4300_ _3937_/X _8265_/Q _4304_/S vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4231_ _4231_/A vssd1 vssd1 vccd1 vccd1 _8295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4162_ _4162_/A vssd1 vssd1 vccd1 vccd1 _8348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4093_ _8360_/Q _4010_/X _4093_/S vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__mux2_1
X_7921_ _7921_/CLK _7921_/D vssd1 vssd1 vccd1 vccd1 _7921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7852_ _8060_/CLK _7852_/D vssd1 vssd1 vccd1 vccd1 _7852_/Q sky130_fd_sc_hd__dfxtp_1
X_7783_ _7783_/CLK _7783_/D vssd1 vssd1 vccd1 vccd1 _7783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _4995_/A vssd1 vssd1 vccd1 vccd1 _8098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6803_ _6803_/A _6803_/B vssd1 vssd1 vccd1 vccd1 _6803_/X sky130_fd_sc_hd__and2_1
X_3946_ _4287_/A vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__buf_2
X_8404_ _8404_/CLK _8404_/D vssd1 vssd1 vccd1 vccd1 _8404_/Q sky130_fd_sc_hd__dfxtp_1
X_3877_ _8447_/Q vssd1 vssd1 vccd1 vccd1 _3877_/X sky130_fd_sc_hd__buf_2
X_5616_ _5616_/A vssd1 vssd1 vccd1 vccd1 _7921_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3377_ clkbuf_0__3377_/X vssd1 vssd1 vccd1 vccd1 _6841__383/A sky130_fd_sc_hd__clkbuf_4
X_5547_ _7948_/Q _4984_/X _5549_/S vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__mux2_1
X_8335_ _8335_/CLK _8335_/D vssd1 vssd1 vccd1 vccd1 _8335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3414_ _6983_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3414_/X sky130_fd_sc_hd__clkbuf_16
X_8266_ _8266_/CLK _8266_/D vssd1 vssd1 vccd1 vccd1 _8266_/Q sky130_fd_sc_hd__dfxtp_1
X_5478_ _8002_/Q _4359_/A _5482_/S vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4429_ _4428_/X _8215_/Q _4429_/S vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__mux2_1
X_7217_ _7217_/A _7217_/B _7217_/C vssd1 vssd1 vccd1 vccd1 _7292_/A sky130_fd_sc_hd__nand3_1
Xclkbuf_0__3276_ _6683_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3276_/X sky130_fd_sc_hd__clkbuf_16
X_8197_ _8197_/CLK _8197_/D vssd1 vssd1 vccd1 vccd1 _8197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7148_ _8300_/Q _8299_/Q _8298_/Q _8297_/Q vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__and4_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8520__219 vssd1 vssd1 vccd1 vccd1 _8520__219/HI core0Index[6] sky130_fd_sc_hd__conb_1
XFILLER_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6975__470 _6975__470/A vssd1 vssd1 vccd1 vccd1 _8151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6570__284 _6571__285/A vssd1 vssd1 vccd1 vccd1 _7924_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4780_ _4780_/A vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3231_ clkbuf_0__3231_/X vssd1 vssd1 vccd1 vccd1 _6578_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6450_ _6450_/A vssd1 vssd1 vccd1 vccd1 _7842_/D sky130_fd_sc_hd__clkbuf_1
X_5401_ _5401_/A vssd1 vssd1 vccd1 vccd1 _8041_/D sky130_fd_sc_hd__clkbuf_1
X_6381_ _7692_/A _6390_/B _6387_/C vssd1 vssd1 vccd1 vccd1 _6381_/X sky130_fd_sc_hd__and3_1
X_5332_ _5338_/A _5332_/B vssd1 vssd1 vccd1 vccd1 _5332_/Y sky130_fd_sc_hd__nand2_1
X_8120_ _8120_/CLK _8120_/D vssd1 vssd1 vccd1 vccd1 _8120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8051_ _8051_/CLK _8051_/D vssd1 vssd1 vccd1 vccd1 _8051_/Q sky130_fd_sc_hd__dfxtp_1
X_5263_ _5174_/X _5261_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _5263_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3061_ _6266_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3061_/X sky130_fd_sc_hd__clkbuf_16
X_5194_ _8368_/Q _5178_/X _5179_/X _8360_/Q _5037_/A vssd1 vssd1 vccd1 vccd1 _5194_/X
+ sky130_fd_sc_hd__o221a_1
X_4214_ _4214_/A vssd1 vssd1 vccd1 vccd1 _8329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _8353_/Q _4144_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4076_ _4076_/A vssd1 vssd1 vccd1 vccd1 _8368_/D sky130_fd_sc_hd__clkbuf_1
X_7904_ _7904_/CLK _7904_/D vssd1 vssd1 vccd1 vccd1 _7904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7835_ _8497_/CLK _7835_/D vssd1 vssd1 vccd1 vccd1 _7835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4978_ _8066_/Q vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__clkbuf_4
X_7766_ _8308_/CLK _7766_/D vssd1 vssd1 vccd1 vccd1 _7766_/Q sky130_fd_sc_hd__dfxtp_1
X_3929_ _3928_/X _8455_/Q _3935_/S vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__mux2_1
X_7697_ _7695_/Y _7696_/Y _6194_/X vssd1 vssd1 vccd1 vccd1 _8490_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1_0__3429_ clkbuf_0__3429_/X vssd1 vssd1 vccd1 vccd1 _7064__541/A sky130_fd_sc_hd__clkbuf_4
X_6648_ _7970_/Q _5933_/A _6652_/S vssd1 vssd1 vccd1 vccd1 _6649_/A sky130_fd_sc_hd__mux2_1
X_7129__93 _7131__95/A vssd1 vssd1 vccd1 vccd1 _8274_/CLK sky130_fd_sc_hd__inv_2
X_8318_ _8442_/CLK _8318_/D vssd1 vssd1 vccd1 vccd1 _8318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8249_ _8249_/CLK _8249_/D vssd1 vssd1 vccd1 vccd1 _8249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7447__20 _7447__20/A vssd1 vssd1 vccd1 vccd1 _8406_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7003__492 _7004__493/A vssd1 vssd1 vccd1 vccd1 _8173_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8542__241 vssd1 vssd1 vccd1 vccd1 _8542__241/HI partID[5] sky130_fd_sc_hd__conb_1
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5950_ _5950_/A vssd1 vssd1 vccd1 vccd1 _5950_/X sky130_fd_sc_hd__clkbuf_1
X_6282__214 _6282__214/A vssd1 vssd1 vccd1 vccd1 _7806_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4901_ _4911_/C vssd1 vssd1 vccd1 vccd1 _4901_/Y sky130_fd_sc_hd__inv_2
X_5881_ _5881_/A vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__clkbuf_1
X_4832_ _4801_/X _7978_/Q _7882_/Q _4769_/X _4794_/A vssd1 vssd1 vccd1 vccd1 _4832_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ _4760_/X _7915_/Q _4762_/X _7923_/Q _4715_/X vssd1 vssd1 vccd1 vccd1 _4763_/X
+ sky130_fd_sc_hd__o221a_1
X_7551_ _8428_/Q _7510_/B _7544_/X _7498_/B vssd1 vssd1 vccd1 vccd1 _7552_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__clkbuf_2
X_7482_ _8490_/Q _7492_/B _7477_/X _7478_/Y _7481_/X vssd1 vssd1 vccd1 vccd1 _7486_/C
+ sky130_fd_sc_hd__a2111o_1
X_6433_ _7835_/Q _5958_/A _6433_/S vssd1 vssd1 vccd1 vccd1 _6434_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6364_ _4608_/A _4608_/B _8017_/Q _6292_/B vssd1 vssd1 vccd1 vccd1 _6364_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8103_ _8103_/CLK _8103_/D vssd1 vssd1 vccd1 vccd1 _8103_/Q sky130_fd_sc_hd__dfxtp_1
X_7421__174 _7422__175/A vssd1 vssd1 vccd1 vccd1 _8385_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6295_ _7831_/Q _7839_/Q _7840_/Q vssd1 vssd1 vccd1 vccd1 _7658_/A sky130_fd_sc_hd__or3_1
X_5315_ _8078_/Q _5087_/A _4025_/B _5282_/X vssd1 vssd1 vccd1 vccd1 _8078_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8034_ _8034_/CLK _8034_/D vssd1 vssd1 vccd1 vccd1 _8034_/Q sky130_fd_sc_hd__dfxtp_1
X_5246_ _5246_/A vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5177_ _8408_/Q _8146_/Q _5301_/S vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _8127_/Q _4781_/A _4114_/Y vssd1 vssd1 vccd1 vccd1 _4608_/A sky130_fd_sc_hd__o21ai_2
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4059_ _4059_/A vssd1 vssd1 vccd1 vccd1 _8375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6521__245 _6521__245/A vssd1 vssd1 vccd1 vccd1 _7885_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _8017_/CLK _7818_/D vssd1 vssd1 vccd1 vccd1 _7818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7749_ _8483_/CLK _7749_/D vssd1 vssd1 vccd1 vccd1 _7749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8526__225 vssd1 vssd1 vccd1 vccd1 _8526__225/HI core1Index[5] sky130_fd_sc_hd__conb_1
X_6682__330 _6682__330/A vssd1 vssd1 vccd1 vccd1 _7994_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6834__377 _6836__379/A vssd1 vssd1 vccd1 vccd1 _8045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6988__480 _6988__480/A vssd1 vssd1 vccd1 vccd1 _8161_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730__364 _6731__365/A vssd1 vssd1 vccd1 vccd1 _8031_/CLK sky130_fd_sc_hd__inv_2
X_7123__88 _7123__88/A vssd1 vssd1 vccd1 vccd1 _8269_/CLK sky130_fd_sc_hd__inv_2
X_5100_ _7798_/Q _8006_/Q _8285_/Q _8033_/Q _5060_/X _5052_/X vssd1 vssd1 vccd1 vccd1
+ _5100_/X sky130_fd_sc_hd__mux4_1
X_6080_ _6080_/A vssd1 vssd1 vccd1 vccd1 _6107_/A sky130_fd_sc_hd__buf_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__clkbuf_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7441__15 _7441__15/A vssd1 vssd1 vccd1 vccd1 _8401_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6982_ _7044_/A vssd1 vssd1 vccd1 vccd1 _6982_/X sky130_fd_sc_hd__buf_1
X_5933_ _5933_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__or2_1
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5864_ _6207_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__and2_1
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4815_ _4760_/X _7914_/Q _4814_/X _7922_/Q _4715_/X vssd1 vssd1 vccd1 vccd1 _4815_/X
+ sky130_fd_sc_hd__o221a_1
X_7603_ _7603_/A _7675_/B vssd1 vssd1 vccd1 vccd1 _7604_/C sky130_fd_sc_hd__and2_1
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5795_ _7792_/Q _4365_/A _5795_/S vssd1 vssd1 vccd1 vccd1 _5796_/A sky130_fd_sc_hd__mux2_1
X_7534_ _7534_/A _7534_/B vssd1 vssd1 vccd1 vccd1 _8420_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4746_ _4746_/A vssd1 vssd1 vccd1 vccd1 _4926_/B sky130_fd_sc_hd__clkbuf_2
X_7465_ _7492_/A _7465_/B _7465_/C vssd1 vssd1 vccd1 vccd1 _7465_/X sky130_fd_sc_hd__and3_1
X_4677_ _4903_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _4678_/A sky130_fd_sc_hd__and2_1
XFILLER_103_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6416_ _8483_/Q vssd1 vssd1 vccd1 vccd1 _6419_/A sky130_fd_sc_hd__inv_2
XFILLER_1_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6347_ _8138_/Q _6318_/A _6319_/X vssd1 vssd1 vccd1 vccd1 _6347_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3059_ clkbuf_0__3059_/X vssd1 vssd1 vccd1 vccd1 _6264__200/A sky130_fd_sc_hd__clkbuf_4
X_6278_ _6278_/A vssd1 vssd1 vccd1 vccd1 _6278_/X sky130_fd_sc_hd__buf_1
Xinput106 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__buf_6
X_5229_ _5224_/A _5226_/X _5228_/X _5048_/X vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__o211a_1
X_8017_ _8017_/CLK _8017_/D vssd1 vssd1 vccd1 vccd1 _8017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3413_ clkbuf_0__3413_/X vssd1 vssd1 vccd1 vccd1 _7007_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6681__329/A sky130_fd_sc_hd__clkbuf_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7370__132 _7370__132/A vssd1 vssd1 vccd1 vccd1 _8343_/CLK sky130_fd_sc_hd__inv_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _8145_/Q _4448_/X _4604_/S vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__mux2_1
X_5580_ _5580_/A vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__clkbuf_2
X_4531_ _4365_/X _8175_/Q _4531_/S vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4462_ _4462_/A vssd1 vssd1 vccd1 vccd1 _8205_/D sky130_fd_sc_hd__clkbuf_1
X_7250_ _7349_/A vssd1 vssd1 vccd1 vccd1 _7250_/X sky130_fd_sc_hd__buf_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6201_ _7971_/Q _6197_/X _6195_/X _6198_/X _7760_/Q vssd1 vssd1 vccd1 vccd1 _7760_/D
+ sky130_fd_sc_hd__o32a_1
X_4393_ _4393_/A vssd1 vssd1 vccd1 vccd1 _8228_/D sky130_fd_sc_hd__clkbuf_1
X_7181_ _7181_/A _7181_/B vssd1 vssd1 vccd1 vccd1 _7182_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6132_ _6915_/A vssd1 vssd1 vccd1 vccd1 _6132_/X sky130_fd_sc_hd__buf_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6063_ _7745_/Q _6063_/B vssd1 vssd1 vccd1 vccd1 _6063_/X sky130_fd_sc_hd__or2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6962__461 _6968__464/A vssd1 vssd1 vccd1 vccd1 _8140_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _4425_/X _8090_/Q _5016_/S vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7058__536 _7059__537/A vssd1 vssd1 vccd1 vccd1 _8217_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7603_/A _6242_/X _6353_/X _6194_/X vssd1 vssd1 vccd1 vccd1 _8142_/D sky130_fd_sc_hd__a211oi_1
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _5916_/A vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3060_ clkbuf_0__3060_/X vssd1 vssd1 vccd1 vccd1 _6491_/A sky130_fd_sc_hd__clkbuf_4
X_6896_ _6896_/A vssd1 vssd1 vccd1 vccd1 _8088_/D sky130_fd_sc_hd__clkbuf_1
X_5847_ _4153_/X _7726_/Q _5849_/S vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5778_ _5778_/A vssd1 vssd1 vccd1 vccd1 _7800_/D sky130_fd_sc_hd__clkbuf_1
X_4729_ _4930_/B _4726_/X _4728_/X vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__a21o_1
X_7517_ _7517_/A _7517_/B vssd1 vssd1 vccd1 vccd1 _7517_/Y sky130_fd_sc_hd__nand2_1
X_8497_ _8497_/CLK _8497_/D vssd1 vssd1 vccd1 vccd1 _8497_/Q sky130_fd_sc_hd__dfxtp_2
X_7448_ _7448_/A vssd1 vssd1 vccd1 vccd1 _7448_/X sky130_fd_sc_hd__buf_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7638__45 _7638__45/A vssd1 vssd1 vccd1 vccd1 _8468_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898__411 _6900__413/A vssd1 vssd1 vccd1 vccd1 _8089_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6534__255 _6534__255/A vssd1 vssd1 vccd1 vccd1 _7895_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6750_ _8427_/Q _6808_/A _6808_/B _6808_/C vssd1 vssd1 vccd1 vccd1 _7484_/B sky130_fd_sc_hd__nand4_1
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ _8408_/Q _3883_/X _3962_/S vssd1 vssd1 vccd1 vccd1 _3963_/A sky130_fd_sc_hd__mux2_1
X_5701_ _7883_/Q _4987_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__mux2_1
X_3893_ _8466_/Q _3892_/X _3893_/S vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__mux2_1
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _7914_/D sky130_fd_sc_hd__clkbuf_1
X_8420_ _8425_/CLK _8420_/D vssd1 vssd1 vccd1 vccd1 _8420_/Q sky130_fd_sc_hd__dfxtp_1
X_5563_ _5562_/X _7942_/Q _5572_/S vssd1 vssd1 vccd1 vccd1 _5564_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3430_ _7069_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3430_/X sky130_fd_sc_hd__clkbuf_16
X_8351_ _8351_/CLK _8351_/D vssd1 vssd1 vccd1 vccd1 _8351_/Q sky130_fd_sc_hd__dfxtp_1
X_4514_ _4514_/A vssd1 vssd1 vccd1 vccd1 _8183_/D sky130_fd_sc_hd__clkbuf_1
X_7302_ _7309_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _8309_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5494_ _5361_/X _7995_/Q _5494_/S vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__mux2_1
X_8282_ _8282_/CLK _8282_/D vssd1 vssd1 vccd1 vccd1 _8282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ _8445_/Q vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__clkbuf_4
X_7233_ _7232_/B _7232_/C _7468_/A vssd1 vssd1 vccd1 vccd1 _7233_/Y sky130_fd_sc_hd__a21oi_1
X_4376_ _4353_/X _8235_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__mux2_1
X_7164_ _7211_/C vssd1 vssd1 vccd1 vccd1 _7217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7377__138 _7379__140/A vssd1 vssd1 vccd1 vccd1 _8349_/CLK sky130_fd_sc_hd__inv_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6115_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6115_/X sky130_fd_sc_hd__and2_1
X_7095_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7095_/X sky130_fd_sc_hd__buf_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6046_ _7816_/Q input33/X _6058_/S vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__mux2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _7997_/CLK _7997_/D vssd1 vssd1 vccd1 vccd1 _7997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6948_ _7044_/A vssd1 vssd1 vccd1 vccd1 _6948_/X sky130_fd_sc_hd__buf_1
X_6879_ _6879_/A vssd1 vssd1 vccd1 vccd1 _6879_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3628_ _7442_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3628_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput207 _6049_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _8295_/Q _4229_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4161_ _8348_/Q _3992_/X _4169_/S vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__mux2_1
X_8506__256 vssd1 vssd1 vccd1 vccd1 partID[10] _8506__256/LO sky130_fd_sc_hd__conb_1
X_4092_ _4092_/A vssd1 vssd1 vccd1 vccd1 _8361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7920_ _7920_/CLK _7920_/D vssd1 vssd1 vccd1 vccd1 _7920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7851_ _8060_/CLK _7851_/D vssd1 vssd1 vccd1 vccd1 _7851_/Q sky130_fd_sc_hd__dfxtp_1
X_6802_ _6802_/A _7462_/B vssd1 vssd1 vccd1 vccd1 _6803_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7782_ _7782_/CLK _7782_/D vssd1 vssd1 vccd1 vccd1 _7782_/Q sky130_fd_sc_hd__dfxtp_1
X_4994_ _8098_/Q _4993_/X _4997_/S vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3945_ _3945_/A vssd1 vssd1 vccd1 vccd1 _8450_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3445_ clkbuf_0__3445_/X vssd1 vssd1 vccd1 vccd1 _7144__105/A sky130_fd_sc_hd__clkbuf_4
X_6664_ _6670_/A vssd1 vssd1 vccd1 vccd1 _6664_/X sky130_fd_sc_hd__buf_1
X_5615_ _5577_/X _7921_/Q _5617_/S vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__mux2_1
X_3876_ _3876_/A vssd1 vssd1 vccd1 vccd1 _8472_/D sky130_fd_sc_hd__clkbuf_1
X_8403_ _8403_/CLK _8403_/D vssd1 vssd1 vccd1 vccd1 _8403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3376_ clkbuf_0__3376_/X vssd1 vssd1 vccd1 vccd1 _6837__380/A sky130_fd_sc_hd__clkbuf_4
X_5546_ _5546_/A vssd1 vssd1 vccd1 vccd1 _7949_/D sky130_fd_sc_hd__clkbuf_1
X_8334_ _8334_/CLK _8334_/D vssd1 vssd1 vccd1 vccd1 _8334_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3413_ _6982_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3413_/X sky130_fd_sc_hd__clkbuf_16
X_5477_ _5477_/A vssd1 vssd1 vccd1 vccd1 _8003_/D sky130_fd_sc_hd__clkbuf_1
X_8265_ _8265_/CLK _8265_/D vssd1 vssd1 vccd1 vccd1 _8265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7216_ _8490_/Q _7216_/B _7292_/B vssd1 vssd1 vccd1 vccd1 _7216_/X sky130_fd_sc_hd__or3b_1
X_4428_ _8060_/Q vssd1 vssd1 vccd1 vccd1 _4428_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3275_ _6677_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3275_/X sky130_fd_sc_hd__clkbuf_16
X_8196_ _8196_/CLK _8196_/D vssd1 vssd1 vccd1 vccd1 _8196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4359_ _4359_/A vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__clkbuf_2
X_7147_ _8315_/Q _8314_/Q _7317_/B _8288_/Q vssd1 vssd1 vccd1 vccd1 _7311_/B sky130_fd_sc_hd__and4_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6029_ _7736_/Q _6044_/B vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__or2_1
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_90 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7015__501 _7015__501/A vssd1 vssd1 vccd1 vccd1 _8182_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3230_ clkbuf_0__3230_/X vssd1 vssd1 vccd1 vccd1 _6554__271/A sky130_fd_sc_hd__clkbuf_4
X_5400_ _5353_/X _8041_/Q _5404_/S vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__mux2_1
X_6380_ _8489_/Q vssd1 vssd1 vccd1 vccd1 _7692_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5331_ _5331_/A vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8050_ _8050_/CLK _8050_/D vssd1 vssd1 vccd1 vccd1 _8050_/Q sky130_fd_sc_hd__dfxtp_1
X_5262_ _8264_/Q _5214_/A _5179_/X _8256_/Q _5037_/A vssd1 vssd1 vccd1 vccd1 _5262_/X
+ sky130_fd_sc_hd__o221a_1
X_7001_ _7007_/A vssd1 vssd1 vccd1 vccd1 _7001_/X sky130_fd_sc_hd__buf_1
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3060_ _6265_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3060_/X sky130_fd_sc_hd__clkbuf_16
X_5193_ _8336_/Q _8344_/Q _5301_/S vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4213_ _8329_/Q _4144_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__mux2_1
X_4144_ _8064_/Q vssd1 vssd1 vccd1 vccd1 _4144_/X sky130_fd_sc_hd__buf_2
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4075_ _3934_/X _8368_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4076_/A sky130_fd_sc_hd__mux2_1
X_7903_ _7903_/CLK _7903_/D vssd1 vssd1 vccd1 vccd1 _7903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7834_ _8497_/CLK _7834_/D vssd1 vssd1 vccd1 vccd1 _7834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7765_ _8308_/CLK _7765_/D vssd1 vssd1 vccd1 vccd1 _7765_/Q sky130_fd_sc_hd__dfxtp_1
X_4977_ _4977_/A vssd1 vssd1 vccd1 vccd1 _8104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7696_ _7696_/A _7699_/B vssd1 vssd1 vccd1 vccd1 _7696_/Y sky130_fd_sc_hd__nand2_1
X_3928_ _8447_/Q vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__buf_4
X_6647_ _6647_/A vssd1 vssd1 vccd1 vccd1 _7969_/D sky130_fd_sc_hd__clkbuf_1
X_3859_ _7842_/Q _7843_/Q _7844_/Q _7841_/Q vssd1 vssd1 vccd1 vccd1 _7652_/D sky130_fd_sc_hd__or4b_1
Xclkbuf_1_1_0__3428_ clkbuf_0__3428_/X vssd1 vssd1 vccd1 vccd1 _7062__540/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578_ _6578_/A vssd1 vssd1 vccd1 vccd1 _6578_/X sky130_fd_sc_hd__buf_1
X_5529_ _5529_/A vssd1 vssd1 vccd1 vccd1 _7980_/D sky130_fd_sc_hd__clkbuf_1
X_8317_ _8442_/CLK _8317_/D vssd1 vssd1 vccd1 vccd1 _8317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8248_ _8248_/CLK _8248_/D vssd1 vssd1 vccd1 vccd1 _8248_/Q sky130_fd_sc_hd__dfxtp_1
X_8179_ _8179_/CLK _8179_/D vssd1 vssd1 vccd1 vccd1 _8179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5880_ _7603_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__or2_1
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4900_ _6854_/A vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__buf_2
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4831_ _4932_/B _4829_/X _4830_/X vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4762_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7550_ _7554_/A _7550_/B vssd1 vssd1 vccd1 vccd1 _8427_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4693_ _8103_/Q _8058_/Q _7942_/Q _8295_/Q _4648_/A _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4693_/X sky130_fd_sc_hd__mux4_1
X_7481_ _7479_/X _7480_/Y _6768_/A _7478_/B vssd1 vssd1 vccd1 vccd1 _7481_/X sky130_fd_sc_hd__a2bb2o_1
X_6432_ _6432_/A vssd1 vssd1 vccd1 vccd1 _7834_/D sky130_fd_sc_hd__clkbuf_1
X_8102_ _8102_/CLK _8102_/D vssd1 vssd1 vccd1 vccd1 _8102_/Q sky130_fd_sc_hd__dfxtp_1
X_6363_ _6289_/X _6361_/X _6362_/X vssd1 vssd1 vccd1 vccd1 _7815_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6294_ _6294_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__or2b_1
X_5314_ _3943_/X _5022_/A _5313_/X _5282_/X vssd1 vssd1 vccd1 vccd1 _8079_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8033_ _8033_/CLK _8033_/D vssd1 vssd1 vccd1 vccd1 _8033_/Q sky130_fd_sc_hd__dfxtp_1
X_5245_ _5334_/B _5234_/X _5237_/X _5244_/X _5031_/X vssd1 vssd1 vccd1 vccd1 _5245_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5176_ _5307_/S vssd1 vssd1 vccd1 vccd1 _5301_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_56_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4127_ _4127_/A vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__buf_2
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4058_ _8375_/Q _4014_/X _4062_/S vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6595__303 _6595__303/A vssd1 vssd1 vccd1 vccd1 _7943_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7817_ _8017_/CLK _7817_/D vssd1 vssd1 vccd1 vccd1 _7817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7748_ _7964_/CLK _7748_/D vssd1 vssd1 vccd1 vccd1 _7748_/Q sky130_fd_sc_hd__dfxtp_1
X_7679_ _7674_/Y _7677_/Y _7678_/X vssd1 vssd1 vccd1 vccd1 _8484_/D sky130_fd_sc_hd__a21oi_1
XFILLER_106_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3627_ clkbuf_0__3627_/X vssd1 vssd1 vccd1 vccd1 _7439__13/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _8072_/Q _5084_/B vssd1 vssd1 vccd1 vccd1 _5031_/A sky130_fd_sc_hd__xor2_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6583__295 _6583__295/A vssd1 vssd1 vccd1 vccd1 _7935_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5932_ _5932_/A vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5863_ _5863_/A vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__buf_2
X_5794_ _5794_/A vssd1 vssd1 vccd1 vccd1 _7793_/D sky130_fd_sc_hd__clkbuf_1
X_7602_ _7602_/A vssd1 vssd1 vccd1 vccd1 _8443_/D sky130_fd_sc_hd__clkbuf_1
X_7533_ _7471_/B _7471_/C _7516_/X _7522_/X _8420_/Q vssd1 vssd1 vccd1 vccd1 _7534_/B
+ sky130_fd_sc_hd__a32oi_1
X_4745_ _4745_/A vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4676_ _4622_/X _4646_/X _4657_/X _4675_/X vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__a31o_1
X_7464_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _7492_/A sky130_fd_sc_hd__inv_2
X_8549__248 vssd1 vssd1 vccd1 vccd1 _8549__248/HI versionID[2] sky130_fd_sc_hd__conb_1
X_6415_ _6294_/A _6415_/B vssd1 vssd1 vccd1 vccd1 _6415_/X sky130_fd_sc_hd__and2b_1
X_6346_ _7478_/A _6293_/A _6355_/A vssd1 vssd1 vccd1 vccd1 _6346_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3058_ clkbuf_0__3058_/X vssd1 vssd1 vccd1 vccd1 _6254__191/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput107 wbs_we_i vssd1 vssd1 vccd1 vccd1 _6228_/C sky130_fd_sc_hd__buf_6
X_8016_ _8498_/CLK _8016_/D vssd1 vssd1 vccd1 vccd1 _8016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5228_ _8233_/Q _5227_/X _5239_/B _8468_/Q vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__o22a_1
X_5159_ _5159_/A vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3412_ clkbuf_0__3412_/X vssd1 vssd1 vccd1 vccd1 _6979__473/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900__413 _6900__413/A vssd1 vssd1 vccd1 vccd1 _8091_/CLK sky130_fd_sc_hd__inv_2
X_6603__310 _6603__310/A vssd1 vssd1 vccd1 vccd1 _7950_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6701_/A sky130_fd_sc_hd__clkbuf_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840__382 _6841__383/A vssd1 vssd1 vccd1 vccd1 _8050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _4530_/A vssd1 vssd1 vccd1 vccd1 _8176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ _4347_/X _8205_/Q _4467_/S vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7180_ _8307_/Q _7193_/B _7193_/C _7217_/C _8308_/Q vssd1 vssd1 vccd1 vccd1 _7181_/B
+ sky130_fd_sc_hd__a41o_1
X_6200_ _7970_/Q _6197_/X _6195_/X _6198_/X _7759_/Q vssd1 vssd1 vccd1 vccd1 _7759_/D
+ sky130_fd_sc_hd__o32a_1
X_4392_ _4350_/X _8228_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__mux2_1
X_6131_ _6131_/A vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__buf_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6062_ _7820_/Q input6/X _6077_/S vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__mux2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5013_/A vssd1 vssd1 vccd1 vccd1 _8091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6964_/A vssd1 vssd1 vccd1 vccd1 _8141_/D sky130_fd_sc_hd__clkbuf_1
X_5915_ _5915_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__or2_4
X_6895_ _8324_/Q _7604_/A _6895_/C _6963_/A vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__and4b_1
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5846_ _5846_/A vssd1 vssd1 vccd1 vccd1 _7727_/D sky130_fd_sc_hd__clkbuf_1
X_5777_ _4156_/X _7800_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4728_ _4663_/X _4727_/X _4883_/A vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__a21o_1
X_7516_ _7491_/X _7490_/A _7577_/B _7572_/C vssd1 vssd1 vccd1 vccd1 _7516_/X sky130_fd_sc_hd__a22o_2
X_8496_ _8496_/CLK _8496_/D vssd1 vssd1 vccd1 vccd1 _8496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4659_ _4659_/A vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _6289_/X _6325_/X _6327_/X _6369_/A vssd1 vssd1 vccd1 vccd1 _6329_/X sky130_fd_sc_hd__a31o_1
XFILLER_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6907__419 _6908__420/A vssd1 vssd1 vccd1 vccd1 _8097_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _8409_/D sky130_fd_sc_hd__clkbuf_1
X_5700_ _5700_/A vssd1 vssd1 vccd1 vccd1 _7884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3892_ _8442_/Q vssd1 vssd1 vccd1 vccd1 _3892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5631_ _7914_/Q _4990_/X _5635_/S vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3392_ clkbuf_0__3392_/X vssd1 vssd1 vccd1 vccd1 _6887__406/A sky130_fd_sc_hd__clkbuf_4
X_5562_ _5562_/A vssd1 vssd1 vccd1 vccd1 _5562_/X sky130_fd_sc_hd__clkbuf_2
X_8350_ _8350_/CLK _8350_/D vssd1 vssd1 vccd1 vccd1 _8350_/Q sky130_fd_sc_hd__dfxtp_1
X_4513_ _8183_/Q _4247_/X _4513_/S vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__mux2_1
X_8281_ _8281_/CLK _8281_/D vssd1 vssd1 vccd1 vccd1 _8281_/Q sky130_fd_sc_hd__dfxtp_1
X_7301_ _8309_/Q _7295_/X _7272_/A _7195_/Y vssd1 vssd1 vccd1 vccd1 _7302_/B sky130_fd_sc_hd__o2bb2a_1
X_5493_ _5493_/A vssd1 vssd1 vccd1 vccd1 _7996_/D sky130_fd_sc_hd__clkbuf_1
X_7232_ _7468_/A _7232_/B _7232_/C vssd1 vssd1 vccd1 vccd1 _7232_/X sky130_fd_sc_hd__and3_1
XFILLER_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4444_ _4444_/A vssd1 vssd1 vccd1 vccd1 _8211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7064__541 _7064__541/A vssd1 vssd1 vccd1 vccd1 _8222_/CLK sky130_fd_sc_hd__inv_2
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _8236_/D sky130_fd_sc_hd__clkbuf_1
X_7163_ _7176_/A vssd1 vssd1 vccd1 vccd1 _7211_/C sky130_fd_sc_hd__clkbuf_2
X_6847__388 _6849__390/A vssd1 vssd1 vccd1 vccd1 _8056_/CLK sky130_fd_sc_hd__inv_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _7759_/Q _6111_/X _6112_/X _6113_/X _6109_/X vssd1 vssd1 vccd1 vccd1 _6114_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6045_ _6034_/X _6043_/X _6044_/X _6037_/X vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__o211a_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6704__348 _6706__350/A vssd1 vssd1 vccd1 vccd1 _8012_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _7996_/CLK _7996_/D vssd1 vssd1 vccd1 vccd1 _7996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5829_ _7777_/Q _5577_/A _5831_/S vssd1 vssd1 vccd1 vccd1 _5830_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3627_ _7436_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3627_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8479_ _8483_/CLK _8479_/D vssd1 vssd1 vccd1 vccd1 _8479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6540__260 _6540__260/A vssd1 vssd1 vccd1 vccd1 _7900_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput208 _6052_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_5_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4175_/S vssd1 vssd1 vccd1 vccd1 _4169_/S sky130_fd_sc_hd__buf_2
XFILLER_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7617__27 _7619__29/A vssd1 vssd1 vccd1 vccd1 _8450_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4091_ _8361_/Q _4006_/X _4093_/S vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7850_ _8141_/CLK _7850_/D vssd1 vssd1 vccd1 vccd1 _7850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6801_ _6800_/Y _6757_/A _6797_/B vssd1 vssd1 vccd1 vccd1 _7462_/B sky130_fd_sc_hd__a21bo_1
X_7781_ _7781_/CLK _7781_/D vssd1 vssd1 vccd1 vccd1 _7781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _8061_/Q vssd1 vssd1 vccd1 vccd1 _4993_/X sky130_fd_sc_hd__buf_2
X_6732_ _6825_/A vssd1 vssd1 vccd1 vccd1 _6732_/X sky130_fd_sc_hd__buf_1
X_3944_ _3943_/X _8450_/Q _3944_/S vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3875_ _8472_/Q _3874_/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3876_/A sky130_fd_sc_hd__mux2_1
X_5614_ _5614_/A vssd1 vssd1 vccd1 vccd1 _7922_/D sky130_fd_sc_hd__clkbuf_1
X_8402_ _8402_/CLK _8402_/D vssd1 vssd1 vccd1 vccd1 _8402_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3375_ clkbuf_0__3375_/X vssd1 vssd1 vccd1 vccd1 _6844_/A sky130_fd_sc_hd__clkbuf_4
X_7383__143 _7384__144/A vssd1 vssd1 vccd1 vccd1 _8354_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3412_ _6976_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3412_/X sky130_fd_sc_hd__clkbuf_16
X_5545_ _7949_/Q _4981_/X _5549_/S vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__mux2_1
X_8333_ _8333_/CLK _8333_/D vssd1 vssd1 vccd1 vccd1 _8333_/Q sky130_fd_sc_hd__dfxtp_1
X_5476_ _8003_/Q _4356_/A _5476_/S vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__mux2_1
X_8264_ _8264_/CLK _8264_/D vssd1 vssd1 vccd1 vccd1 _8264_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3274_ _6676_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3274_/X sky130_fd_sc_hd__clkbuf_16
X_8195_ _8195_/CLK _8195_/D vssd1 vssd1 vccd1 vccd1 _8195_/Q sky130_fd_sc_hd__dfxtp_1
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _8216_/D sky130_fd_sc_hd__clkbuf_1
X_7215_ _7184_/A _7176_/A _7193_/C _8306_/Q vssd1 vssd1 vccd1 vccd1 _7292_/B sky130_fd_sc_hd__a31o_1
X_7146_ _7345_/S vssd1 vssd1 vccd1 vccd1 _7331_/A sky130_fd_sc_hd__clkbuf_2
X_4358_ _4358_/A vssd1 vssd1 vccd1 vccd1 _8242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _7083_/A vssd1 vssd1 vccd1 vccd1 _7077_/X sky130_fd_sc_hd__buf_1
X_4289_ _4304_/S vssd1 vssd1 vccd1 vccd1 _4298_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6028_ _6085_/A vssd1 vssd1 vccd1 vccd1 _6044_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_104_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ _7979_/CLK _7979_/D vssd1 vssd1 vccd1 vccd1 _7979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_80 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_91 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5330_/A vssd1 vssd1 vccd1 vccd1 _8073_/D sky130_fd_sc_hd__clkbuf_1
X_5261_ _8240_/Q _8248_/Q _5261_/S vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4212_ _4212_/A vssd1 vssd1 vccd1 vccd1 _8330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5192_ _8392_/Q _5189_/X _5152_/A _5191_/X vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__o211a_1
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4143_ _4143_/A vssd1 vssd1 vccd1 vccd1 _8354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4074_ _4074_/A vssd1 vssd1 vccd1 vccd1 _8369_/D sky130_fd_sc_hd__clkbuf_1
X_7902_ _7902_/CLK _7902_/D vssd1 vssd1 vccd1 vccd1 _7902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7833_ _8497_/CLK _7833_/D vssd1 vssd1 vccd1 vccd1 _7833_/Q sky130_fd_sc_hd__dfxtp_1
X_7764_ _8433_/CLK _7764_/D vssd1 vssd1 vccd1 vccd1 _7764_/Q sky130_fd_sc_hd__dfxtp_1
X_4976_ _8104_/Q _4973_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__mux2_1
X_6715_ _6715_/A vssd1 vssd1 vccd1 vccd1 _8018_/D sky130_fd_sc_hd__clkbuf_1
X_3927_ _3927_/A vssd1 vssd1 vccd1 vccd1 _8456_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3427_ clkbuf_0__3427_/X vssd1 vssd1 vccd1 vccd1 _7054__533/A sky130_fd_sc_hd__clkbuf_4
X_7695_ _8490_/Q _7698_/B vssd1 vssd1 vccd1 vccd1 _7695_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3858_ _7849_/Q _7850_/Q _7851_/Q _7852_/Q vssd1 vssd1 vccd1 vccd1 _7652_/C sky130_fd_sc_hd__or4_2
X_6646_ _7969_/Q _5931_/A _6652_/S vssd1 vssd1 vccd1 vccd1 _6647_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5528_ _5357_/X _7980_/Q _5530_/S vssd1 vssd1 vccd1 vccd1 _5529_/A sky130_fd_sc_hd__mux2_1
X_8316_ _8442_/CLK _8316_/D vssd1 vssd1 vccd1 vccd1 _8316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _5459_/A vssd1 vssd1 vccd1 vccd1 _8011_/D sky130_fd_sc_hd__clkbuf_1
X_8247_ _8247_/CLK _8247_/D vssd1 vssd1 vccd1 vccd1 _8247_/Q sky130_fd_sc_hd__dfxtp_1
X_8178_ _8178_/CLK _8178_/D vssd1 vssd1 vccd1 vccd1 _8178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7080__53 _7082__55/A vssd1 vssd1 vccd1 vccd1 _8234_/CLK sky130_fd_sc_hd__inv_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7010__498 _7012__500/A vssd1 vssd1 vccd1 vccd1 _8179_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7135__98 _7136__99/A vssd1 vssd1 vccd1 vccd1 _8279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7453__25 _7453__25/A vssd1 vssd1 vccd1 vccd1 _8411_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_0_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_4830_ _8185_/Q _4778_/X _4765_/A _8161_/Q _4740_/S vssd1 vssd1 vccd1 vccd1 _4830_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__clkbuf_2
X_4692_ _8197_/Q _7998_/Q _7934_/Q _7894_/Q _4648_/A _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4692_/X sky130_fd_sc_hd__mux4_1
X_7480_ _7479_/B _7479_/C _7197_/A vssd1 vssd1 vccd1 vccd1 _7480_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8510__209 vssd1 vssd1 vccd1 vccd1 _8510__209/HI caravel_irq[0] sky130_fd_sc_hd__conb_1
X_6431_ _7834_/Q _5956_/A _6433_/S vssd1 vssd1 vccd1 vccd1 _6432_/A sky130_fd_sc_hd__mux2_1
X_6362_ _7815_/Q _6401_/A _6192_/X vssd1 vssd1 vccd1 vccd1 _6362_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8101_ _8101_/CLK _8101_/D vssd1 vssd1 vccd1 vccd1 _8101_/Q sky130_fd_sc_hd__dfxtp_1
X_5313_ _8079_/Q _5025_/A _5246_/A _5312_/X _5088_/A vssd1 vssd1 vccd1 vccd1 _5313_/X
+ sky130_fd_sc_hd__a221o_1
X_6293_ _6293_/A vssd1 vssd1 vccd1 vccd1 _6293_/X sky130_fd_sc_hd__clkbuf_2
X_8032_ _8032_/CLK _8032_/D vssd1 vssd1 vccd1 vccd1 _8032_/Q sky130_fd_sc_hd__dfxtp_1
X_6926__433 _6926__433/A vssd1 vssd1 vccd1 vccd1 _8111_/CLK sky130_fd_sc_hd__inv_2
X_5244_ _5336_/B _5240_/X _5243_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__a211o_1
X_5175_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5307_/S sky130_fd_sc_hd__buf_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4126_ _4123_/Y _4607_/C _4911_/B vssd1 vssd1 vccd1 vccd1 _4129_/C sky130_fd_sc_hd__o21ba_1
XFILLER_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A vssd1 vssd1 vccd1 vccd1 _8376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7816_ _8017_/CLK _7816_/D vssd1 vssd1 vccd1 vccd1 _7816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4959_ _8111_/Q _4229_/X _4965_/S vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7747_ _8425_/CLK _7747_/D vssd1 vssd1 vccd1 vccd1 _7747_/Q sky130_fd_sc_hd__dfxtp_1
X_7678_ _7678_/A vssd1 vssd1 vccd1 vccd1 _7678_/X sky130_fd_sc_hd__clkbuf_2
X_6629_ _6629_/A vssd1 vssd1 vccd1 vccd1 _7961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3626_ clkbuf_0__3626_/X vssd1 vssd1 vccd1 vccd1 _7432__7/A sky130_fd_sc_hd__clkbuf_4
X_7396__153 _7396__153/A vssd1 vssd1 vccd1 vccd1 _8364_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _5931_/A _5939_/B vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__or2_1
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ _6228_/C _5866_/B vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__and2_1
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4813_ _4749_/X _7802_/Q _7727_/Q _4753_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4813_/X
+ sky130_fd_sc_hd__a221o_1
X_5793_ _7793_/Q _4362_/A _5795_/S vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__mux2_1
X_7601_ _7604_/A _7604_/B _7601_/C vssd1 vssd1 vccd1 vccd1 _7602_/A sky130_fd_sc_hd__and3_1
X_7532_ _7534_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _8419_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _4416_/X _4610_/X _4743_/X _4682_/X vssd1 vssd1 vccd1 vccd1 _8137_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4675_ _4661_/X _4666_/X _4672_/X _4673_/X _4746_/A vssd1 vssd1 vccd1 vccd1 _4675_/X
+ sky130_fd_sc_hd__o221a_1
X_7463_ _7680_/A _7498_/B _7461_/X _7462_/X vssd1 vssd1 vccd1 vccd1 _7487_/C sky130_fd_sc_hd__o211ai_1
X_7028__512 _7029__513/A vssd1 vssd1 vccd1 vccd1 _8193_/CLK sky130_fd_sc_hd__inv_2
X_6414_ _7829_/Q _6343_/X _6378_/X vssd1 vssd1 vccd1 vccd1 _7829_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6345_ _6768_/A vssd1 vssd1 vccd1 vccd1 _7478_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3057_ clkbuf_0__3057_/X vssd1 vssd1 vccd1 vccd1 _6252__190/A sky130_fd_sc_hd__clkbuf_4
X_8015_ _8015_/CLK _8015_/D vssd1 vssd1 vccd1 vccd1 _8015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5227_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _6975__470/A sky130_fd_sc_hd__clkbuf_4
X_5158_ _3931_/X _5022_/X _5157_/X _5091_/X vssd1 vssd1 vccd1 vccd1 _8083_/D sky130_fd_sc_hd__o211a_1
XFILLER_72_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4109_ _7603_/A _6242_/A _6206_/A vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__a21oi_2
X_5089_ _8086_/Q _5024_/X _5331_/A _5086_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5089_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6672__322/A sky130_fd_sc_hd__clkbuf_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8532__231 vssd1 vssd1 vccd1 vccd1 _8532__231/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7404__160 _7404__160/A vssd1 vssd1 vccd1 vccd1 _8371_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4460_ _4460_/A vssd1 vssd1 vccd1 vccd1 _8206_/D sky130_fd_sc_hd__clkbuf_1
X_4391_ _4391_/A vssd1 vssd1 vccd1 vccd1 _8229_/D sky130_fd_sc_hd__clkbuf_1
X_6130_ _6130_/A vssd1 vssd1 vccd1 vccd1 _7724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6061_ _6061_/A vssd1 vssd1 vccd1 vccd1 _6077_/S sky130_fd_sc_hd__buf_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _4422_/X _8091_/Q _5016_/S vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963_ _6963_/A _8035_/Q _6963_/C vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__and3_1
X_5914_ _5914_/A vssd1 vssd1 vccd1 vccd1 _5914_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6894_ _6419_/A _7649_/B _6293_/X _7613_/C vssd1 vssd1 vccd1 vccd1 _8087_/D sky130_fd_sc_hd__o211a_1
X_5845_ _4150_/X _7727_/Q _5849_/S vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__mux2_1
X_8516__215 vssd1 vssd1 vccd1 vccd1 _8516__215/HI core0Index[2] sky130_fd_sc_hd__conb_1
XFILLER_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5776_ _5776_/A vssd1 vssd1 vccd1 vccd1 _7801_/D sky130_fd_sc_hd__clkbuf_1
X_6260__196 _6263__199/A vssd1 vssd1 vccd1 vccd1 _7788_/CLK sky130_fd_sc_hd__inv_2
X_7347__114 _7348__115/A vssd1 vssd1 vccd1 vccd1 _8325_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7515_ _7504_/A _7490_/Y _7511_/D _7514_/X vssd1 vssd1 vccd1 vccd1 _8414_/D sky130_fd_sc_hd__o211a_1
X_8495_ _8496_/CLK _8495_/D vssd1 vssd1 vccd1 vccd1 _8495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4727_ _8163_/Q _8155_/Q _8117_/Q _8187_/Q _4650_/X _4651_/X vssd1 vssd1 vccd1 vccd1
+ _4727_/X sky130_fd_sc_hd__mux4_2
X_4658_ _4798_/A vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput90 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__buf_4
XFILLER_107_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4589_ _4604_/S vssd1 vssd1 vccd1 vccd1 _4598_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6328_ _6328_/A vssd1 vssd1 vccd1 vccd1 _6369_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6259_/A vssd1 vssd1 vccd1 vccd1 _6259_/X sky130_fd_sc_hd__buf_1
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6939__443 _6941__445/A vssd1 vssd1 vccd1 vccd1 _8122_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3960_ _8409_/Q _3880_/X _3962_/S vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3891_ _3891_/A vssd1 vssd1 vccd1 vccd1 _8467_/D sky130_fd_sc_hd__clkbuf_1
X_5630_ _5630_/A vssd1 vssd1 vccd1 vccd1 _7915_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3391_ clkbuf_0__3391_/X vssd1 vssd1 vccd1 vccd1 _6882__402/A sky130_fd_sc_hd__clkbuf_4
X_5561_ _5561_/A vssd1 vssd1 vccd1 vccd1 _7943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5492_ _5357_/X _7996_/Q _5494_/S vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__mux2_1
X_8280_ _8280_/CLK _8280_/D vssd1 vssd1 vccd1 vccd1 _8280_/Q sky130_fd_sc_hd__dfxtp_1
X_4512_ _4512_/A vssd1 vssd1 vccd1 vccd1 _8184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7300_ _7309_/A _7300_/B vssd1 vssd1 vccd1 vccd1 _8308_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7231_ _7195_/A _7195_/B _7459_/A vssd1 vssd1 vccd1 vccd1 _7231_/Y sky130_fd_sc_hd__a21oi_1
X_4443_ _8211_/Q _4442_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__mux2_1
X_4374_ _4350_/X _8236_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__mux2_1
X_7162_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _7468_/A sky130_fd_sc_hd__inv_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6113_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__and2_1
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6044_ _7740_/Q _6044_/B vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__or2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7995_ _7995_/CLK _7995_/D vssd1 vssd1 vccd1 vccd1 _7995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5828_ _5828_/A vssd1 vssd1 vccd1 vccd1 _7778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3626_ _7430_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3626_/X sky130_fd_sc_hd__clkbuf_16
X_5759_ _7857_/Q _5577_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5760_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8478_ _8478_/CLK _8478_/D vssd1 vssd1 vccd1 vccd1 _8478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7087__59 _7088__60/A vssd1 vssd1 vccd1 vccd1 _8240_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3239_ clkbuf_0__3239_/X vssd1 vssd1 vccd1 vccd1 _6597__305/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6913__424 _6914__425/A vssd1 vssd1 vccd1 vccd1 _8102_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4090_ _4090_/A vssd1 vssd1 vccd1 vccd1 _8362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6920__428 _6922__430/A vssd1 vssd1 vccd1 vccd1 _8106_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _8424_/Q vssd1 vssd1 vccd1 vccd1 _6800_/Y sky130_fd_sc_hd__inv_2
X_7780_ _7780_/CLK _7780_/D vssd1 vssd1 vccd1 vccd1 _7780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4992_ _4992_/A vssd1 vssd1 vccd1 vccd1 _8099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ _8442_/Q vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__clkbuf_4
X_3874_ _8448_/Q vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3443_ clkbuf_0__3443_/X vssd1 vssd1 vccd1 vccd1 _7134__97/A sky130_fd_sc_hd__clkbuf_4
X_5613_ _5574_/X _7922_/Q _5617_/S vssd1 vssd1 vccd1 vccd1 _5614_/A sky130_fd_sc_hd__mux2_1
X_8401_ _8401_/CLK _8401_/D vssd1 vssd1 vccd1 vccd1 _8401_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3374_ clkbuf_0__3374_/X vssd1 vssd1 vccd1 vccd1 _6830__375/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3411_ _6970_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3411_/X sky130_fd_sc_hd__clkbuf_16
X_8332_ _8332_/CLK _8332_/D vssd1 vssd1 vccd1 vccd1 _8332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5544_ _5544_/A vssd1 vssd1 vccd1 vccd1 _7950_/D sky130_fd_sc_hd__clkbuf_1
X_6517__241 _6518__242/A vssd1 vssd1 vccd1 vccd1 _7881_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5475_ _5475_/A vssd1 vssd1 vccd1 vccd1 _8004_/D sky130_fd_sc_hd__clkbuf_1
X_8263_ _8263_/CLK _8263_/D vssd1 vssd1 vccd1 vccd1 _8263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8194_ _8194_/CLK _8194_/D vssd1 vssd1 vccd1 vccd1 _8194_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3273_ _6670_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3273_/X sky130_fd_sc_hd__clkbuf_16
X_4426_ _4425_/X _8216_/Q _4429_/S vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__mux2_1
X_7214_ _8494_/Q _7241_/A _7241_/B vssd1 vssd1 vccd1 vccd1 _7214_/X sky130_fd_sc_hd__and3_1
X_7145_ _7600_/A _6242_/X _6157_/A vssd1 vssd1 vccd1 vccd1 _7345_/S sky130_fd_sc_hd__a21oi_4
X_4357_ _4356_/X _8242_/Q _4357_/S vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7107_/A vssd1 vssd1 vccd1 vccd1 _7076_/X sky130_fd_sc_hd__buf_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4288_ _4515_/A _4343_/B vssd1 vssd1 vccd1 vccd1 _4304_/S sky130_fd_sc_hd__or2_4
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _7811_/Q input28/X _6039_/S vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7978_ _7978_/CLK _7978_/D vssd1 vssd1 vccd1 vccd1 _7978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6942_/A vssd1 vssd1 vccd1 vccd1 _6929_/X sky130_fd_sc_hd__buf_1
XFILLER_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8447_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_70 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7622__31 _7624__33/A vssd1 vssd1 vccd1 vccd1 _8454_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_92 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_81 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _5224_/A _5258_/X _5259_/X vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6139__180 _6139__180/A vssd1 vssd1 vccd1 vccd1 _7729_/CLK sky130_fd_sc_hd__inv_2
X_4211_ _8330_/Q _4141_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__mux2_1
X_5191_ _8400_/Q _5046_/B _5190_/X _5305_/A vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__o22a_1
X_7022__507 _7024__509/A vssd1 vssd1 vccd1 vccd1 _8188_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ _8354_/Q _4141_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4143_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4073_ _3931_/X _8369_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__mux2_1
X_7901_ _7901_/CLK _7901_/D vssd1 vssd1 vccd1 vccd1 _7901_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_opt_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7832_ _8497_/CLK _7832_/D vssd1 vssd1 vccd1 vccd1 _7832_/Q sky130_fd_sc_hd__dfxtp_2
X_4975_ _4997_/S vssd1 vssd1 vccd1 vccd1 _4988_/S sky130_fd_sc_hd__buf_2
X_7763_ _8433_/CLK _7763_/D vssd1 vssd1 vccd1 vccd1 _7763_/Q sky130_fd_sc_hd__dfxtp_1
X_3926_ _3925_/X _8456_/Q _3935_/S vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__mux2_1
X_6714_ _6410_/C _6624_/A _6714_/S vssd1 vssd1 vccd1 vccd1 _6715_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3426_ clkbuf_0__3426_/X vssd1 vssd1 vccd1 vccd1 _7050__530/A sky130_fd_sc_hd__clkbuf_4
X_7694_ _7692_/Y _7693_/Y _7678_/X vssd1 vssd1 vccd1 vccd1 _8489_/D sky130_fd_sc_hd__a21oi_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6645_ _6645_/A vssd1 vssd1 vccd1 vccd1 _7968_/D sky130_fd_sc_hd__clkbuf_1
X_3857_ _7845_/Q _7846_/Q _7847_/Q _7848_/Q vssd1 vssd1 vccd1 vccd1 _7652_/B sky130_fd_sc_hd__or4_1
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5527_ _5527_/A vssd1 vssd1 vccd1 vccd1 _7981_/D sky130_fd_sc_hd__clkbuf_1
X_8315_ _8315_/CLK _8315_/D vssd1 vssd1 vccd1 vccd1 _8315_/Q sky130_fd_sc_hd__dfxtp_1
X_8246_ _8246_/CLK _8246_/D vssd1 vssd1 vccd1 vccd1 _8246_/Q sky130_fd_sc_hd__dfxtp_1
X_5458_ _8011_/Q _4445_/X _5458_/S vssd1 vssd1 vccd1 vccd1 _5459_/A sky130_fd_sc_hd__mux2_1
X_5389_ _5389_/A vssd1 vssd1 vccd1 vccd1 _8046_/D sky130_fd_sc_hd__clkbuf_1
X_8177_ _8177_/CLK _8177_/D vssd1 vssd1 vccd1 vccd1 _8177_/Q sky130_fd_sc_hd__dfxtp_1
X_4409_ _4409_/A vssd1 vssd1 vccd1 vccd1 _8222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7438__12 _7439__13/A vssd1 vssd1 vccd1 vccd1 _8398_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6878__400 _6878__400/A vssd1 vssd1 vccd1 vccd1 _8076_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4789_/A vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4691_ _4637_/X _4688_/X _4690_/X vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__a21o_1
X_6430_ _6430_/A vssd1 vssd1 vccd1 vccd1 _7833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6361_ _6359_/X _6293_/X _6371_/A _6355_/X _6360_/X vssd1 vssd1 vccd1 vccd1 _6361_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8100_ _8100_/CLK _8100_/D vssd1 vssd1 vccd1 vccd1 _8100_/Q sky130_fd_sc_hd__dfxtp_1
X_5312_ _5031_/A _5290_/X _5297_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6292_ _8016_/Q _6292_/B vssd1 vssd1 vccd1 vccd1 _6293_/A sky130_fd_sc_hd__and2_1
XFILLER_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8031_ _8031_/CLK _8031_/D vssd1 vssd1 vccd1 vccd1 _8031_/Q sky130_fd_sc_hd__dfxtp_1
X_5243_ _5220_/X _5241_/X _5242_/X vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5174_ _5305_/A vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__buf_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _8130_/Q _4653_/A vssd1 vssd1 vccd1 vccd1 _4607_/C sky130_fd_sc_hd__xor2_1
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4056_ _8376_/Q _4010_/X _4056_/S vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7815_ _8017_/CLK _7815_/D vssd1 vssd1 vccd1 vccd1 _7815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4958_ _4958_/A vssd1 vssd1 vccd1 vccd1 _8112_/D sky130_fd_sc_hd__clkbuf_1
X_7746_ _8489_/CLK _7746_/D vssd1 vssd1 vccd1 vccd1 _7746_/Q sky130_fd_sc_hd__dfxtp_1
X_3909_ _3909_/A vssd1 vssd1 vccd1 vccd1 _8461_/D sky130_fd_sc_hd__clkbuf_1
X_4889_ _4932_/B _4887_/X _4888_/X vssd1 vssd1 vccd1 vccd1 _4889_/X sky130_fd_sc_hd__o21a_1
X_7677_ _7677_/A _7693_/B vssd1 vssd1 vccd1 vccd1 _7677_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__3409_ clkbuf_0__3409_/X vssd1 vssd1 vccd1 vccd1 _6969__465/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6628_ _5913_/A _7961_/Q _6634_/S vssd1 vssd1 vccd1 vccd1 _6629_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6559_ _6559_/A vssd1 vssd1 vccd1 vccd1 _6559_/X sky130_fd_sc_hd__buf_1
X_8229_ _8229_/CLK _8229_/D vssd1 vssd1 vccd1 vccd1 _8229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3239_ _6592_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3239_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3625_ clkbuf_0__3625_/X vssd1 vssd1 vccd1 vccd1 _7429__5/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6496__225 _6496__225/A vssd1 vssd1 vccd1 vccd1 _7865_/CLK sky130_fd_sc_hd__inv_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5939_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _5861_/A vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7600_ _7600_/A _7675_/B vssd1 vssd1 vccd1 vccd1 _7601_/C sky130_fd_sc_hd__and2_1
X_5792_ _5792_/A vssd1 vssd1 vccd1 vccd1 _7794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4812_ _4419_/X _4610_/X _4811_/X _4682_/X vssd1 vssd1 vccd1 vccd1 _8136_/D sky130_fd_sc_hd__o211a_1
X_7531_ _8419_/Q _7530_/X _7527_/X _7478_/B vssd1 vssd1 vccd1 vccd1 _7532_/B sky130_fd_sc_hd__o2bb2a_1
X_4743_ _4612_/X _8137_/Q _4924_/A _4742_/X _4678_/X vssd1 vssd1 vccd1 vccd1 _4743_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7462_ _7692_/A _7462_/B vssd1 vssd1 vccd1 vccd1 _7462_/X sky130_fd_sc_hd__xor2_1
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4674_ _8126_/Q _4674_/B vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__xnor2_4
X_6413_ _7828_/Q _6401_/X _6371_/A _6412_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _7828_/D
+ sky130_fd_sc_hd__a221o_1
X_7393_ _7417_/A vssd1 vssd1 vccd1 vccd1 _7393_/X sky130_fd_sc_hd__buf_1
X_6344_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _6768_/A sky130_fd_sc_hd__buf_2
XFILLER_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8014_ _8014_/CLK _8014_/D vssd1 vssd1 vccd1 vccd1 _8014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6666__317 _6667__318/A vssd1 vssd1 vccd1 vccd1 _7981_/CLK sky130_fd_sc_hd__inv_2
X_5226_ _8201_/Q _8209_/Q _5241_/S vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5157_ _8083_/Q _5024_/X _5246_/A _5156_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5157_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4108_ _5853_/B _7659_/A _7659_/B _4108_/D vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__and4_1
X_5088_ _5088_/A vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6669__320/A sky130_fd_sc_hd__clkbuf_4
X_4039_ _8383_/Q _4014_/X _4043_/S vssd1 vssd1 vccd1 vccd1 _4040_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7729_ _7729_/CLK _7729_/D vssd1 vssd1 vccd1 vccd1 _7729_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7113__80 _7113__80/A vssd1 vssd1 vccd1 vccd1 _8261_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _4347_/X _8229_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4391_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6511__236 _6514__239/A vssd1 vssd1 vccd1 vccd1 _7876_/CLK sky130_fd_sc_hd__inv_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6060_ _6053_/X _6058_/X _6059_/X _6056_/X vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__o211a_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _8092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _5913_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__or2_4
X_6893_ _7615_/C vssd1 vssd1 vccd1 vccd1 _7613_/C sky130_fd_sc_hd__clkbuf_2
X_5844_ _5844_/A vssd1 vssd1 vccd1 vccd1 _7728_/D sky130_fd_sc_hd__clkbuf_1
X_5775_ _4153_/X _7801_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__mux2_1
X_7514_ _7582_/A vssd1 vssd1 vccd1 vccd1 _7514_/X sky130_fd_sc_hd__buf_2
X_4726_ _8329_/Q _8219_/Q _7876_/Q _8353_/Q _4648_/X _4633_/X vssd1 vssd1 vccd1 vccd1
+ _4726_/X sky130_fd_sc_hd__mux4_1
X_8494_ _8498_/CLK _8494_/D vssd1 vssd1 vccd1 vccd1 _8494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4657_ _4637_/X _4649_/X _4656_/X vssd1 vssd1 vccd1 vccd1 _4657_/X sky130_fd_sc_hd__a21o_1
Xinput80 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__clkbuf_2
Xinput91 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _5939_/A sky130_fd_sc_hd__buf_4
X_4588_ _4588_/A _5430_/B vssd1 vssd1 vccd1 vccd1 _4604_/S sky130_fd_sc_hd__nor2_2
X_6327_ _8475_/Q _6311_/X _6326_/X _6306_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _6327_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5209_ _5224_/A vssd1 vssd1 vccd1 vccd1 _5338_/B sky130_fd_sc_hd__clkbuf_2
X_6189_ _6184_/X _7964_/Q _6186_/X _6188_/X _7753_/Q vssd1 vssd1 vccd1 vccd1 _7753_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7629__37 _7629__37/A vssd1 vssd1 vccd1 vccd1 _8460_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8539__238 vssd1 vssd1 vccd1 vccd1 _8539__238/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _8467_/Q _3889_/X _3893_/S vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3390_ clkbuf_0__3390_/X vssd1 vssd1 vccd1 vccd1 _6909_/A sky130_fd_sc_hd__clkbuf_4
X_5560_ _5557_/X _7943_/Q _5572_/S vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__mux2_1
X_5491_ _5491_/A vssd1 vssd1 vccd1 vccd1 _7997_/D sky130_fd_sc_hd__clkbuf_1
X_4511_ _8184_/Q _4244_/X _4513_/S vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__mux2_1
X_4442_ _8446_/Q vssd1 vssd1 vccd1 vccd1 _4442_/X sky130_fd_sc_hd__buf_2
X_7230_ _8288_/Q vssd1 vssd1 vccd1 vccd1 _7320_/B sky130_fd_sc_hd__inv_2
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4373_ _4373_/A vssd1 vssd1 vccd1 vccd1 _8237_/D sky130_fd_sc_hd__clkbuf_1
X_7161_ _7161_/A _7236_/C _7161_/C vssd1 vssd1 vccd1 vccd1 _7222_/B sky130_fd_sc_hd__and3_1
XFILLER_112_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6112_/A vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _7815_/Q input32/X _6058_/S vssd1 vssd1 vccd1 vccd1 _6043_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7994_ _7994_/CLK _7994_/D vssd1 vssd1 vccd1 vccd1 _7994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7071__547 _7073__549/A vssd1 vssd1 vccd1 vccd1 _8228_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5827_ _7778_/Q _5574_/A _5831_/S vssd1 vssd1 vccd1 vccd1 _5828_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3625_ _7424_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3625_/X sky130_fd_sc_hd__clkbuf_16
X_5758_ _5758_/A vssd1 vssd1 vccd1 vccd1 _7858_/D sky130_fd_sc_hd__clkbuf_1
X_4709_ _8049_/Q _8041_/Q _7869_/Q _8110_/Q _4648_/X _4640_/X vssd1 vssd1 vccd1 vccd1
+ _4709_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8477_ _8478_/CLK _8477_/D vssd1 vssd1 vccd1 vccd1 _8477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5689_ _7888_/Q _4996_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679__327 _6682__330/A vssd1 vssd1 vccd1 vccd1 _7991_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3238_ clkbuf_0__3238_/X vssd1 vssd1 vccd1 vccd1 _6670_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _8099_/Q _4990_/X _4997_/S vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _3942_/A vssd1 vssd1 vccd1 vccd1 _8451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3873_ _3873_/A vssd1 vssd1 vccd1 vccd1 _8473_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3442_ clkbuf_0__3442_/X vssd1 vssd1 vccd1 vccd1 _7131__95/A sky130_fd_sc_hd__clkbuf_4
X_5612_ _5612_/A vssd1 vssd1 vccd1 vccd1 _7923_/D sky130_fd_sc_hd__clkbuf_1
X_6592_ _6598_/A vssd1 vssd1 vccd1 vccd1 _6592_/X sky130_fd_sc_hd__buf_1
X_8400_ _8400_/CLK _8400_/D vssd1 vssd1 vccd1 vccd1 _8400_/Q sky130_fd_sc_hd__dfxtp_1
X_5543_ _7950_/Q _4978_/X _5549_/S vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__mux2_1
X_8331_ _8331_/CLK _8331_/D vssd1 vssd1 vccd1 vccd1 _8331_/Q sky130_fd_sc_hd__dfxtp_1
X_8262_ _8262_/CLK _8262_/D vssd1 vssd1 vccd1 vccd1 _8262_/Q sky130_fd_sc_hd__dfxtp_1
X_5474_ _8004_/Q _4353_/A _5476_/S vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__mux2_1
X_8193_ _8193_/CLK _8193_/D vssd1 vssd1 vccd1 vccd1 _8193_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3272_ _6664_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3272_/X sky130_fd_sc_hd__clkbuf_16
X_7213_ _7241_/A _7241_/B _6768_/A vssd1 vssd1 vccd1 vccd1 _7213_/Y sky130_fd_sc_hd__a21oi_1
X_4425_ _8061_/Q vssd1 vssd1 vccd1 vccd1 _4425_/X sky130_fd_sc_hd__buf_2
X_4356_ _4356_/A vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7075_ _7075_/A vssd1 vssd1 vccd1 vccd1 _7075_/X sky130_fd_sc_hd__buf_1
X_4287_ _4287_/A _4287_/B _3972_/B vssd1 vssd1 vccd1 vccd1 _4343_/B sky130_fd_sc_hd__or3b_4
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6026_ _6009_/X _6024_/X _6025_/X _6018_/X vssd1 vssd1 vccd1 vccd1 _6026_/X sky130_fd_sc_hd__o211a_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092__63 _7092__63/A vssd1 vssd1 vccd1 vccd1 _8244_/CLK sky130_fd_sc_hd__inv_2
X_7390__149 _7391__150/A vssd1 vssd1 vccd1 vccd1 _8360_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _7977_/CLK _7977_/D vssd1 vssd1 vccd1 vccd1 _7977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6859_ _8437_/Q _6863_/B vssd1 vssd1 vccd1 vccd1 _6860_/A sky130_fd_sc_hd__and2_1
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_71 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_60 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_93 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_82 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6579__291 _6580__292/A vssd1 vssd1 vccd1 vccd1 _7931_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _4210_/A vssd1 vssd1 vccd1 vccd1 _8331_/D sky130_fd_sc_hd__clkbuf_1
X_5190_ _7787_/Q _8384_/Q _5190_/S vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4141_ _8065_/Q vssd1 vssd1 vccd1 vccd1 _4141_/X sky130_fd_sc_hd__buf_2
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _4072_/A vssd1 vssd1 vccd1 vccd1 _8370_/D sky130_fd_sc_hd__clkbuf_1
X_7900_ _7900_/CLK _7900_/D vssd1 vssd1 vccd1 vccd1 _7900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7831_ _8499_/CLK _7831_/D vssd1 vssd1 vccd1 vccd1 _7831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _5815_/A _5558_/A vssd1 vssd1 vccd1 vccd1 _4997_/S sky130_fd_sc_hd__nor2_2
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7762_ _8433_/CLK _7762_/D vssd1 vssd1 vccd1 vccd1 _7762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3925_ _8448_/Q vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__buf_4
X_7693_ _7693_/A _7693_/B vssd1 vssd1 vccd1 vccd1 _7693_/Y sky130_fd_sc_hd__nand2_1
X_6713_ _6713_/A vssd1 vssd1 vccd1 vccd1 _8017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3425_ clkbuf_0__3425_/X vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__clkbuf_4
X_6644_ _7968_/Q _5928_/A _6652_/S vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__mux2_1
X_3856_ _7854_/Q _7853_/Q vssd1 vssd1 vccd1 vccd1 _7652_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3287_ clkbuf_0__3287_/X vssd1 vssd1 vccd1 vccd1 _6734__367/A sky130_fd_sc_hd__clkbuf_4
X_5526_ _5353_/X _7981_/Q _5530_/S vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__mux2_1
X_8314_ _8315_/CLK _8314_/D vssd1 vssd1 vccd1 vccd1 _8314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8245_ _8245_/CLK _8245_/D vssd1 vssd1 vccd1 vccd1 _8245_/Q sky130_fd_sc_hd__dfxtp_1
X_5457_ _5457_/A vssd1 vssd1 vccd1 vccd1 _8012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4408_ _4404_/X _8222_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__mux2_1
X_5388_ _5365_/X _8046_/Q _5392_/S vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__mux2_1
X_8176_ _8176_/CLK _8176_/D vssd1 vssd1 vccd1 vccd1 _8176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4339_ _4339_/A vssd1 vssd1 vccd1 vccd1 _8248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4627_/A _4689_/X _4721_/A vssd1 vssd1 vccd1 vccd1 _4690_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6360_ _8140_/Q _6318_/X _6353_/X vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__a21o_1
X_5311_ _5278_/A _5300_/X _5303_/X _5310_/X _5332_/B vssd1 vssd1 vccd1 vccd1 _5311_/X
+ sky130_fd_sc_hd__o311a_1
X_6885__405 _6885__405/A vssd1 vssd1 vccd1 vccd1 _8081_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8030_ _8030_/CLK _8030_/D vssd1 vssd1 vccd1 vccd1 _8030_/Q sky130_fd_sc_hd__dfxtp_1
X_6291_ _6291_/A vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__clkbuf_2
X_5242_ _8367_/Q _5214_/A _5239_/B _8359_/Q _5074_/X vssd1 vssd1 vccd1 vccd1 _5242_/X
+ sky130_fd_sc_hd__o221a_1
X_5173_ _8234_/Q _5163_/X _5295_/A _5169_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _5173_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _8125_/Q vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__clkbuf_4
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_4055_ _4055_/A vssd1 vssd1 vccd1 vccd1 _8377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7814_ _8481_/CLK _7814_/D vssd1 vssd1 vccd1 vccd1 _7814_/Q sky130_fd_sc_hd__dfxtp_1
X_4957_ _8112_/Q _4223_/X _4965_/S vssd1 vssd1 vccd1 vccd1 _4958_/A sky130_fd_sc_hd__mux2_1
X_7745_ _8489_/CLK _7745_/D vssd1 vssd1 vccd1 vccd1 _7745_/Q sky130_fd_sc_hd__dfxtp_1
X_6933__439 _6934__440/A vssd1 vssd1 vccd1 vccd1 _8117_/CLK sky130_fd_sc_hd__inv_2
X_3908_ _8461_/Q _3883_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3909_/A sky130_fd_sc_hd__mux2_1
X_4888_ _8349_/Q _4619_/A _4803_/X _8325_/Q _4798_/X vssd1 vssd1 vccd1 vccd1 _4888_/X
+ sky130_fd_sc_hd__o221a_1
X_7676_ _7699_/B vssd1 vssd1 vccd1 vccd1 _7693_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6627_ _6627_/A vssd1 vssd1 vccd1 vccd1 _7960_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3408_ clkbuf_0__3408_/X vssd1 vssd1 vccd1 vccd1 _6960__460/A sky130_fd_sc_hd__clkbuf_4
X_3839_ _8087_/Q _3918_/A vssd1 vssd1 vccd1 vccd1 _5328_/B sky130_fd_sc_hd__and2_1
XFILLER_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5509_ _5509_/A vssd1 vssd1 vccd1 vccd1 _7989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8228_ _8228_/CLK _8228_/D vssd1 vssd1 vccd1 vccd1 _8228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3238_ _6591_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3238_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3624_ clkbuf_0__3624_/X vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__clkbuf_4
X_8159_ _8159_/CLK _8159_/D vssd1 vssd1 vccd1 vccd1 _8159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5860_ _6423_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__and2_1
XFILLER_46_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4612_/X _8136_/Q _4925_/A _4810_/X _4678_/X vssd1 vssd1 vccd1 vccd1 _4811_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5791_ _7794_/Q _4359_/A _5795_/S vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__mux2_1
X_4742_ _4622_/X _4729_/X _4733_/X _4741_/X vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__a31o_1
X_7530_ _7557_/B vssd1 vssd1 vccd1 vccd1 _7530_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4721_/A vssd1 vssd1 vccd1 vccd1 _4673_/X sky130_fd_sc_hd__clkbuf_2
X_7461_ _7689_/A _7461_/B vssd1 vssd1 vccd1 vccd1 _7461_/X sky130_fd_sc_hd__xor2_1
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6412_ _8479_/Q _6412_/B _8018_/Q vssd1 vssd1 vccd1 vccd1 _6412_/X sky130_fd_sc_hd__and3_1
X_7392_ _7392_/A vssd1 vssd1 vccd1 vccd1 _7392_/X sky130_fd_sc_hd__buf_1
X_6343_ _6343_/A vssd1 vssd1 vccd1 vccd1 _6343_/X sky130_fd_sc_hd__buf_2
XFILLER_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8013_ _8013_/CLK _8013_/D vssd1 vssd1 vccd1 vccd1 _8013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5225_ _8177_/Q _5214_/X _5216_/X _8169_/Q _5099_/X vssd1 vssd1 vccd1 vccd1 _5225_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5031_/X _5143_/X _5147_/X _5155_/X vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__a31o_2
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _5087_/A _7323_/A vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__and2_1
X_4107_ _8127_/Q vssd1 vssd1 vccd1 vccd1 _4903_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4038_ _4038_/A vssd1 vssd1 vccd1 vccd1 _8384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7035__518 _7037__520/A vssd1 vssd1 vccd1 vccd1 _8199_/CLK sky130_fd_sc_hd__inv_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5989_ _7964_/Q _5993_/B vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__and2_2
X_7728_ _7728_/CLK _7728_/D vssd1 vssd1 vccd1 vccd1 _7728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659_ _7659_/A _7659_/B _7659_/C vssd1 vssd1 vccd1 vccd1 _7704_/B sky130_fd_sc_hd__and3_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput190 _6100_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4419_/X _8092_/Q _5010_/S vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6961_ _6976_/A vssd1 vssd1 vccd1 vccd1 _6961_/X sky130_fd_sc_hd__buf_1
X_5912_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6892_ _6892_/A _7604_/B vssd1 vssd1 vccd1 vccd1 _7615_/C sky130_fd_sc_hd__and2_1
X_5843_ _4147_/X _7728_/Q _5843_/S vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5774_ _5774_/A vssd1 vssd1 vccd1 vccd1 _7802_/D sky130_fd_sc_hd__clkbuf_1
X_7427__3 _7429__5/A vssd1 vssd1 vccd1 vccd1 _8389_/CLK sky130_fd_sc_hd__inv_2
X_6672__322 _6672__322/A vssd1 vssd1 vccd1 vccd1 _7986_/CLK sky130_fd_sc_hd__inv_2
X_7513_ _7575_/A vssd1 vssd1 vccd1 vccd1 _7582_/A sky130_fd_sc_hd__clkbuf_2
X_8493_ _8498_/CLK _8493_/D vssd1 vssd1 vccd1 vccd1 _8493_/Q sky130_fd_sc_hd__dfxtp_1
X_4725_ _4413_/X _4610_/X _4724_/X _4682_/X vssd1 vssd1 vccd1 vccd1 _8138_/D sky130_fd_sc_hd__o211a_1
XFILLER_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4656_ _4627_/A _4652_/X _4883_/A vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__a21o_1
X_4587_ _4587_/A vssd1 vssd1 vccd1 vccd1 _8151_/D sky130_fd_sc_hd__clkbuf_1
Xinput81 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _7600_/A sky130_fd_sc_hd__buf_6
Xinput70 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _7597_/A sky130_fd_sc_hd__buf_8
XFILLER_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput92 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _7603_/A sky130_fd_sc_hd__buf_6
X_6326_ _8135_/Q _6318_/X _6319_/X vssd1 vssd1 vccd1 vccd1 _6326_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7099__69 _7100__70/A vssd1 vssd1 vccd1 vccd1 _8250_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5220_/A vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__buf_2
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6188_/X sky130_fd_sc_hd__clkbuf_2
X_5139_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6978__472 _6979__473/A vssd1 vssd1 vccd1 vccd1 _8153_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6573__286 _6574__287/A vssd1 vssd1 vccd1 vccd1 _7926_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6946__449 _6947__450/A vssd1 vssd1 vccd1 vccd1 _8128_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5490_ _5353_/X _7997_/Q _5494_/S vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__mux2_1
X_4510_ _4510_/A vssd1 vssd1 vccd1 vccd1 _8185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4441_ _4441_/A vssd1 vssd1 vccd1 vccd1 _8212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7160_ _8485_/Q _7305_/A _7305_/B vssd1 vssd1 vccd1 vccd1 _7161_/C sky130_fd_sc_hd__nand3b_1
X_4372_ _4347_/X _8237_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__clkbuf_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6061_/A vssd1 vssd1 vccd1 vccd1 _6058_/S sky130_fd_sc_hd__buf_2
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8522__221 vssd1 vssd1 vccd1 vccd1 _8522__221/HI core1Index[1] sky130_fd_sc_hd__conb_1
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7993_ _7993_/CLK _7993_/D vssd1 vssd1 vccd1 vccd1 _7993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5826_ _5826_/A vssd1 vssd1 vccd1 vccd1 _7779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3624_ _7423_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3624_/X sky130_fd_sc_hd__clkbuf_16
X_5757_ _7858_/Q _5574_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__mux2_1
X_4708_ _4930_/B _4705_/X _4707_/X vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__a21o_1
X_8476_ _8497_/CLK _8476_/D vssd1 vssd1 vccd1 vccd1 _8476_/Q sky130_fd_sc_hd__dfxtp_1
X_5688_ _5688_/A vssd1 vssd1 vccd1 vccd1 _7889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4639_ _4670_/A vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7289_ _7289_/A _7289_/B vssd1 vssd1 vccd1 vccd1 _7289_/Y sky130_fd_sc_hd__nand2_1
X_6309_ _8133_/Q _6318_/A _6353_/A vssd1 vssd1 vccd1 vccd1 _6309_/X sky130_fd_sc_hd__a21o_1
X_7634__41 _7635__42/A vssd1 vssd1 vccd1 vccd1 _8464_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3237_ clkbuf_0__3237_/X vssd1 vssd1 vccd1 vccd1 _6879_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952__453 _6952__453/A vssd1 vssd1 vccd1 vccd1 _8132_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7048__528 _7048__528/A vssd1 vssd1 vccd1 vccd1 _8209_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4990_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _4990_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3441_ clkbuf_0__3441_/X vssd1 vssd1 vccd1 vccd1 _7123__88/A sky130_fd_sc_hd__clkbuf_4
X_3941_ _3940_/X _8451_/Q _3944_/S vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3872_ _8473_/Q _3812_/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5611_ _5571_/X _7923_/Q _5611_/S vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__mux2_1
X_6591_ _6879_/A vssd1 vssd1 vccd1 vccd1 _6591_/X sky130_fd_sc_hd__buf_1
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5542_ _5542_/A vssd1 vssd1 vccd1 vccd1 _7951_/D sky130_fd_sc_hd__clkbuf_1
X_8330_ _8330_/CLK _8330_/D vssd1 vssd1 vccd1 vccd1 _8330_/Q sky130_fd_sc_hd__dfxtp_1
X_8261_ _8261_/CLK _8261_/D vssd1 vssd1 vccd1 vccd1 _8261_/Q sky130_fd_sc_hd__dfxtp_1
X_5473_ _5473_/A vssd1 vssd1 vccd1 vccd1 _8005_/D sky130_fd_sc_hd__clkbuf_1
X_8192_ _8192_/CLK _8192_/D vssd1 vssd1 vccd1 vccd1 _8192_/Q sky130_fd_sc_hd__dfxtp_1
X_7212_ _8301_/Q _7211_/C _8302_/Q vssd1 vssd1 vccd1 vccd1 _7241_/B sky130_fd_sc_hd__a21o_1
X_4424_ _4424_/A vssd1 vssd1 vccd1 vccd1 _8217_/D sky130_fd_sc_hd__clkbuf_1
X_4355_ _4355_/A vssd1 vssd1 vccd1 vccd1 _8243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4286_/A vssd1 vssd1 vccd1 vccd1 _8271_/D sky130_fd_sc_hd__clkbuf_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6025_ _7735_/Q _6025_/B vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__or2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6524__247 _6524__247/A vssd1 vssd1 vccd1 vccd1 _7887_/CLK sky130_fd_sc_hd__inv_2
X_7976_ _7976_/CLK _7976_/D vssd1 vssd1 vccd1 vccd1 _7976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6858_ _6858_/A vssd1 vssd1 vccd1 vccd1 _8062_/D sky130_fd_sc_hd__clkbuf_1
X_5809_ _3886_/X _7786_/Q _5813_/S vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6789_ _6789_/A _6789_/B _6789_/C vssd1 vssd1 vccd1 vccd1 _7468_/B sky130_fd_sc_hd__nand3_2
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8459_ _8459_/CLK _8459_/D vssd1 vssd1 vccd1 vccd1 _8459_/Q sky130_fd_sc_hd__dfxtp_1
X_6685__332 _6685__332/A vssd1 vssd1 vccd1 vccd1 _7996_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_61 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_50 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_83 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_72 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_94 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6733__366 _6734__367/A vssd1 vssd1 vccd1 vccd1 _8033_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4140_ _4140_/A vssd1 vssd1 vccd1 vccd1 _8355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4071_ _3928_/X _8370_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7830_ _8017_/CLK _7830_/D vssd1 vssd1 vccd1 vccd1 _7830_/Q sky130_fd_sc_hd__dfxtp_1
X_6959__459 _6960__460/A vssd1 vssd1 vccd1 vccd1 _8138_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4973_ _8067_/Q vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__clkbuf_4
X_7761_ _8441_/CLK _7761_/D vssd1 vssd1 vccd1 vccd1 _7761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3924_ _3924_/A vssd1 vssd1 vccd1 vccd1 _8457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7692_ _7692_/A _7692_/B vssd1 vssd1 vccd1 vccd1 _7692_/Y sky130_fd_sc_hd__nand2_1
X_6712_ _6387_/C _6606_/A _6714_/S vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3424_ clkbuf_0__3424_/X vssd1 vssd1 vccd1 vccd1 _7043__525/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6643_ _6658_/S vssd1 vssd1 vccd1 vccd1 _6652_/S sky130_fd_sc_hd__buf_2
X_3855_ _7654_/A _6287_/A vssd1 vssd1 vccd1 vccd1 _7659_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3286_ clkbuf_0__3286_/X vssd1 vssd1 vccd1 vccd1 _6731__365/A sky130_fd_sc_hd__clkbuf_4
X_5525_ _5525_/A vssd1 vssd1 vccd1 vccd1 _7982_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_22_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8489_/CLK sky130_fd_sc_hd__clkbuf_16
X_8313_ _8315_/CLK _8313_/D vssd1 vssd1 vccd1 vccd1 _8313_/Q sky130_fd_sc_hd__dfxtp_1
X_8244_ _8244_/CLK _8244_/D vssd1 vssd1 vccd1 vccd1 _8244_/Q sky130_fd_sc_hd__dfxtp_1
X_5456_ _8012_/Q _4442_/X _5458_/S vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4407_ _4429_/S vssd1 vssd1 vccd1 vccd1 _4420_/S sky130_fd_sc_hd__buf_2
X_6530__251 _6531__252/A vssd1 vssd1 vccd1 vccd1 _7891_/CLK sky130_fd_sc_hd__inv_2
X_5387_ _5387_/A vssd1 vssd1 vccd1 vccd1 _8047_/D sky130_fd_sc_hd__clkbuf_1
X_8175_ _8175_/CLK _8175_/D vssd1 vssd1 vccd1 vccd1 _8175_/Q sky130_fd_sc_hd__dfxtp_1
X_7126_ _7132_/A vssd1 vssd1 vccd1 vccd1 _7126_/X sky130_fd_sc_hd__buf_1
X_4338_ _8248_/Q _4197_/X _4340_/S vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _5502_/B _5448_/B vssd1 vssd1 vccd1 vccd1 _4285_/S sky130_fd_sc_hd__nor2_4
X_7057_ _7057_/A vssd1 vssd1 vccd1 vccd1 _7057_/X sky130_fd_sc_hd__buf_1
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _6008_/A vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7959_ _8425_/CLK _7959_/D vssd1 vssd1 vccd1 vccd1 _7959_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5310_ _5305_/X _5306_/X _5113_/X _5309_/X vssd1 vssd1 vccd1 vccd1 _5310_/X sky130_fd_sc_hd__a211o_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6290_ _8499_/Q vssd1 vssd1 vccd1 vccd1 _7207_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5241_ _8335_/Q _8343_/Q _5241_/S vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__mux2_1
X_5172_ _8469_/Q _5285_/B vssd1 vssd1 vccd1 vccd1 _5172_/X sky130_fd_sc_hd__or2_1
XFILLER_68_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7444__17 _7445__18/A vssd1 vssd1 vccd1 vccd1 _8403_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4123_ _8128_/Q _8127_/Q _4113_/B vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__a21oi_1
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ _8377_/Q _4006_/X _4056_/S vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7813_ _8017_/CLK _7813_/D vssd1 vssd1 vccd1 vccd1 _7813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7744_ _8490_/CLK _7744_/D vssd1 vssd1 vccd1 vccd1 _7744_/Q sky130_fd_sc_hd__dfxtp_1
X_6972__467 _6973__468/A vssd1 vssd1 vccd1 vccd1 _8148_/CLK sky130_fd_sc_hd__inv_2
X_4956_ _4971_/S vssd1 vssd1 vccd1 vccd1 _4965_/S sky130_fd_sc_hd__buf_2
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _8462_/D sky130_fd_sc_hd__clkbuf_1
X_4887_ _8215_/Q _4801_/X _4787_/X _7872_/Q vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__a22o_1
X_7675_ _8017_/Q _7675_/B _7701_/B vssd1 vssd1 vccd1 vccd1 _7699_/B sky130_fd_sc_hd__and3_1
X_6626_ _5911_/A _7960_/Q _6634_/S vssd1 vssd1 vccd1 vccd1 _6627_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3407_ clkbuf_0__3407_/X vssd1 vssd1 vccd1 vccd1 _6954__455/A sky130_fd_sc_hd__clkbuf_4
X_3838_ _3838_/A _3838_/B _3838_/C _3838_/D vssd1 vssd1 vccd1 vccd1 _3918_/A sky130_fd_sc_hd__or4_1
X_5508_ _7989_/Q _4350_/A _5512_/S vssd1 vssd1 vccd1 vccd1 _5509_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8227_ _8227_/CLK _8227_/D vssd1 vssd1 vccd1 vccd1 _8227_/Q sky130_fd_sc_hd__dfxtp_1
X_5439_ _5439_/A vssd1 vssd1 vccd1 vccd1 _8023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7125__90 _7125__90/A vssd1 vssd1 vccd1 vccd1 _8271_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3237_ _6590_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3237_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3623_ clkbuf_0__3623_/X vssd1 vssd1 vccd1 vccd1 _7419__172/A sky130_fd_sc_hd__clkbuf_4
X_8158_ _8158_/CLK _8158_/D vssd1 vssd1 vccd1 vccd1 _8158_/Q sky130_fd_sc_hd__dfxtp_1
X_8089_ _8089_/CLK _8089_/D vssd1 vssd1 vccd1 vccd1 _8089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8502__252 vssd1 vssd1 vccd1 vccd1 partID[2] _8502__252/LO sky130_fd_sc_hd__conb_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6537__257 _6539__259/A vssd1 vssd1 vccd1 vccd1 _7897_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4810_ _4926_/B _4774_/X _4786_/X _4809_/X vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__a31o_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6891__410 _6891__410/A vssd1 vssd1 vccd1 vccd1 _8086_/CLK sky130_fd_sc_hd__inv_2
X_5790_ _5790_/A vssd1 vssd1 vccd1 vccd1 _7795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4735_/X _4737_/X _4740_/X _4721_/X _4746_/A vssd1 vssd1 vccd1 vccd1 _4741_/X
+ sky130_fd_sc_hd__o221a_1
X_4672_ _4668_/X _4671_/X _4735_/A vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__mux2_1
X_7460_ _7557_/A _7460_/B vssd1 vssd1 vccd1 vccd1 _7487_/B sky130_fd_sc_hd__nand2_1
X_6411_ _7827_/Q _6401_/X _6371_/A _6410_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _7827_/D
+ sky130_fd_sc_hd__a221o_1
X_6342_ _7812_/Q _6286_/X _6341_/X vssd1 vssd1 vccd1 vccd1 _7812_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8012_ _8012_/CLK _8012_/D vssd1 vssd1 vccd1 vccd1 _8012_/Q sky130_fd_sc_hd__dfxtp_1
X_5224_ _5224_/A _5224_/B vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__or2_1
X_5155_ _5187_/A _5150_/X _5152_/X _5154_/X _5159_/A vssd1 vssd1 vccd1 vccd1 _5155_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5086_ _5031_/X _5058_/X _5068_/X _5085_/X vssd1 vssd1 vccd1 vccd1 _5086_/X sky130_fd_sc_hd__a31o_2
X_4106_ _8128_/Q vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4037_ _8384_/Q _4010_/X _4037_/S vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5988_ _5988_/A vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__clkbuf_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7727_ _7727_/CLK _7727_/D vssd1 vssd1 vccd1 vccd1 _7727_/Q sky130_fd_sc_hd__dfxtp_1
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _8120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7658_ _7658_/A vssd1 vssd1 vccd1 vccd1 _7659_/C sky130_fd_sc_hd__clkinv_2
X_6609_ _6609_/A vssd1 vssd1 vccd1 vccd1 _7952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7589_ _8438_/Q _7595_/B vssd1 vssd1 vccd1 vccd1 _7589_/X sky130_fd_sc_hd__or2_1
XFILLER_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput180 _6064_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput191 _6102_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
XFILLER_102_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3399_ clkbuf_0__3399_/X vssd1 vssd1 vccd1 vccd1 _7044_/A sky130_fd_sc_hd__clkbuf_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7379__140 _7379__140/A vssd1 vssd1 vccd1 vccd1 _8351_/CLK sky130_fd_sc_hd__inv_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5911_ _5911_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__or2_4
X_5842_ _5842_/A vssd1 vssd1 vccd1 vccd1 _7729_/D sky130_fd_sc_hd__clkbuf_1
X_5773_ _4150_/X _7802_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7512_ _7512_/A vssd1 vssd1 vccd1 vccd1 _8413_/D sky130_fd_sc_hd__clkbuf_1
X_4724_ _4612_/X _8138_/Q _4924_/A _4723_/X _4678_/X vssd1 vssd1 vccd1 vccd1 _4724_/X
+ sky130_fd_sc_hd__a221o_1
X_8492_ _8496_/CLK _8492_/D vssd1 vssd1 vccd1 vccd1 _8492_/Q sky130_fd_sc_hd__dfxtp_1
X_4655_ _4721_/A vssd1 vssd1 vccd1 vccd1 _4883_/A sky130_fd_sc_hd__buf_2
XFILLER_116_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7374_ _7380_/A vssd1 vssd1 vccd1 vccd1 _7374_/X sky130_fd_sc_hd__buf_1
X_4586_ _4428_/X _8151_/Q _4586_/S vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__mux2_1
Xinput71 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _7693_/A sky130_fd_sc_hd__buf_4
Xinput82 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__clkbuf_2
Xinput60 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _3844_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_107_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput93 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__buf_4
X_6325_ _6774_/A _6293_/A _6299_/X vssd1 vssd1 vccd1 vccd1 _6325_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7041__523 _7041__523/A vssd1 vssd1 vccd1 vccd1 _8204_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__clkbuf_2
X_6187_ _6184_/X _7963_/Q _6186_/X _6180_/X _7752_/Q vssd1 vssd1 vccd1 vccd1 _7752_/D
+ sky130_fd_sc_hd__o32a_1
X_5138_ _3928_/X _5022_/X _5137_/X _5091_/X vssd1 vssd1 vccd1 vccd1 _8084_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5069_ _5108_/A vssd1 vssd1 vccd1 vccd1 _5152_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6985__477 _6985__477/A vssd1 vssd1 vccd1 vccd1 _8158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _8212_/Q _4439_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4371_ _4371_/A vssd1 vssd1 vccd1 vccd1 _8238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6110_ _7758_/Q _6095_/X _6099_/X _6108_/X _6109_/X vssd1 vssd1 vccd1 vccd1 _6110_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6034_/X _6039_/X _6040_/X _6037_/X vssd1 vssd1 vccd1 vccd1 _6041_/X sky130_fd_sc_hd__o211a_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7992_ _7992_/CLK _7992_/D vssd1 vssd1 vccd1 vccd1 _7992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5825_ _7779_/Q _5571_/A _5825_/S vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5756_ _5756_/A vssd1 vssd1 vccd1 vccd1 _7859_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3623_ _7417_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3623_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5687_ _7889_/Q _4993_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__mux2_1
X_4707_ _4637_/X _4706_/X _4883_/A vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__a21o_1
X_8475_ _8481_/CLK _8475_/D vssd1 vssd1 vccd1 vccd1 _8475_/Q sky130_fd_sc_hd__dfxtp_1
X_4638_ _4650_/A vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__buf_2
X_7360__125 _7360__125/A vssd1 vssd1 vccd1 vccd1 _8336_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4569_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5655_/A sky130_fd_sc_hd__clkbuf_2
X_7288_ _7297_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _8304_/D sky130_fd_sc_hd__nor2_1
X_6308_ _6312_/B _6308_/B vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__or2_1
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6239_ _8287_/Q vssd1 vssd1 vccd1 vccd1 _7320_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7006__495 _7006__495/A vssd1 vssd1 vccd1 vccd1 _8176_/CLK sky130_fd_sc_hd__inv_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3236_ clkbuf_0__3236_/X vssd1 vssd1 vccd1 vccd1 _6588__299/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8545__244 vssd1 vssd1 vccd1 vccd1 _8545__244/HI partID[12] sky130_fd_sc_hd__conb_1
XFILLER_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3940_ _8443_/Q vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3440_ clkbuf_0__3440_/X vssd1 vssd1 vccd1 vccd1 _7119__85/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3871_ _3893_/S vssd1 vssd1 vccd1 vccd1 _3884_/S sky130_fd_sc_hd__buf_2
XFILLER_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5610_ _5610_/A vssd1 vssd1 vccd1 vccd1 _7924_/D sky130_fd_sc_hd__clkbuf_1
X_6590_ _6915_/A vssd1 vssd1 vccd1 vccd1 _6590_/X sky130_fd_sc_hd__buf_1
X_5541_ _7951_/Q _4973_/X _5549_/S vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8260_ _8260_/CLK _8260_/D vssd1 vssd1 vccd1 vccd1 _8260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5472_ _8005_/Q _4350_/A _5476_/S vssd1 vssd1 vccd1 vccd1 _5473_/A sky130_fd_sc_hd__mux2_1
X_7211_ _7211_/A _7211_/B _7211_/C vssd1 vssd1 vccd1 vccd1 _7241_/A sky130_fd_sc_hd__nand3_2
X_8191_ _8191_/CLK _8191_/D vssd1 vssd1 vccd1 vccd1 _8191_/Q sky130_fd_sc_hd__dfxtp_1
X_4423_ _4422_/X _8217_/Q _4429_/S vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__mux2_1
X_4354_ _4353_/X _8243_/Q _4357_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__mux2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4285_ _8271_/Q _4200_/X _4285_/S vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__mux2_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _7810_/Q input25/X _6039_/S vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__mux2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7975_ _8441_/CLK _7975_/D vssd1 vssd1 vccd1 vccd1 _7975_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6857_ _8436_/Q _6863_/B vssd1 vssd1 vccd1 vccd1 _6858_/A sky130_fd_sc_hd__and2_1
X_5808_ _5808_/A vssd1 vssd1 vccd1 vccd1 _7787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6788_ _6767_/Y _6768_/X _6781_/X _6785_/X _6787_/X vssd1 vssd1 vccd1 vccd1 _6794_/C
+ sky130_fd_sc_hd__o2111a_1
X_5739_ _7866_/Q _5574_/A _5743_/S vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8458_ _8458_/CLK _8458_/D vssd1 vssd1 vccd1 vccd1 _8458_/Q sky130_fd_sc_hd__dfxtp_1
X_8389_ _8389_/CLK _8389_/D vssd1 vssd1 vccd1 vccd1 _8389_/Q sky130_fd_sc_hd__dfxtp_1
X_8529__228 vssd1 vssd1 vccd1 vccd1 _8529__228/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6869__392 _6872__395/A vssd1 vssd1 vccd1 vccd1 _8068_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3399_ _6915_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3399_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_40 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_51 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_62 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_84 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_73 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_95 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054__533 _7054__533/A vssd1 vssd1 vccd1 vccd1 _8214_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3219_ clkbuf_0__3219_/X vssd1 vssd1 vccd1 vccd1 _6510_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7456__26 _7620__30/A vssd1 vssd1 vccd1 vccd1 _8412_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6586__297 _6588__299/A vssd1 vssd1 vccd1 vccd1 _7937_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4070_ _4070_/A vssd1 vssd1 vccd1 vccd1 _8371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A vssd1 vssd1 vccd1 vccd1 _8105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7760_ _8433_/CLK _7760_/D vssd1 vssd1 vccd1 vccd1 _7760_/Q sky130_fd_sc_hd__dfxtp_1
X_3923_ _3916_/X _8457_/Q _3935_/S vssd1 vssd1 vccd1 vccd1 _3924_/A sky130_fd_sc_hd__mux2_1
X_7691_ _7689_/Y _7690_/Y _7678_/X vssd1 vssd1 vccd1 vccd1 _8488_/D sky130_fd_sc_hd__a21oi_1
X_6711_ _6711_/A vssd1 vssd1 vccd1 vccd1 _8016_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3423_ clkbuf_0__3423_/X vssd1 vssd1 vccd1 vccd1 _7034__517/A sky130_fd_sc_hd__clkbuf_4
X_6642_ _6642_/A _6642_/B vssd1 vssd1 vccd1 vccd1 _6658_/S sky130_fd_sc_hd__and2_4
X_3854_ _6415_/B _6294_/A vssd1 vssd1 vccd1 vccd1 _6287_/A sky130_fd_sc_hd__or2b_1
X_8312_ _8499_/CLK _8312_/D vssd1 vssd1 vccd1 vccd1 _8312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3285_ clkbuf_0__3285_/X vssd1 vssd1 vccd1 vccd1 _6723__358/A sky130_fd_sc_hd__clkbuf_4
X_5524_ _5349_/X _7982_/Q _5530_/S vssd1 vssd1 vccd1 vccd1 _5525_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5455_ _5455_/A vssd1 vssd1 vccd1 vccd1 _8013_/D sky130_fd_sc_hd__clkbuf_1
X_8243_ _8243_/CLK _8243_/D vssd1 vssd1 vccd1 vccd1 _8243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8174_ _8174_/CLK _8174_/D vssd1 vssd1 vccd1 vccd1 _8174_/Q sky130_fd_sc_hd__dfxtp_1
X_4406_ _5709_/A _5833_/A vssd1 vssd1 vccd1 vccd1 _4429_/S sky130_fd_sc_hd__or2_2
X_5386_ _5361_/X _8047_/Q _5386_/S vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4337_ _4337_/A vssd1 vssd1 vccd1 vccd1 _8249_/D sky130_fd_sc_hd__clkbuf_1
X_4268_ _4268_/A vssd1 vssd1 vccd1 vccd1 _8279_/D sky130_fd_sc_hd__clkbuf_1
X_6007_ _6007_/A vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__clkbuf_1
X_4199_ _4199_/A vssd1 vssd1 vccd1 vccd1 _8334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7958_ _8496_/CLK _7958_/D vssd1 vssd1 vccd1 vccd1 _7958_/Q sky130_fd_sc_hd__dfxtp_1
X_7889_ _7889_/CLK _7889_/D vssd1 vssd1 vccd1 vccd1 _7889_/Q sky130_fd_sc_hd__dfxtp_1
X_6909_ _6909_/A vssd1 vssd1 vccd1 vccd1 _6909_/X sky130_fd_sc_hd__buf_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7373__135 _7373__135/A vssd1 vssd1 vccd1 vccd1 _8346_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _8399_/Q _5163_/X _5224_/A _5238_/X _5239_/X vssd1 vssd1 vccd1 vccd1 _5240_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256__193 _6258__195/A vssd1 vssd1 vccd1 vccd1 _7785_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5171_ _5215_/A vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4118_/X _4120_/Y _4607_/B vssd1 vssd1 vccd1 vccd1 _4129_/B sky130_fd_sc_hd__mux2_1
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _8378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7812_ _8497_/CLK _7812_/D vssd1 vssd1 vccd1 vccd1 _7812_/Q sky130_fd_sc_hd__dfxtp_1
X_4955_ _5539_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _4971_/S sky130_fd_sc_hd__nor2_2
X_7743_ _8490_/CLK _7743_/D vssd1 vssd1 vccd1 vccd1 _7743_/Q sky130_fd_sc_hd__dfxtp_1
X_3906_ _8462_/Q _3880_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4886_ _4757_/X _4884_/X _4885_/X vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1_0__3406_ clkbuf_0__3406_/X vssd1 vssd1 vccd1 vccd1 _6970_/A sky130_fd_sc_hd__clkbuf_4
X_7674_ _8484_/Q _7692_/B vssd1 vssd1 vccd1 vccd1 _7674_/Y sky130_fd_sc_hd__nand2_1
X_6625_ _6640_/S vssd1 vssd1 vccd1 vccd1 _6634_/S sky130_fd_sc_hd__clkbuf_2
X_3837_ _8074_/Q _3920_/B _5018_/A _3836_/Y vssd1 vssd1 vccd1 vccd1 _3838_/D sky130_fd_sc_hd__a31o_1
XFILLER_118_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _5507_/A vssd1 vssd1 vccd1 vccd1 _7990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8226_ _8226_/CLK _8226_/D vssd1 vssd1 vccd1 vccd1 _8226_/Q sky130_fd_sc_hd__dfxtp_1
X_5438_ _8023_/Q _4442_/X _5440_/S vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3236_ _6584_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3236_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3622_ clkbuf_0__3622_/X vssd1 vssd1 vccd1 vccd1 _7416__170/A sky130_fd_sc_hd__clkbuf_4
X_5369_ _5577_/A vssd1 vssd1 vccd1 vccd1 _5369_/X sky130_fd_sc_hd__clkbuf_2
X_8157_ _8157_/CLK _8157_/D vssd1 vssd1 vccd1 vccd1 _8157_/Q sky130_fd_sc_hd__dfxtp_1
X_7108_ _7120_/A vssd1 vssd1 vccd1 vccd1 _7108_/X sky130_fd_sc_hd__buf_1
X_8088_ _8442_/CLK _8088_/D vssd1 vssd1 vccd1 vccd1 _8088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6698__343 _6698__343/A vssd1 vssd1 vccd1 vccd1 _8007_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4738_/X _4739_/X _4740_/S vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4671_ _8198_/Q _7999_/Q _7935_/Q _7895_/Q _4669_/X _4670_/X vssd1 vssd1 vccd1 vccd1
+ _4671_/X sky130_fd_sc_hd__mux4_1
X_6410_ _8480_/Q _6412_/B _6410_/C vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__and3_1
X_6341_ _6289_/A _6338_/X _6340_/X _6369_/A vssd1 vssd1 vccd1 vccd1 _6341_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6272_ _6278_/A vssd1 vssd1 vccd1 vccd1 _6272_/X sky130_fd_sc_hd__buf_1
XFILLER_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8011_ _8011_/CLK _8011_/D vssd1 vssd1 vccd1 vccd1 _8011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5223_ _8407_/Q _8145_/Q _5261_/S vssd1 vssd1 vccd1 vccd1 _5224_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5154_ _5074_/X _5153_/X _5113_/X vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4105_ _4475_/B _5538_/B _5538_/A vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__or3b_2
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5085_ _5072_/X _5077_/X _5082_/X _5083_/X _5159_/A vssd1 vssd1 vccd1 vccd1 _5085_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4036_ _4036_/A vssd1 vssd1 vccd1 vccd1 _8385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5987_ _7963_/Q _5993_/B vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__and2_2
XFILLER_40_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7726_ _7726_/CLK _7726_/D vssd1 vssd1 vccd1 vccd1 _7726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4938_ _8120_/Q _4223_/X _4946_/S vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__mux2_1
X_7657_ _7703_/A vssd1 vssd1 vccd1 vccd1 _7657_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4869_ _4613_/A _8134_/Q _4925_/A _4868_/X _4678_/A vssd1 vssd1 vccd1 vccd1 _4869_/X
+ sky130_fd_sc_hd__a221o_1
X_6608_ _7699_/A _7952_/Q _6616_/S vssd1 vssd1 vccd1 vccd1 _6609_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7588_ _8438_/Q _7578_/X _7587_/X _7582_/X vssd1 vssd1 vccd1 vccd1 _8437_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput170 _5865_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8209_ _8209_/CLK _8209_/D vssd1 vssd1 vccd1 vccd1 _8209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3219_ _6497_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3219_/X sky130_fd_sc_hd__clkbuf_16
Xoutput181 _6068_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput192 _6104_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6543__262 _6544__263/A vssd1 vssd1 vccd1 vccd1 _7902_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3398_ clkbuf_0__3398_/X vssd1 vssd1 vccd1 vccd1 _6911__422/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8509__259 vssd1 vssd1 vccd1 vccd1 partID[15] _8509__259/LO sky130_fd_sc_hd__conb_1
X_6849__390 _6849__390/A vssd1 vssd1 vccd1 vccd1 _8058_/CLK sky130_fd_sc_hd__inv_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6706__350 _6706__350/A vssd1 vssd1 vccd1 vccd1 _8014_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5910_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _4144_/X _7729_/Q _5843_/S vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__mux2_1
X_5772_ _5772_/A vssd1 vssd1 vccd1 vccd1 _7803_/D sky130_fd_sc_hd__clkbuf_1
X_4723_ _4622_/X _4708_/X _4712_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__a31o_1
X_7511_ _7490_/Y _7575_/A _7511_/C _7511_/D vssd1 vssd1 vccd1 vccd1 _7512_/A sky130_fd_sc_hd__and4b_1
X_8491_ _8498_/CLK _8491_/D vssd1 vssd1 vccd1 vccd1 _8491_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7442_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7442_/X sky130_fd_sc_hd__buf_1
X_4654_ _4674_/B _4654_/B vssd1 vssd1 vccd1 vccd1 _4721_/A sky130_fd_sc_hd__nor2_2
Xinput50 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _3842_/C sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _7690_/A sky130_fd_sc_hd__buf_4
X_4585_ _4585_/A vssd1 vssd1 vccd1 vccd1 _8152_/D sky130_fd_sc_hd__clkbuf_1
Xinput83 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__buf_4
X_6324_ _8497_/Q vssd1 vssd1 vccd1 vccd1 _6774_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5206_ _3934_/X _5022_/X _5205_/X _5091_/X vssd1 vssd1 vccd1 vccd1 _8082_/D sky130_fd_sc_hd__o211a_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6486__216 _6488__218/A vssd1 vssd1 vccd1 vccd1 _7856_/CLK sky130_fd_sc_hd__inv_2
X_6186_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6186_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5137_ _8084_/Q _5024_/X _5331_/A _5136_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5137_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _5038_/X _5061_/X _5067_/X vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _8390_/Q _4018_/X _4023_/S vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7709_ _7611_/A _7707_/B _7704_/Y vssd1 vssd1 vccd1 vccd1 _7709_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7018__504 _7019__505/A vssd1 vssd1 vccd1 vccd1 _8185_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4342_/X _8238_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4371_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6040_ _7739_/Q _6044_/B vssd1 vssd1 vccd1 vccd1 _6040_/X sky130_fd_sc_hd__or2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7991_ _7991_/CLK _7991_/D vssd1 vssd1 vccd1 vccd1 _7991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ _6942_/A vssd1 vssd1 vccd1 vccd1 _6942_/X sky130_fd_sc_hd__buf_1
XFILLER_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6600__307 _6600__307/A vssd1 vssd1 vccd1 vccd1 _7947_/CLK sky130_fd_sc_hd__inv_2
X_6873_ _6873_/A vssd1 vssd1 vccd1 vccd1 _6873_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_16_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8425_/CLK sky130_fd_sc_hd__clkbuf_16
X_5824_ _5824_/A vssd1 vssd1 vccd1 vccd1 _7780_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3622_ _7411_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3622_/X sky130_fd_sc_hd__clkbuf_16
X_5755_ _7859_/Q _5571_/A _5755_/S vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5686_ _5686_/A vssd1 vssd1 vccd1 vccd1 _7890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8474_ _8478_/CLK _8474_/D vssd1 vssd1 vccd1 vccd1 _8474_/Q sky130_fd_sc_hd__dfxtp_1
X_4706_ _8164_/Q _8156_/Q _8118_/Q _8188_/Q _4650_/X _4651_/X vssd1 vssd1 vccd1 vccd1
+ _4706_/X sky130_fd_sc_hd__mux4_2
X_4637_ _4740_/S vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__clkbuf_2
X_6830__375 _6830__375/A vssd1 vssd1 vccd1 vccd1 _8043_/CLK sky130_fd_sc_hd__inv_2
X_4568_ _4568_/A vssd1 vssd1 vccd1 vccd1 _8159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4499_ _8190_/Q _4223_/X _4507_/S vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__mux2_1
X_7287_ _8304_/Q _7280_/X _7286_/X _7172_/B vssd1 vssd1 vccd1 vccd1 _7288_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6307_ _6310_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _6318_/A sky130_fd_sc_hd__nor2_1
X_6238_ _8315_/Q _6238_/B vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__and2b_1
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3235_ clkbuf_0__3235_/X vssd1 vssd1 vccd1 vccd1 _6580__292/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6991__482 _6991__482/A vssd1 vssd1 vccd1 vccd1 _8163_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6250__188 _6252__190/A vssd1 vssd1 vccd1 vccd1 _7780_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7640__46 _7644__50/A vssd1 vssd1 vccd1 vccd1 _8469_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3870_ _4457_/A _4083_/A vssd1 vssd1 vccd1 vccd1 _3893_/S sky130_fd_sc_hd__nor2_2
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5540_ _5555_/S vssd1 vssd1 vccd1 vccd1 _5549_/S sky130_fd_sc_hd__buf_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5471_ _5471_/A vssd1 vssd1 vccd1 vccd1 _8006_/D sky130_fd_sc_hd__clkbuf_1
X_7210_ _8487_/Q _7195_/Y _7197_/X _7200_/X _7209_/X vssd1 vssd1 vccd1 vccd1 _7210_/X
+ sky130_fd_sc_hd__o2111a_1
X_4422_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__clkbuf_2
X_8190_ _8190_/CLK _8190_/D vssd1 vssd1 vccd1 vccd1 _8190_/Q sky130_fd_sc_hd__dfxtp_1
X_4353_ _4353_/A vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__buf_2
X_4284_ _4284_/A vssd1 vssd1 vccd1 vccd1 _8272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _6061_/A vssd1 vssd1 vccd1 vccd1 _6039_/S sky130_fd_sc_hd__buf_2
XFILLER_100_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7974_ _8439_/CLK _7974_/D vssd1 vssd1 vccd1 vccd1 _7974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6856_ _6856_/A vssd1 vssd1 vccd1 vccd1 _8061_/D sky130_fd_sc_hd__clkbuf_1
X_3999_ _8395_/Q _3998_/X _4011_/S vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__mux2_1
X_5807_ _3883_/X _7787_/Q _5807_/S vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__mux2_1
X_6787_ _7197_/A _7478_/B vssd1 vssd1 vccd1 vccd1 _6787_/X sky130_fd_sc_hd__xor2_1
X_5738_ _5738_/A vssd1 vssd1 vccd1 vccd1 _7867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5577_/X _7897_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5670_/A sky130_fd_sc_hd__mux2_1
X_8457_ _8457_/CLK _8457_/D vssd1 vssd1 vccd1 vccd1 _8457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8388_ _8388_/CLK _8388_/D vssd1 vssd1 vccd1 vccd1 _8388_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3398_ _6909_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3398_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7339_ _8321_/Q _7343_/B vssd1 vssd1 vccd1 vccd1 _7339_/X sky130_fd_sc_hd__or2_1
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_52 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_30 _6108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_41 _6117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_63 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_85 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_74 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_96 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6499__226 _6500__227/A vssd1 vssd1 vccd1 vccd1 _7866_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3218_ clkbuf_0__3218_/X vssd1 vssd1 vccd1 vccd1 _6496__225/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6692__338 _6692__338/A vssd1 vssd1 vccd1 vccd1 _8002_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8512__211 vssd1 vssd1 vccd1 vccd1 _8512__211/HI caravel_irq[2] sky130_fd_sc_hd__conb_1
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998__488 _6999__489/A vssd1 vssd1 vccd1 vccd1 _8169_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ _8105_/Q _4247_/X _4971_/S vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__mux2_1
X_3922_ _3944_/S vssd1 vssd1 vccd1 vccd1 _3935_/S sky130_fd_sc_hd__buf_2
X_7690_ _7690_/A _7693_/B vssd1 vssd1 vccd1 vccd1 _7690_/Y sky130_fd_sc_hd__nand2_1
X_6710_ _8016_/Q _6207_/A _6714_/S vssd1 vssd1 vccd1 vccd1 _6711_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3422_ clkbuf_0__3422_/X vssd1 vssd1 vccd1 vccd1 _7031__515/A sky130_fd_sc_hd__clkbuf_4
X_6641_ _6641_/A vssd1 vssd1 vccd1 vccd1 _7967_/D sky130_fd_sc_hd__clkbuf_1
X_3853_ _7853_/Q vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6572_ _6578_/A vssd1 vssd1 vccd1 vccd1 _6572_/X sky130_fd_sc_hd__buf_1
X_8311_ _8499_/CLK _8311_/D vssd1 vssd1 vccd1 vccd1 _8311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5523_ _5523_/A vssd1 vssd1 vccd1 vccd1 _7983_/D sky130_fd_sc_hd__clkbuf_1
X_5454_ _8013_/Q _4439_/X _5458_/S vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__mux2_1
X_8242_ _8242_/CLK _8242_/D vssd1 vssd1 vccd1 vccd1 _8242_/Q sky130_fd_sc_hd__dfxtp_1
X_8173_ _8173_/CLK _8173_/D vssd1 vssd1 vccd1 vccd1 _8173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5385_ _5385_/A vssd1 vssd1 vccd1 vccd1 _8048_/D sky130_fd_sc_hd__clkbuf_1
X_4405_ _4903_/B _4405_/B _4904_/A vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__or3b_4
X_4336_ _8249_/Q _4194_/X _4340_/S vssd1 vssd1 vccd1 vccd1 _4337_/A sky130_fd_sc_hd__mux2_1
X_4267_ _8279_/Q _4200_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6006_ _7971_/Q _6006_/B vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__and2_1
X_4198_ _8334_/Q _4197_/X _4201_/S vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__mux2_1
X_6268__202 _6268__202/A vssd1 vssd1 vccd1 vccd1 _7794_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7957_ _8489_/CLK _7957_/D vssd1 vssd1 vccd1 vccd1 _7957_/Q sky130_fd_sc_hd__dfxtp_1
X_7888_ _7888_/CLK _7888_/D vssd1 vssd1 vccd1 vccd1 _7888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7407__162 _7410__165/A vssd1 vssd1 vccd1 vccd1 _8373_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6843__385 _6843__385/A vssd1 vssd1 vccd1 vccd1 _8053_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6507__233 _6508__234/A vssd1 vssd1 vccd1 vccd1 _7873_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6700__345 _6700__345/A vssd1 vssd1 vccd1 vccd1 _8009_/CLK sky130_fd_sc_hd__inv_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3430_ clkbuf_0__3430_/X vssd1 vssd1 vccd1 vccd1 _7074__550/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5170_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4121_ _8131_/Q _8126_/Q vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__xor2_1
X_4052_ _8378_/Q _4002_/X _4056_/S vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7811_ _8497_/CLK _7811_/D vssd1 vssd1 vccd1 vccd1 _7811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4954_ _4999_/C _4999_/B _4999_/A vssd1 vssd1 vccd1 vccd1 _5727_/B sky130_fd_sc_hd__nand3b_4
X_7742_ _8490_/CLK _7742_/D vssd1 vssd1 vccd1 vccd1 _7742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3905_ _3905_/A vssd1 vssd1 vccd1 vccd1 _8463_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3628_ clkbuf_0__3628_/X vssd1 vssd1 vccd1 vccd1 _7447__20/A sky130_fd_sc_hd__clkbuf_16
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _8183_/Q _4789_/A _4790_/X _8159_/Q _4715_/A vssd1 vssd1 vccd1 vccd1 _4885_/X
+ sky130_fd_sc_hd__o221a_1
X_7673_ _7698_/B vssd1 vssd1 vccd1 vccd1 _7692_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3405_ clkbuf_0__3405_/X vssd1 vssd1 vccd1 vccd1 _6944__447/A sky130_fd_sc_hd__clkbuf_4
X_6624_ _6624_/A _6642_/B vssd1 vssd1 vccd1 vccd1 _6640_/S sky130_fd_sc_hd__nand2_2
X_3836_ _5019_/B _5316_/A _3826_/Y vssd1 vssd1 vccd1 vccd1 _3836_/Y sky130_fd_sc_hd__a21oi_1
X_6716__352 _6718__354/A vssd1 vssd1 vccd1 vccd1 _8019_/CLK sky130_fd_sc_hd__inv_2
X_5506_ _7990_/Q _4347_/A _5512_/S vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8225_ _8225_/CLK _8225_/D vssd1 vssd1 vccd1 vccd1 _8225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5437_ _5437_/A vssd1 vssd1 vccd1 vccd1 _8024_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3235_ _6578_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3235_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5368_ _8061_/Q vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3621_ clkbuf_0__3621_/X vssd1 vssd1 vccd1 vccd1 _7409__164/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8156_ _8156_/CLK _8156_/D vssd1 vssd1 vccd1 vccd1 _8156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7107_ _7107_/A vssd1 vssd1 vccd1 vccd1 _7107_/X sky130_fd_sc_hd__buf_1
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _8257_/D sky130_fd_sc_hd__clkbuf_1
X_5299_ _8263_/Q _5178_/X _5285_/B _8255_/Q _5098_/A vssd1 vssd1 vccd1 vccd1 _5299_/X
+ sky130_fd_sc_hd__o221a_1
X_8087_ _8478_/CLK _8087_/D vssd1 vssd1 vccd1 vccd1 _8087_/Q sky130_fd_sc_hd__dfxtp_1
X_7038_ _7038_/A vssd1 vssd1 vccd1 vccd1 _7038_/X sky130_fd_sc_hd__buf_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7131__95 _7131__95/A vssd1 vssd1 vccd1 vccd1 _8276_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4670_/A vssd1 vssd1 vccd1 vccd1 _4670_/X sky130_fd_sc_hd__buf_2
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7067__544 _7068__545/A vssd1 vssd1 vccd1 vccd1 _8225_/CLK sky130_fd_sc_hd__inv_2
X_6340_ _8477_/Q _6311_/X _6339_/X _6306_/X _6352_/A vssd1 vssd1 vccd1 vccd1 _6340_/X
+ sky130_fd_sc_hd__a221o_1
X_8010_ _8010_/CLK _8010_/D vssd1 vssd1 vccd1 vccd1 _8010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _8375_/Q _5216_/X _5336_/B _5221_/X vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__o211a_1
X_5153_ _8171_/Q _8147_/Q _8409_/Q _8179_/Q _5123_/A _5111_/X vssd1 vssd1 vccd1 vccd1
+ _5153_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ _8131_/Q vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _8072_/Q _5084_/B vssd1 vssd1 vccd1 vccd1 _5159_/A sky130_fd_sc_hd__xnor2_4
X_4035_ _8385_/Q _4006_/X _4037_/S vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _5986_/A vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__clkbuf_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7725_ _7725_/CLK _7725_/D vssd1 vssd1 vccd1 vccd1 _7725_/Q sky130_fd_sc_hd__dfxtp_1
X_4937_ _4952_/S vssd1 vssd1 vccd1 vccd1 _4946_/S sky130_fd_sc_hd__buf_2
X_4868_ _4926_/B _4848_/X _4854_/X _4867_/X vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7656_ _7656_/A vssd1 vssd1 vccd1 vccd1 _7656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6607_ _6622_/S vssd1 vssd1 vccd1 vccd1 _6616_/S sky130_fd_sc_hd__clkbuf_2
X_3819_ _8073_/Q vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ _8352_/Q _4619_/A _4765_/A _8328_/Q _4798_/X vssd1 vssd1 vccd1 vccd1 _4799_/X
+ sky130_fd_sc_hd__o221a_1
X_7587_ _8437_/Q _7595_/B vssd1 vssd1 vccd1 vccd1 _7587_/X sky130_fd_sc_hd__or2_1
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6469_ _7851_/Q _7966_/Q _6714_/S vssd1 vssd1 vccd1 vccd1 _6470_/A sky130_fd_sc_hd__mux2_1
Xoutput160 _5881_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8208_ _8208_/CLK _8208_/D vssd1 vssd1 vccd1 vccd1 _8208_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput171 _5867_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
Xclkbuf_0__3218_ _6491_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3218_/X sky130_fd_sc_hd__clkbuf_16
Xoutput182 _6071_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput193 _6106_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
X_8139_ _8139_/CLK _8139_/D vssd1 vssd1 vccd1 vccd1 _8139_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3550_ clkbuf_0__3550_/X vssd1 vssd1 vccd1 vccd1 _7259__113/A sky130_fd_sc_hd__clkbuf_16
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3397_ clkbuf_0__3397_/X vssd1 vssd1 vccd1 vccd1 _6906__418/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7104__73 _7104__73/A vssd1 vssd1 vccd1 vccd1 _8254_/CLK sky130_fd_sc_hd__inv_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _7730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5771_ _4147_/X _7803_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5772_/A sky130_fd_sc_hd__mux2_1
X_4722_ _4714_/X _4717_/X _4720_/X _4721_/X _4746_/A vssd1 vssd1 vccd1 vccd1 _4722_/X
+ sky130_fd_sc_hd__o221a_1
X_8490_ _8490_/CLK _8490_/D vssd1 vssd1 vccd1 vccd1 _8490_/Q sky130_fd_sc_hd__dfxtp_2
X_7510_ _7510_/A _7510_/B vssd1 vssd1 vccd1 vccd1 _7511_/D sky130_fd_sc_hd__nand2_1
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4653_ _4653_/A _4653_/B vssd1 vssd1 vccd1 vccd1 _4654_/B sky130_fd_sc_hd__nor2_1
Xinput40 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__buf_4
Xinput51 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _3846_/B sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__clkbuf_8
X_4584_ _4425_/X _8152_/Q _4586_/S vssd1 vssd1 vccd1 vccd1 _4585_/A sky130_fd_sc_hd__mux2_1
Xinput95 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _7607_/A sky130_fd_sc_hd__buf_6
Xinput84 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6323_ _7809_/Q _6286_/X _6322_/X vssd1 vssd1 vccd1 vccd1 _7809_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5205_ _8082_/Q _5025_/A _5246_/A _5204_/X _5088_/A vssd1 vssd1 vccd1 vccd1 _5205_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6185_ _6184_/X _7962_/Q _6178_/X _6180_/X _7751_/Q vssd1 vssd1 vccd1 vccd1 _7751_/D
+ sky130_fd_sc_hd__o32a_1
X_5136_ _5031_/X _5122_/X _5127_/X _5135_/X vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__a31o_2
X_5067_ _5062_/X _5065_/X _5104_/A vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4362_/A vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _5969_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__and2_1
XFILLER_80_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7708_ _6792_/A _7704_/Y _7707_/X _6194_/X vssd1 vssd1 vccd1 vccd1 _8493_/D sky130_fd_sc_hd__a211o_1
XFILLER_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7639_ _7639_/A vssd1 vssd1 vccd1 vccd1 _7639_/X sky130_fd_sc_hd__buf_1
XFILLER_21_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7259__113 _7259__113/A vssd1 vssd1 vccd1 vccd1 _8296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6922__430 _6922__430/A vssd1 vssd1 vccd1 vccd1 _8108_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7990_ _7990_/CLK _7990_/D vssd1 vssd1 vccd1 vccd1 _7990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5823_ _7780_/Q _5568_/A _5825_/S vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3621_ _7405_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3621_/X sky130_fd_sc_hd__clkbuf_16
X_5754_ _5754_/A vssd1 vssd1 vccd1 vccd1 _7860_/D sky130_fd_sc_hd__clkbuf_1
X_8473_ _8473_/CLK _8473_/D vssd1 vssd1 vccd1 vccd1 _8473_/Q sky130_fd_sc_hd__dfxtp_1
X_5685_ _7890_/Q _4990_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__mux2_1
X_6492__221 _6494__223/A vssd1 vssd1 vccd1 vccd1 _7861_/CLK sky130_fd_sc_hd__inv_2
X_4705_ _8330_/Q _8220_/Q _7877_/Q _8354_/Q _4630_/X _4633_/X vssd1 vssd1 vccd1 vccd1
+ _4705_/X sky130_fd_sc_hd__mux4_1
X_7424_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7424_/X sky130_fd_sc_hd__buf_1
X_4636_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4740_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7355_ _7355_/A vssd1 vssd1 vccd1 vccd1 _7355_/X sky130_fd_sc_hd__buf_1
X_4567_ _4428_/X _8159_/Q _4567_/S vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__mux2_1
X_6306_ _6355_/B vssd1 vssd1 vccd1 vccd1 _6306_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4498_ _4513_/S vssd1 vssd1 vccd1 vccd1 _4507_/S sky130_fd_sc_hd__buf_2
X_7286_ _7286_/A vssd1 vssd1 vccd1 vccd1 _7286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6237_ _8316_/Q _8317_/Q _8318_/Q _8319_/Q _8313_/Q _8314_/Q vssd1 vssd1 vccd1 vccd1
+ _6238_/B sky130_fd_sc_hd__mux4_1
X_7401__157 _7401__157/A vssd1 vssd1 vccd1 vccd1 _8368_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6167_/X _7952_/Q _6161_/X _6163_/X _7741_/Q vssd1 vssd1 vccd1 vccd1 _7741_/D
+ sky130_fd_sc_hd__o32a_1
X_5119_ _8362_/Q _8346_/Q _8338_/Q _8370_/Q _5060_/X _5044_/X vssd1 vssd1 vccd1 vccd1
+ _5119_/X sky130_fd_sc_hd__mux4_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6099_ _6112_/A vssd1 vssd1 vccd1 vccd1 _6099_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3234_ clkbuf_0__3234_/X vssd1 vssd1 vccd1 vccd1 _6577__290/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6501__228 _6503__230/A vssd1 vssd1 vccd1 vccd1 _7868_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6556__273 _6558__275/A vssd1 vssd1 vccd1 vccd1 _7913_/CLK sky130_fd_sc_hd__inv_2
X_5470_ _8006_/Q _4347_/A _5476_/S vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4421_ _4421_/A vssd1 vssd1 vccd1 vccd1 _8218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _4352_/A vssd1 vssd1 vccd1 vccd1 _8244_/D sky130_fd_sc_hd__clkbuf_1
X_4283_ _8272_/Q _4197_/X _4285_/S vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6022_ _6009_/X _6020_/X _6021_/X _6018_/X vssd1 vssd1 vccd1 vccd1 _6022_/X sky130_fd_sc_hd__o211a_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7973_ _8441_/CLK _7973_/D vssd1 vssd1 vccd1 vccd1 _7973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6855_ _8435_/Q _6863_/B vssd1 vssd1 vccd1 vccd1 _6856_/A sky130_fd_sc_hd__and2_1
X_3998_ _4347_/A vssd1 vssd1 vccd1 vccd1 _3998_/X sky130_fd_sc_hd__buf_2
X_5806_ _5806_/A vssd1 vssd1 vccd1 vccd1 _7788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6786_ _8419_/Q _6786_/B vssd1 vssd1 vccd1 vccd1 _7478_/B sky130_fd_sc_hd__xnor2_2
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5737_ _7867_/Q _5571_/A _5737_/S vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__mux2_1
X_8456_ _8456_/CLK _8456_/D vssd1 vssd1 vccd1 vccd1 _8456_/Q sky130_fd_sc_hd__dfxtp_1
X_5668_ _5668_/A vssd1 vssd1 vccd1 vccd1 _7898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5599_ _5580_/X _7928_/Q _5599_/S vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__mux2_1
X_8387_ _8387_/CLK _8387_/D vssd1 vssd1 vccd1 vccd1 _8387_/Q sky130_fd_sc_hd__dfxtp_1
X_4619_ _4619_/A _4755_/A vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3397_ _6903_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3397_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7338_ _8083_/Q _7324_/A _7326_/X _7337_/X _7331_/X vssd1 vssd1 vccd1 vccd1 _8320_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7269_ _7282_/A _7269_/B vssd1 vssd1 vccd1 vccd1 _8298_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_31 _6108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_20 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_42 _6117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_75 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_86 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_64 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_53 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_97 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3217_ clkbuf_0__3217_/X vssd1 vssd1 vccd1 vccd1 _6488__218/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6876__398 _6876__398/A vssd1 vssd1 vccd1 vccd1 _8074_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8442_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7061__539 _7062__540/A vssd1 vssd1 vccd1 vccd1 _8220_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _4970_/A vssd1 vssd1 vccd1 vccd1 _8106_/D sky130_fd_sc_hd__clkbuf_1
X_3921_ _5502_/A _5412_/A vssd1 vssd1 vccd1 vccd1 _3944_/S sky130_fd_sc_hd__or2_2
XFILLER_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3852_ _7854_/Q vssd1 vssd1 vccd1 vccd1 _6415_/B sky130_fd_sc_hd__clkbuf_1
X_6640_ _5926_/A _7967_/Q _6640_/S vssd1 vssd1 vccd1 vccd1 _6641_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5522_ _5343_/X _7983_/Q _5530_/S vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__mux2_1
X_8310_ _8498_/CLK _8310_/D vssd1 vssd1 vccd1 vccd1 _8310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _5453_/A vssd1 vssd1 vccd1 vccd1 _8014_/D sky130_fd_sc_hd__clkbuf_1
X_8241_ _8241_/CLK _8241_/D vssd1 vssd1 vccd1 vccd1 _8241_/Q sky130_fd_sc_hd__dfxtp_1
X_8172_ _8172_/CLK _8172_/D vssd1 vssd1 vccd1 vccd1 _8172_/Q sky130_fd_sc_hd__dfxtp_1
X_5384_ _5357_/X _8048_/Q _5386_/S vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__mux2_1
X_4404_ _8067_/Q vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__buf_2
X_4335_ _4335_/A vssd1 vssd1 vccd1 vccd1 _8250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4266_ _4266_/A vssd1 vssd1 vccd1 vccd1 _8280_/D sky130_fd_sc_hd__clkbuf_1
X_6005_ _6005_/A vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__clkbuf_1
X_4197_ _8443_/Q vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2998_ clkbuf_0__2998_/X vssd1 vssd1 vccd1 vccd1 _6143__183/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7956_ _8489_/CLK _7956_/D vssd1 vssd1 vccd1 vccd1 _7956_/Q sky130_fd_sc_hd__dfxtp_1
X_7887_ _7887_/CLK _7887_/D vssd1 vssd1 vccd1 vccd1 _7887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6838_ _6844_/A vssd1 vssd1 vccd1 vccd1 _6838_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3619_ clkbuf_0__3619_/X vssd1 vssd1 vccd1 vccd1 _7396__153/A sky130_fd_sc_hd__clkbuf_4
X_8535__234 vssd1 vssd1 vccd1 vccd1 _8535__234/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6769_ _8417_/Q vssd1 vssd1 vccd1 vccd1 _6782_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8439_ _8439_/CLK _8439_/D vssd1 vssd1 vccd1 vccd1 _8439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4120_ _8130_/Q _4120_/B _4911_/B vssd1 vssd1 vccd1 vccd1 _4120_/Y sky130_fd_sc_hd__nand3_1
X_4051_ _4051_/A vssd1 vssd1 vccd1 vccd1 _8379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7810_ _8499_/CLK _7810_/D vssd1 vssd1 vccd1 vccd1 _7810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4953_ _4953_/A vssd1 vssd1 vccd1 vccd1 _8113_/D sky130_fd_sc_hd__clkbuf_1
X_8519__218 vssd1 vssd1 vccd1 vccd1 _8519__218/HI core0Index[5] sky130_fd_sc_hd__conb_1
X_7741_ _8490_/CLK _7741_/D vssd1 vssd1 vccd1 vccd1 _7741_/Q sky130_fd_sc_hd__dfxtp_1
X_3904_ _8463_/Q _3877_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7672_ _7672_/A _7704_/B vssd1 vssd1 vccd1 vccd1 _7698_/B sky130_fd_sc_hd__nand2_2
X_6263__199 _6263__199/A vssd1 vssd1 vccd1 vccd1 _7791_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4884_ _8151_/Q _4770_/X _4787_/X _8113_/Q vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1_0__3404_ clkbuf_0__3404_/X vssd1 vssd1 vccd1 vccd1 _6937__442/A sky130_fd_sc_hd__clkbuf_4
X_6623_ _6623_/A vssd1 vssd1 vccd1 vccd1 _7959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3835_ _3832_/Y _3834_/X _5316_/A vssd1 vssd1 vccd1 vccd1 _3838_/C sky130_fd_sc_hd__a21oi_1
X_5505_ _5505_/A vssd1 vssd1 vccd1 vccd1 _7991_/D sky130_fd_sc_hd__clkbuf_1
X_6485_ _6491_/A vssd1 vssd1 vccd1 vccd1 _6485_/X sky130_fd_sc_hd__buf_1
XFILLER_9_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5436_ _8024_/Q _4439_/X _5440_/S vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__mux2_1
X_8224_ _8224_/CLK _8224_/D vssd1 vssd1 vccd1 vccd1 _8224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3234_ _6572_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3234_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5367_ _5367_/A vssd1 vssd1 vccd1 vccd1 _8054_/D sky130_fd_sc_hd__clkbuf_1
X_8155_ _8155_/CLK _8155_/D vssd1 vssd1 vccd1 vccd1 _8155_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3620_ clkbuf_0__3620_/X vssd1 vssd1 vccd1 vccd1 _7404__160/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4318_ _8257_/Q _4194_/X _4322_/S vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__mux2_1
X_5298_ _8239_/Q _8247_/Q _5301_/S vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8086_ _8086_/CLK _8086_/D vssd1 vssd1 vccd1 vccd1 _8086_/Q sky130_fd_sc_hd__dfxtp_1
X_6569__283 _6569__283/A vssd1 vssd1 vccd1 vccd1 _7923_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4249_/A vssd1 vssd1 vccd1 vccd1 _8289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7253__108 _7255__110/A vssd1 vssd1 vccd1 vccd1 _8291_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7939_ _7939_/CLK _7939_/D vssd1 vssd1 vccd1 vccd1 _7939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7116__82 _7118__84/A vssd1 vssd1 vccd1 vccd1 _8263_/CLK sky130_fd_sc_hd__inv_2
X_6136__177 _6138__179/A vssd1 vssd1 vccd1 vccd1 _7726_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5221_ _8225_/Q _5046_/B _5219_/X _5220_/X vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5152_ _5152_/A _5152_/B vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__and2_1
XFILLER_102_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7432__7 _7432__7/A vssd1 vssd1 vccd1 vccd1 _8393_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7356__121 _7356__121/A vssd1 vssd1 vccd1 vccd1 _8332_/CLK sky130_fd_sc_hd__inv_2
X_4103_ _8129_/Q vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__clkbuf_2
X_5083_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _4034_/A vssd1 vssd1 vccd1 vccd1 _8386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7724_ _8017_/CLK _7724_/D vssd1 vssd1 vccd1 vccd1 _7724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _7962_/Q _5993_/B vssd1 vssd1 vccd1 vccd1 _5986_/A sky130_fd_sc_hd__and2_2
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936_ _4936_/A _5727_/A vssd1 vssd1 vccd1 vccd1 _4952_/S sky130_fd_sc_hd__nor2_2
X_4867_ _4721_/X _4857_/X _4860_/X _4866_/X _4622_/A vssd1 vssd1 vccd1 vccd1 _4867_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7655_ _8018_/Q _7701_/B vssd1 vssd1 vccd1 vccd1 _7656_/A sky130_fd_sc_hd__and2_1
X_6606_ _6606_/A _6642_/B vssd1 vssd1 vccd1 vccd1 _6622_/S sky130_fd_sc_hd__nand2_2
X_7586_ _7586_/A vssd1 vssd1 vccd1 vccd1 _7595_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _8074_/Q vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4798_ _4798_/A vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6468_ _6468_/A vssd1 vssd1 vccd1 vccd1 _6714_/S sky130_fd_sc_hd__buf_4
Xoutput150 _5921_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput161 _5942_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
X_5419_ _5419_/A vssd1 vssd1 vccd1 vccd1 _8032_/D sky130_fd_sc_hd__clkbuf_1
X_8207_ _8207_/CLK _8207_/D vssd1 vssd1 vccd1 vccd1 _8207_/Q sky130_fd_sc_hd__dfxtp_1
X_6399_ _8484_/Q _6408_/B _7672_/A vssd1 vssd1 vccd1 vccd1 _6399_/X sky130_fd_sc_hd__and3_1
Xoutput172 _5871_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3217_ _6485_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3217_/X sky130_fd_sc_hd__clkbuf_16
Xoutput194 _6110_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput183 _6076_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
X_8138_ _8138_/CLK _8138_/D vssd1 vssd1 vccd1 vccd1 _8138_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8069_ _8069_/CLK _8069_/D vssd1 vssd1 vccd1 vccd1 _8069_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3396_ clkbuf_0__3396_/X vssd1 vssd1 vccd1 vccd1 _6900__413/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6550__268 _6552__270/A vssd1 vssd1 vccd1 vccd1 _7908_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5770_ _5770_/A vssd1 vssd1 vccd1 vccd1 _7804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__buf_2
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4652_ _8332_/Q _8222_/Q _7879_/Q _8356_/Q _4650_/X _4651_/X vssd1 vssd1 vccd1 vccd1
+ _4652_/X sky130_fd_sc_hd__mux4_1
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__clkbuf_1
Xinput63 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__buf_4
Xinput41 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _5974_/A sky130_fd_sc_hd__buf_4
X_4583_ _4583_/A vssd1 vssd1 vccd1 vccd1 _8153_/D sky130_fd_sc_hd__clkbuf_1
Xinput96 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _7609_/A sky130_fd_sc_hd__buf_4
Xinput74 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _7684_/A sky130_fd_sc_hd__buf_4
Xinput85 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6322_ _6289_/X _6317_/X _6321_/X _6192_/X vssd1 vssd1 vccd1 vccd1 _6322_/X sky130_fd_sc_hd__a31o_1
X_6253_ _6259_/A vssd1 vssd1 vccd1 vccd1 _6253_/X sky130_fd_sc_hd__buf_1
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5204_ _5332_/B _5183_/X _5187_/X _5203_/X vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__a31o_1
XFILLER_97_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6184_ _6328_/A vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__clkbuf_2
X_5135_ _5187_/A _5130_/X _5132_/X _5134_/X _5159_/A vssd1 vssd1 vccd1 vccd1 _5135_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7110__77 _7110__77/A vssd1 vssd1 vccd1 vccd1 _8258_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5066_ _5084_/B _5066_/B vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4017_ _8443_/Q vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__buf_2
X_5968_ _5968_/A vssd1 vssd1 vccd1 vccd1 _5968_/X sky130_fd_sc_hd__clkbuf_1
X_4919_ _4999_/C _4921_/A _4918_/Y vssd1 vssd1 vccd1 vccd1 _8129_/D sky130_fd_sc_hd__o21a_1
X_7707_ _7707_/A _7707_/B _7707_/C vssd1 vssd1 vccd1 vccd1 _7707_/X sky130_fd_sc_hd__and3_1
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5899_ _5899_/A vssd1 vssd1 vccd1 vccd1 _5899_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7569_ _6820_/C _7564_/Y _7568_/X _7556_/X vssd1 vssd1 vccd1 vccd1 _7569_/X sky130_fd_sc_hd__a211o_1
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6881__401 _6882__402/A vssd1 vssd1 vccd1 vccd1 _8077_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6729__363 _6731__365/A vssd1 vssd1 vccd1 vccd1 _8030_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3379_ clkbuf_0__3379_/X vssd1 vssd1 vccd1 vccd1 _6872__395/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5822_ _5822_/A vssd1 vssd1 vccd1 vccd1 _7781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _7860_/Q _5568_/A _5755_/S vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3620_ _7399_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3620_/X sky130_fd_sc_hd__clkbuf_16
X_4704_ _4410_/X _4610_/X _4703_/X _4682_/X vssd1 vssd1 vccd1 vccd1 _8139_/D sky130_fd_sc_hd__o211a_1
X_8472_ _8472_/CLK _8472_/D vssd1 vssd1 vccd1 vccd1 _8472_/Q sky130_fd_sc_hd__dfxtp_1
X_5684_ _5684_/A vssd1 vssd1 vccd1 vccd1 _7891_/D sky130_fd_sc_hd__clkbuf_1
X_7423_ _7454_/A vssd1 vssd1 vccd1 vccd1 _7423_/X sky130_fd_sc_hd__buf_1
X_4635_ _4766_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__nor2_1
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _8160_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_opt_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6305_ _6296_/A _6418_/B _6310_/B vssd1 vssd1 vccd1 vccd1 _6355_/B sky130_fd_sc_hd__o21a_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4497_ _5539_/A _4936_/A vssd1 vssd1 vccd1 vccd1 _4513_/S sky130_fd_sc_hd__nor2_2
X_7285_ _7297_/A _7285_/B vssd1 vssd1 vccd1 vccd1 _8303_/D sky130_fd_sc_hd__nor2_1
X_6236_ _8320_/Q _8321_/Q _8322_/Q _8323_/Q _7317_/B _8314_/Q vssd1 vssd1 vccd1 vccd1
+ _6236_/X sky130_fd_sc_hd__mux4_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _7678_/A vssd1 vssd1 vccd1 vccd1 _6167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _3925_/X _5022_/X _5117_/X _5091_/X vssd1 vssd1 vccd1 vccd1 _8085_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6098_ _7829_/Q _6129_/C _7703_/A vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__a21bo_2
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5049_ _5196_/S vssd1 vssd1 vccd1 vccd1 _5190_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3233_ clkbuf_0__3233_/X vssd1 vssd1 vccd1 vccd1 _6569__283/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7369__131 _7370__132/A vssd1 vssd1 vccd1 vccd1 _8342_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7625__34 _7626__35/A vssd1 vssd1 vccd1 vccd1 _8457_/CLK sky130_fd_sc_hd__inv_2
X_6662__314 _6663__315/A vssd1 vssd1 vccd1 vccd1 _7978_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6888__407 _6891__410/A vssd1 vssd1 vccd1 vccd1 _8083_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4420_ _4419_/X _8218_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6968__464 _6968__464/A vssd1 vssd1 vccd1 vccd1 _8145_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4351_ _4350_/X _8244_/Q _4357_/S vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4282_ _4282_/A vssd1 vssd1 vccd1 vccd1 _8273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6021_ _7734_/Q _6025_/B vssd1 vssd1 vccd1 vccd1 _6021_/X sky130_fd_sc_hd__or2_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7972_ _8439_/CLK _7972_/D vssd1 vssd1 vccd1 vccd1 _7972_/Q sky130_fd_sc_hd__dfxtp_1
X_6563__278 _6563__278/A vssd1 vssd1 vccd1 vccd1 _7918_/CLK sky130_fd_sc_hd__inv_2
X_6923_ _6942_/A vssd1 vssd1 vccd1 vccd1 _6923_/X sky130_fd_sc_hd__buf_1
XFILLER_23_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6854_ _6854_/A vssd1 vssd1 vccd1 vccd1 _6863_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3997_ _8448_/Q vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__buf_2
X_5805_ _3880_/X _7788_/Q _5807_/S vssd1 vssd1 vccd1 vccd1 _5806_/A sky130_fd_sc_hd__mux2_1
X_6785_ _7200_/A _6785_/B vssd1 vssd1 vccd1 vccd1 _6785_/X sky130_fd_sc_hd__xor2_1
X_5736_ _5736_/A vssd1 vssd1 vccd1 vccd1 _7868_/D sky130_fd_sc_hd__clkbuf_1
X_5667_ _5574_/X _7898_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5668_/A sky130_fd_sc_hd__mux2_1
X_8455_ _8455_/CLK _8455_/D vssd1 vssd1 vccd1 vccd1 _8455_/Q sky130_fd_sc_hd__dfxtp_1
X_4618_ _4623_/B vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__clkbuf_2
X_5598_ _5598_/A vssd1 vssd1 vccd1 vccd1 _7929_/D sky130_fd_sc_hd__clkbuf_1
X_8386_ _8386_/CLK _8386_/D vssd1 vssd1 vccd1 vccd1 _8386_/Q sky130_fd_sc_hd__dfxtp_1
X_4549_ _8167_/Q _4454_/X _4549_/S vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__mux2_1
X_7337_ _8320_/Q _7337_/B vssd1 vssd1 vccd1 vccd1 _7337_/X sky130_fd_sc_hd__or2_1
Xclkbuf_0__3396_ _6897_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3396_/X sky130_fd_sc_hd__clkbuf_16
X_7268_ _7261_/B _7206_/B _7262_/Y _7264_/X _8298_/Q vssd1 vssd1 vccd1 vccd1 _7269_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6219_ _7611_/A _7770_/Q _6223_/S vssd1 vssd1 vccd1 vccd1 _6220_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7199_ _8300_/Q _7273_/A vssd1 vssd1 vccd1 vccd1 _7200_/B sky130_fd_sc_hd__xor2_1
XINSDIODE2_10 _7703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_43 _6117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_32 _6108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_21 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_54 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_76 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_65 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_98 _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_87 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7350__116 _7351__117/A vssd1 vssd1 vccd1 vccd1 _8327_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3949_/A _3920_/B _4025_/B _3948_/A vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__or4b_2
X_3851_ _7833_/Q _7834_/Q _6301_/B vssd1 vssd1 vccd1 vccd1 _7654_/A sky130_fd_sc_hd__or3_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5521_ _5536_/S vssd1 vssd1 vccd1 vccd1 _5530_/S sky130_fd_sc_hd__buf_2
X_8240_ _8240_/CLK _8240_/D vssd1 vssd1 vccd1 vccd1 _8240_/Q sky130_fd_sc_hd__dfxtp_1
X_5452_ _8014_/Q _4436_/X _5458_/S vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__mux2_1
X_8171_ _8171_/CLK _8171_/D vssd1 vssd1 vccd1 vccd1 _8171_/Q sky130_fd_sc_hd__dfxtp_1
X_5383_ _5383_/A vssd1 vssd1 vccd1 vccd1 _8049_/D sky130_fd_sc_hd__clkbuf_1
X_4403_ _4403_/A vssd1 vssd1 vccd1 vccd1 _8223_/D sky130_fd_sc_hd__clkbuf_1
X_4334_ _8250_/Q _4191_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6004_ _7970_/Q _6006_/B vssd1 vssd1 vccd1 vccd1 _6005_/A sky130_fd_sc_hd__and2_1
X_4265_ _8280_/Q _4197_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__mux2_1
X_4196_ _4196_/A vssd1 vssd1 vccd1 vccd1 _8335_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2997_ clkbuf_0__2997_/X vssd1 vssd1 vccd1 vccd1 _6139__180/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7955_ _8490_/CLK _7955_/D vssd1 vssd1 vccd1 vccd1 _7955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7886_ _7886_/CLK _7886_/D vssd1 vssd1 vccd1 vccd1 _7886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3618_ clkbuf_0__3618_/X vssd1 vssd1 vccd1 vccd1 _7411_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3549_ clkbuf_0__3549_/X vssd1 vssd1 vccd1 vccd1 _7255__110/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6768_ _6768_/A _7471_/B _7471_/C vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__and3_1
X_6275__208 _6275__208/A vssd1 vssd1 vccd1 vccd1 _7800_/CLK sky130_fd_sc_hd__inv_2
X_5719_ _4147_/X _7875_/Q _5719_/S vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__mux2_1
X_8438_ _8439_/CLK _8438_/D vssd1 vssd1 vccd1 vccd1 _8438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8369_ _8369_/CLK _8369_/D vssd1 vssd1 vccd1 vccd1 _8369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3379_ _6850_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3379_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7414__168 _7414__168/A vssd1 vssd1 vccd1 vccd1 _8379_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6514__239 _6514__239/A vssd1 vssd1 vccd1 vccd1 _7879_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ _8379_/Q _3998_/X _4056_/S vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037__520 _7037__520/A vssd1 vssd1 vccd1 vccd1 _8201_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _8113_/Q _4247_/X _4952_/S vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__mux2_1
X_7740_ _8490_/CLK _7740_/D vssd1 vssd1 vccd1 vccd1 _7740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _8464_/D sky130_fd_sc_hd__clkbuf_1
X_4883_ _4883_/A _4883_/B _4883_/C vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__or3_1
X_7671_ _8483_/Q _7656_/X _7670_/X _7662_/X vssd1 vssd1 vccd1 vccd1 _8483_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6622_ _7677_/A _7959_/Q _6622_/S vssd1 vssd1 vccd1 vccd1 _6623_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3834_ _8074_/Q _3920_/B _5018_/A vssd1 vssd1 vccd1 vccd1 _3834_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0__3403_ clkbuf_0__3403_/X vssd1 vssd1 vccd1 vccd1 _6934__440/A sky130_fd_sc_hd__clkbuf_4
X_6553_ _6553_/A vssd1 vssd1 vccd1 vccd1 _6553_/X sky130_fd_sc_hd__buf_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5504_ _7991_/Q _4342_/A _5512_/S vssd1 vssd1 vccd1 vccd1 _5505_/A sky130_fd_sc_hd__mux2_1
X_6484_ _6149_/X _6231_/B _7649_/A vssd1 vssd1 vccd1 vccd1 _7855_/D sky130_fd_sc_hd__a21oi_1
X_5435_ _5435_/A vssd1 vssd1 vccd1 vccd1 _8025_/D sky130_fd_sc_hd__clkbuf_1
X_8223_ _8223_/CLK _8223_/D vssd1 vssd1 vccd1 vccd1 _8223_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3233_ _6566_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3233_/X sky130_fd_sc_hd__clkbuf_16
X_7142__103 _7144__105/A vssd1 vssd1 vccd1 vccd1 _8284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5366_ _5365_/X _8054_/Q _5374_/S vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__mux2_1
X_8154_ _8154_/CLK _8154_/D vssd1 vssd1 vccd1 vccd1 _8154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4317_ _4317_/A vssd1 vssd1 vccd1 vccd1 _8258_/D sky130_fd_sc_hd__clkbuf_1
X_5297_ _5048_/X _5293_/X _5295_/X _5296_/X _5056_/X vssd1 vssd1 vccd1 vccd1 _5297_/X
+ sky130_fd_sc_hd__a221o_1
X_8085_ _8085_/CLK _8085_/D vssd1 vssd1 vccd1 vccd1 _8085_/Q sky130_fd_sc_hd__dfxtp_1
X_4248_ _8289_/Q _4247_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6723__358 _6723__358/A vssd1 vssd1 vccd1 vccd1 _8025_/CLK sky130_fd_sc_hd__inv_2
X_4179_ _4201_/S vssd1 vssd1 vccd1 vccd1 _4192_/S sky130_fd_sc_hd__buf_2
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7938_ _7938_/CLK _7938_/D vssd1 vssd1 vccd1 vccd1 _7938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7869_ _7869_/CLK _7869_/D vssd1 vssd1 vccd1 vccd1 _7869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5220_/A vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5151_ _8470_/Q _8211_/Q _8203_/Q _8235_/Q _5060_/A _5044_/A vssd1 vssd1 vccd1 vccd1
+ _5152_/B sky130_fd_sc_hd__mux4_1
X_5082_ _5079_/X _5081_/X _5152_/A vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _8130_/Q vssd1 vssd1 vccd1 vccd1 _4475_/B sky130_fd_sc_hd__clkbuf_2
X_4033_ _8386_/Q _4002_/X _4037_/S vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__mux2_1
X_6826__371 _6827__372/A vssd1 vssd1 vccd1 vccd1 _8039_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5993_/B sky130_fd_sc_hd__clkbuf_4
X_7723_ _7723_/A vssd1 vssd1 vccd1 vccd1 _8499_/D sky130_fd_sc_hd__clkbuf_1
X_4935_ _4630_/X _4924_/X _4934_/Y vssd1 vssd1 vccd1 vccd1 _8122_/D sky130_fd_sc_hd__a21oi_1
X_4866_ _4861_/X _4862_/X _4773_/A _4865_/X vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__a211o_1
X_7654_ _7654_/A _7654_/B _7654_/C _7654_/D vssd1 vssd1 vccd1 vccd1 _7701_/B sky130_fd_sc_hd__nor4_4
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4797_ _8218_/Q _4795_/X _4796_/X _7875_/Q vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__a22o_1
X_3817_ _4287_/A _5319_/A _3972_/B vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__or3_2
X_7585_ _8437_/Q _7578_/X _7584_/X _7582_/X vssd1 vssd1 vccd1 vccd1 _8436_/D sky130_fd_sc_hd__o211a_1
X_7363__126 _7367__130/A vssd1 vssd1 vccd1 vccd1 _8337_/CLK sky130_fd_sc_hd__inv_2
X_6467_ _6467_/A vssd1 vssd1 vccd1 vccd1 _7850_/D sky130_fd_sc_hd__clkbuf_1
Xoutput151 _5923_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
X_8206_ _8206_/CLK _8206_/D vssd1 vssd1 vccd1 vccd1 _8206_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput140 _5901_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
X_5418_ _3877_/X _8032_/Q _5422_/S vssd1 vssd1 vccd1 vccd1 _5419_/A sky130_fd_sc_hd__mux2_1
X_6398_ _7822_/Q _6383_/X _6393_/X _6397_/X _6391_/X vssd1 vssd1 vccd1 vccd1 _7822_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput162 _5944_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput173 _5873_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
X_5349_ _5562_/A vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__clkbuf_2
Xoutput184 _6079_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput195 _6114_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8137_ _8137_/CLK _8137_/D vssd1 vssd1 vccd1 vccd1 _8137_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8068_ _8068_/CLK _8068_/D vssd1 vssd1 vccd1 vccd1 _8068_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6142__182 _6143__183/A vssd1 vssd1 vccd1 vccd1 _7731_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4720_ _4718_/X _4719_/X _4740_/S vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__mux2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4651_ _4670_/A vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__buf_2
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__clkbuf_4
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
Xinput53 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _3846_/D sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__buf_4
Xinput42 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__buf_4
X_4582_ _4422_/X _8153_/Q _4586_/S vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput75 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _7681_/A sky130_fd_sc_hd__buf_4
Xinput86 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _5928_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput97 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _7611_/A sky130_fd_sc_hd__buf_4
X_6321_ _8474_/Q _6311_/X _6320_/X _6306_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _6321_/X
+ sky130_fd_sc_hd__a221o_1
X_5203_ _5187_/A _5192_/X _5195_/X _5202_/X _5031_/A vssd1 vssd1 vccd1 vccd1 _5203_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6183_ _6176_/X _7961_/Q _6178_/X _6180_/X _7750_/Q vssd1 vssd1 vccd1 vccd1 _7750_/D
+ sky130_fd_sc_hd__o32a_1
X_5134_ _5038_/A _5133_/X _5113_/X vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _8396_/Q _8388_/Q _7791_/Q _8404_/Q _5063_/X _5064_/X vssd1 vssd1 vccd1 vccd1
+ _5065_/X sky130_fd_sc_hd__mux4_1
X_4016_ _4016_/A vssd1 vssd1 vccd1 vccd1 _8391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5967_ _5967_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5968_/A sky130_fd_sc_hd__and2_1
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7706_ _6359_/X _7707_/C _7705_/X _6421_/X vssd1 vssd1 vccd1 vccd1 _8492_/D sky130_fd_sc_hd__o211a_1
X_4918_ _4911_/B _4911_/C _6963_/C vssd1 vssd1 vccd1 vccd1 _4918_/Y sky130_fd_sc_hd__a21boi_1
X_5898_ _7693_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__or2_1
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4849_ _4753_/X _8053_/Q _7937_/Q _4796_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _4849_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7568_ _8432_/Q _7563_/A _7567_/Y vssd1 vssd1 vccd1 vccd1 _7568_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7499_ _7499_/A _7499_/B _7499_/C vssd1 vssd1 vccd1 vccd1 _7500_/D sky130_fd_sc_hd__and3_1
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3378_ clkbuf_0__3378_/X vssd1 vssd1 vccd1 vccd1 _6846__387/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5821_ _7781_/Q _5565_/A _5825_/S vssd1 vssd1 vccd1 vccd1 _5822_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5752_ _5752_/A vssd1 vssd1 vccd1 vccd1 _7861_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3550_ _7256_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3550_/X sky130_fd_sc_hd__clkbuf_16
X_4703_ _4612_/X _8139_/Q _4924_/A _4702_/X _4678_/X vssd1 vssd1 vccd1 vccd1 _4703_/X
+ sky130_fd_sc_hd__a221o_1
X_8471_ _8471_/CLK _8471_/D vssd1 vssd1 vccd1 vccd1 _8471_/Q sky130_fd_sc_hd__dfxtp_1
X_5683_ _7891_/Q _4987_/X _5683_/S vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4634_ _8051_/Q _8043_/Q _7871_/Q _8112_/Q _4630_/X _4633_/X vssd1 vssd1 vccd1 vccd1
+ _4634_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4565_ _4425_/X _8160_/Q _4567_/S vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6304_ _6304_/A _7654_/A _6304_/C _6297_/B vssd1 vssd1 vccd1 vccd1 _6310_/B sky130_fd_sc_hd__or4b_1
XFILLER_89_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4496_ _4475_/B _4999_/C _4999_/A vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__nand3b_2
X_7284_ _8303_/Q _7280_/X _7272_/X _7192_/B vssd1 vssd1 vccd1 vccd1 _7285_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _8313_/Q vssd1 vssd1 vccd1 vccd1 _7317_/B sky130_fd_sc_hd__clkbuf_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6159_/X _7772_/Q _6161_/X _6163_/X _7740_/Q vssd1 vssd1 vccd1 vccd1 _7740_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6473_/A vssd1 vssd1 vccd1 vccd1 _7703_/A sky130_fd_sc_hd__clkbuf_4
X_5117_ _8085_/Q _5024_/X _5331_/A _5116_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5117_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5048_ _5062_/A vssd1 vssd1 vccd1 vccd1 _5048_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3232_ clkbuf_0__3232_/X vssd1 vssd1 vccd1 vccd1 _6565__280/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6839__381 _6841__383/A vssd1 vssd1 vccd1 vccd1 _8049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7031__515 _7031__515/A vssd1 vssd1 vccd1 vccd1 _8196_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4350_/A vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4281_ _8273_/Q _4194_/X _4285_/S vssd1 vssd1 vccd1 vccd1 _4282_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _7809_/Q input14/X _6123_/B vssd1 vssd1 vccd1 vccd1 _6020_/X sky130_fd_sc_hd__mux2_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7971_ _8439_/CLK _7971_/D vssd1 vssd1 vccd1 vccd1 _7971_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6853_ _6853_/A vssd1 vssd1 vccd1 vccd1 _8060_/D sky130_fd_sc_hd__clkbuf_1
X_5804_ _5804_/A vssd1 vssd1 vccd1 vccd1 _7789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3996_ _3996_/A vssd1 vssd1 vccd1 vccd1 _8396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6784_ _7479_/B _7479_/C vssd1 vssd1 vccd1 vccd1 _6785_/B sky130_fd_sc_hd__nand2_1
X_5735_ _7868_/Q _5568_/A _5737_/S vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5666_ _5666_/A vssd1 vssd1 vccd1 vccd1 _7899_/D sky130_fd_sc_hd__clkbuf_1
X_8454_ _8454_/CLK _8454_/D vssd1 vssd1 vccd1 vccd1 _8454_/Q sky130_fd_sc_hd__dfxtp_1
X_4617_ _8123_/Q _8122_/Q vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__nand2_1
X_7405_ _7417_/A vssd1 vssd1 vccd1 vccd1 _7405_/X sky130_fd_sc_hd__buf_1
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5597_ _5577_/X _7929_/Q _5599_/S vssd1 vssd1 vccd1 vccd1 _5598_/A sky130_fd_sc_hd__mux2_1
X_8385_ _8385_/CLK _8385_/D vssd1 vssd1 vccd1 vccd1 _8385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4548_ _4548_/A vssd1 vssd1 vccd1 vccd1 _8168_/D sky130_fd_sc_hd__clkbuf_1
X_7336_ _8082_/Q _7648_/B _7326_/X _7335_/X _7331_/X vssd1 vssd1 vccd1 vccd1 _8319_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_116_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _4479_/A vssd1 vssd1 vccd1 vccd1 _8198_/D sky130_fd_sc_hd__clkbuf_1
X_7267_ _7321_/A vssd1 vssd1 vccd1 vccd1 _7282_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6218_ _6218_/A vssd1 vssd1 vccd1 vccd1 _7769_/D sky130_fd_sc_hd__clkbuf_1
X_7198_ _8299_/Q _8298_/Q _8297_/Q vssd1 vssd1 vccd1 vccd1 _7273_/A sky130_fd_sc_hd__nand3_2
XINSDIODE2_22 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6149_ _6161_/A vssd1 vssd1 vccd1 vccd1 _6149_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_33 _6113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_11 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_44 _6117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_66 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_77 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_55 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_88 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_99 _5943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _7835_/Q _7836_/Q _7837_/Q _7838_/Q vssd1 vssd1 vccd1 vccd1 _6301_/B sky130_fd_sc_hd__or4_1
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5520_ _5655_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5536_/S sky130_fd_sc_hd__or2_2
XFILLER_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5451_ _5451_/A vssd1 vssd1 vccd1 vccd1 _8015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8170_ _8170_/CLK _8170_/D vssd1 vssd1 vccd1 vccd1 _8170_/Q sky130_fd_sc_hd__dfxtp_1
X_5382_ _5353_/X _8049_/Q _5386_/S vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__mux2_1
X_4402_ _4365_/X _8223_/Q _4402_/S vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__mux2_1
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _8251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4264_ _4264_/A vssd1 vssd1 vccd1 vccd1 _8281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6003_ _6003_/A vssd1 vssd1 vccd1 vccd1 _6003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4195_ _8335_/Q _4194_/X _4201_/S vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2996_ clkbuf_0__2996_/X vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__clkbuf_4
X_7954_ _8490_/CLK _7954_/D vssd1 vssd1 vccd1 vccd1 _7954_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7885_ _7885_/CLK _7885_/D vssd1 vssd1 vccd1 vccd1 _7885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3617_ clkbuf_0__3617_/X vssd1 vssd1 vccd1 vccd1 _7391__150/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6767_ _7471_/B _7471_/C _6768_/A vssd1 vssd1 vccd1 vccd1 _6767_/Y sky130_fd_sc_hd__a21oi_1
X_3979_ _3928_/X _8402_/Q _3983_/S vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__mux2_1
X_5718_ _5718_/A vssd1 vssd1 vccd1 vccd1 _7876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _5574_/X _7906_/Q _5653_/S vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__mux2_1
X_7128__92 _7128__92/A vssd1 vssd1 vccd1 vccd1 _8273_/CLK sky130_fd_sc_hd__inv_2
X_8437_ _8439_/CLK _8437_/D vssd1 vssd1 vccd1 vccd1 _8437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8368_ _8368_/CLK _8368_/D vssd1 vssd1 vccd1 vccd1 _8368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7319_ _8314_/Q _7315_/Y _7318_/X _7248_/X vssd1 vssd1 vccd1 vccd1 _8314_/D sky130_fd_sc_hd__o211a_1
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3378_ _6844_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3378_/X sky130_fd_sc_hd__clkbuf_16
X_8299_ _8315_/CLK _8299_/D vssd1 vssd1 vccd1 vccd1 _8299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6709__351 _6719__355/A vssd1 vssd1 vccd1 vccd1 _8015_/CLK sky130_fd_sc_hd__inv_2
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7002__491 _7004__493/A vssd1 vssd1 vccd1 vccd1 _8172_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4951_ _4951_/A vssd1 vssd1 vccd1 vccd1 _8114_/D sky130_fd_sc_hd__clkbuf_1
X_3902_ _8464_/Q _3874_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__mux2_1
X_4882_ _4783_/X _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _4883_/C sky130_fd_sc_hd__o21a_1
X_7670_ _5911_/A _7657_/X _7660_/Y vssd1 vssd1 vccd1 vccd1 _7670_/X sky130_fd_sc_hd__a21o_1
X_6675__325 _6675__325/A vssd1 vssd1 vccd1 vccd1 _7989_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3402_ clkbuf_0__3402_/X vssd1 vssd1 vccd1 vccd1 _6926__433/A sky130_fd_sc_hd__clkbuf_4
X_3833_ _8075_/Q _8070_/Q vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__xnor2_1
X_6621_ _6621_/A vssd1 vssd1 vccd1 vccd1 _7958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5503_ _5518_/S vssd1 vssd1 vccd1 vccd1 _5512_/S sky130_fd_sc_hd__buf_2
X_6483_ _7722_/A vssd1 vssd1 vccd1 vccd1 _7649_/A sky130_fd_sc_hd__clkbuf_4
X_5434_ _8025_/Q _4436_/X _5440_/S vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__mux2_1
X_8222_ _8222_/CLK _8222_/D vssd1 vssd1 vccd1 vccd1 _8222_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3232_ _6560_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3232_/X sky130_fd_sc_hd__clkbuf_16
X_8153_ _8153_/CLK _8153_/D vssd1 vssd1 vccd1 vccd1 _8153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5365_ _5574_/A vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4316_ _8258_/Q _4191_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__mux2_1
X_5296_ _5214_/A _8027_/Q _7792_/Q _5239_/B _5074_/X vssd1 vssd1 vccd1 vccd1 _5296_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8084_ _8084_/CLK _8084_/D vssd1 vssd1 vccd1 vccd1 _8084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4247_ _8060_/Q vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8541__240 vssd1 vssd1 vccd1 vccd1 _8541__240/HI partID[3] sky130_fd_sc_hd__conb_1
X_4178_ _5502_/B _4178_/B vssd1 vssd1 vccd1 vccd1 _4201_/S sky130_fd_sc_hd__nor2_2
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7937_ _7937_/CLK _7937_/D vssd1 vssd1 vccd1 vccd1 _7937_/Q sky130_fd_sc_hd__dfxtp_1
X_6281__213 _6282__214/A vssd1 vssd1 vccd1 vccd1 _7805_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _7868_/CLK _7868_/D vssd1 vssd1 vccd1 vccd1 _7868_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6819_ _6819_/A vssd1 vssd1 vccd1 vccd1 _6820_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7799_ _7799_/CLK _7799_/D vssd1 vssd1 vccd1 vccd1 _7799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6576__289 _6577__290/A vssd1 vssd1 vccd1 vccd1 _7929_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7420__173 _7422__175/A vssd1 vssd1 vccd1 vccd1 _8384_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6520__244 _6521__245/A vssd1 vssd1 vccd1 vccd1 _7884_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5150_ _5148_/X _5149_/X _5186_/S vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__mux2_1
X_8525__224 vssd1 vssd1 vccd1 vccd1 _8525__224/HI core1Index[4] sky130_fd_sc_hd__conb_1
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5081_ _8380_/Q _8278_/Q _8015_/Q _8230_/Q _5064_/A _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5081_/X sky130_fd_sc_hd__mux4_1
X_7122__87 _7123__88/A vssd1 vssd1 vccd1 vccd1 _8268_/CLK sky130_fd_sc_hd__inv_2
X_4101_ _8067_/Q vssd1 vssd1 vccd1 vccd1 _4101_/X sky130_fd_sc_hd__buf_2
XFILLER_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4032_ _4032_/A vssd1 vssd1 vccd1 vccd1 _8387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7440__14 _7441__15/A vssd1 vssd1 vccd1 vccd1 _8400_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5983_ _5983_/A vssd1 vssd1 vccd1 vccd1 _5983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7722_ _7722_/A _7722_/B vssd1 vssd1 vccd1 vccd1 _7723_/A sky130_fd_sc_hd__or2_1
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4934_ _4630_/X _4932_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _4934_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_19_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4865_ _8045_/Q _4814_/X _4798_/X _4864_/X vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__o211a_1
X_7653_ _7832_/Q _7658_/A _6292_/B vssd1 vssd1 vccd1 vccd1 _7654_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6604_ _6670_/A vssd1 vssd1 vccd1 vccd1 _6604_/X sky130_fd_sc_hd__buf_1
X_4796_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4796_/X sky130_fd_sc_hd__buf_2
X_3816_ _8075_/Q vssd1 vssd1 vccd1 vccd1 _3972_/B sky130_fd_sc_hd__clkbuf_1
X_7584_ _8436_/Q _7584_/B vssd1 vssd1 vccd1 vccd1 _7584_/X sky130_fd_sc_hd__or2_1
XFILLER_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6535_ _6547_/A vssd1 vssd1 vccd1 vccd1 _6535_/X sky130_fd_sc_hd__buf_1
X_6833__376 _6836__379/A vssd1 vssd1 vccd1 vccd1 _8044_/CLK sky130_fd_sc_hd__inv_2
X_8205_ _8205_/CLK _8205_/D vssd1 vssd1 vccd1 vccd1 _8205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6466_ _7850_/Q _7965_/Q _6466_/S vssd1 vssd1 vccd1 vccd1 _6467_/A sky130_fd_sc_hd__mux2_1
Xoutput152 _5925_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput130 _5953_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput141 _5903_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
X_5417_ _5417_/A vssd1 vssd1 vccd1 vccd1 _8033_/D sky130_fd_sc_hd__clkbuf_1
X_6397_ _7680_/A _6408_/B _7672_/A vssd1 vssd1 vccd1 vccd1 _6397_/X sky130_fd_sc_hd__and3_1
Xoutput174 _5861_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput163 _5883_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
X_5348_ _8066_/Q vssd1 vssd1 vccd1 vccd1 _5562_/A sky130_fd_sc_hd__buf_2
Xoutput185 _6083_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8136_ _8136_/CLK _8136_/D vssd1 vssd1 vccd1 vccd1 _8136_/Q sky130_fd_sc_hd__dfxtp_1
X_7009__497 _7009__497/A vssd1 vssd1 vccd1 vccd1 _8178_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput196 _6116_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
X_8067_ _8439_/CLK _8067_/D vssd1 vssd1 vccd1 vccd1 _8067_/Q sky130_fd_sc_hd__dfxtp_2
X_5279_ _5334_/B _5268_/Y _5271_/Y _5278_/X _5332_/B vssd1 vssd1 vccd1 vccd1 _5280_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_56_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6246__185 _6246__185/A vssd1 vssd1 vccd1 vccd1 _7777_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4650_ _4650_/A vssd1 vssd1 vccd1 vccd1 _4650_/X sky130_fd_sc_hd__clkbuf_4
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _6113_/A sky130_fd_sc_hd__clkbuf_4
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
Xinput54 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _3846_/C sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _6012_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6320_ _8134_/Q _6318_/X _6319_/X vssd1 vssd1 vccd1 vccd1 _6320_/X sky130_fd_sc_hd__a21o_1
X_4581_ _4581_/A vssd1 vssd1 vccd1 vccd1 _8154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput98 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _7707_/A sky130_fd_sc_hd__buf_4
Xinput65 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _5958_/A sky130_fd_sc_hd__buf_4
Xinput76 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _7677_/A sky130_fd_sc_hd__clkbuf_2
Xinput87 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__buf_4
XFILLER_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5202_ _5202_/A _5202_/B _5202_/C vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__or3_1
X_6182_ _6176_/X _7960_/Q _6178_/X _6180_/X _7749_/Q vssd1 vssd1 vccd1 vccd1 _7749_/D
+ sky130_fd_sc_hd__o32a_1
X_5133_ _8172_/Q _8148_/Q _8410_/Q _8180_/Q _5123_/A _5111_/X vssd1 vssd1 vccd1 vccd1
+ _5133_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5064_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5064_/X sky130_fd_sc_hd__buf_2
XFILLER_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4015_ _8391_/Q _4014_/X _4023_/S vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__clkbuf_1
X_5897_ _5943_/B vssd1 vssd1 vccd1 vccd1 _5906_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7705_ _7615_/A _7707_/B _7704_/Y vssd1 vssd1 vccd1 vccd1 _7705_/X sky130_fd_sc_hd__a21o_1
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _8130_/D sky130_fd_sc_hd__clkbuf_1
X_4848_ _4843_/X _4844_/X _4847_/X _4928_/B vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__a211o_1
X_4779_ _8292_/Q _4778_/X _8100_/Q _4762_/X _4696_/S vssd1 vssd1 vccd1 vccd1 _4779_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7567_ _8432_/Q _7563_/A _7577_/A vssd1 vssd1 vccd1 vccd1 _7567_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7498_ _7683_/A _7498_/B vssd1 vssd1 vccd1 vccd1 _7499_/C sky130_fd_sc_hd__xor2_1
XFILLER_106_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6688__335 _6688__335/A vssd1 vssd1 vccd1 vccd1 _7999_/CLK sky130_fd_sc_hd__inv_2
X_6449_ _7842_/Q _5974_/A _6455_/S vssd1 vssd1 vccd1 vccd1 _6450_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7637__44 _7638__45/A vssd1 vssd1 vccd1 vccd1 _8467_/CLK sky130_fd_sc_hd__inv_2
X_8119_ _8119_/CLK _8119_/D vssd1 vssd1 vccd1 vccd1 _8119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3377_ clkbuf_0__3377_/X vssd1 vssd1 vccd1 vccd1 _6843__385/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5820_ _5820_/A vssd1 vssd1 vccd1 vccd1 _7782_/D sky130_fd_sc_hd__clkbuf_1
X_5751_ _7861_/Q _5565_/A _5755_/S vssd1 vssd1 vccd1 vccd1 _5752_/A sky130_fd_sc_hd__mux2_1
X_8470_ _8470_/CLK _8470_/D vssd1 vssd1 vccd1 vccd1 _8470_/Q sky130_fd_sc_hd__dfxtp_1
X_4702_ _4622_/X _4687_/X _4691_/X _4701_/X vssd1 vssd1 vccd1 vccd1 _4702_/X sky130_fd_sc_hd__a31o_1
X_5682_ _5682_/A vssd1 vssd1 vccd1 vccd1 _7892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _4633_/A vssd1 vssd1 vccd1 vccd1 _4633_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4564_ _4564_/A vssd1 vssd1 vccd1 vccd1 _8161_/D sky130_fd_sc_hd__clkbuf_1
X_6533__254 _6534__255/A vssd1 vssd1 vccd1 vccd1 _7894_/CLK sky130_fd_sc_hd__inv_2
X_7283_ _7321_/A vssd1 vssd1 vccd1 vccd1 _7297_/A sky130_fd_sc_hd__clkbuf_2
X_6303_ _7832_/Q vssd1 vssd1 vccd1 vccd1 _6304_/A sky130_fd_sc_hd__clkinv_2
XFILLER_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6234_ _8288_/Q vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__clkbuf_2
X_4495_ _5538_/A vssd1 vssd1 vccd1 vccd1 _4999_/A sky130_fd_sc_hd__buf_2
XFILLER_69_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6159_/X _7771_/Q _6161_/X _6163_/X _7739_/Q vssd1 vssd1 vccd1 vccd1 _7739_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _5031_/X _5097_/X _5103_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__a31o_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6096_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6096_/X sky130_fd_sc_hd__and2_1
X_5047_ _5108_/A vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3231_ clkbuf_0__3231_/X vssd1 vssd1 vccd1 vccd1 _6584_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5949_ _5949_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__and2_1
XFILLER_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7376__137 _7376__137/A vssd1 vssd1 vccd1 vccd1 _8348_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3429_ clkbuf_0__3429_/X vssd1 vssd1 vccd1 vccd1 _7068__545/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3444_ clkbuf_0__3444_/X vssd1 vssd1 vccd1 vccd1 _7349_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4280_ _4280_/A vssd1 vssd1 vccd1 vccd1 _8274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7631__39 _7632__40/A vssd1 vssd1 vccd1 vccd1 _8462_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7970_ _8439_/CLK _7970_/D vssd1 vssd1 vccd1 vccd1 _7970_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6852_ _8434_/Q _6852_/B vssd1 vssd1 vccd1 vccd1 _6853_/A sky130_fd_sc_hd__and2_1
X_5803_ _3877_/X _7789_/Q _5807_/S vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3995_ _8396_/Q _3992_/X _4011_/S vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6783_ _6782_/B _6782_/C _7473_/B _8418_/Q vssd1 vssd1 vccd1 vccd1 _7479_/C sky130_fd_sc_hd__a31o_1
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _5734_/A vssd1 vssd1 vccd1 vccd1 _7869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5665_ _5571_/X _7899_/Q _5665_/S vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__mux2_1
X_8453_ _8453_/CLK _8453_/D vssd1 vssd1 vccd1 vccd1 _8453_/Q sky130_fd_sc_hd__dfxtp_1
X_8384_ _8384_/CLK _8384_/D vssd1 vssd1 vccd1 vccd1 _8384_/Q sky130_fd_sc_hd__dfxtp_1
X_4616_ _4623_/A vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__clkbuf_2
X_5596_ _5596_/A vssd1 vssd1 vccd1 vccd1 _7930_/D sky130_fd_sc_hd__clkbuf_1
X_7335_ _8319_/Q _7337_/B vssd1 vssd1 vccd1 vccd1 _7335_/X sky130_fd_sc_hd__or2_1
X_4547_ _8168_/Q _4451_/X _4549_/S vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__mux2_1
X_4478_ _8198_/Q _4223_/X _4486_/S vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__mux2_1
X_7266_ _7208_/B _7262_/Y _7265_/Y _7248_/X vssd1 vssd1 vccd1 vccd1 _8297_/D sky130_fd_sc_hd__o211a_1
XFILLER_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6217_ _7609_/A _7769_/Q _6217_/S vssd1 vssd1 vccd1 vccd1 _6218_/A sky130_fd_sc_hd__mux2_1
X_7197_ _7197_/A _7197_/B vssd1 vssd1 vccd1 vccd1 _7197_/X sky130_fd_sc_hd__xor2_1
X_6148_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__buf_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8505__255 vssd1 vssd1 vccd1 vccd1 partID[8] _8505__255/LO sky130_fd_sc_hd__conb_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_12 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _6113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_67 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_56 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6072_/X _6077_/X _6078_/X _6075_/X vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__o211a_1
XINSDIODE2_45 _6119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_89 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_78 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3280_ clkbuf_0__3280_/X vssd1 vssd1 vccd1 vccd1 _6825_/A sky130_fd_sc_hd__clkbuf_4
X_5450_ _8015_/Q _4431_/X _5458_/S vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4401_ _4401_/A vssd1 vssd1 vccd1 vccd1 _8224_/D sky130_fd_sc_hd__clkbuf_1
X_5381_ _5381_/A vssd1 vssd1 vccd1 vccd1 _8050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4332_ _8251_/Q _4188_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__mux2_1
X_7120_ _7120_/A vssd1 vssd1 vccd1 vccd1 _7120_/X sky130_fd_sc_hd__buf_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7051_ _7057_/A vssd1 vssd1 vccd1 vccd1 _7051_/X sky130_fd_sc_hd__buf_1
X_4263_ _8281_/Q _4194_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__mux2_1
X_6002_ _7969_/Q _6006_/B vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__and2_1
XFILLER_113_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4194_ _8444_/Q vssd1 vssd1 vccd1 vccd1 _4194_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2995_ clkbuf_0__2995_/X vssd1 vssd1 vccd1 vccd1 _6559_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7953_ _8490_/CLK _7953_/D vssd1 vssd1 vccd1 vccd1 _7953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7884_ _7884_/CLK _7884_/D vssd1 vssd1 vccd1 vccd1 _7884_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3616_ clkbuf_0__3616_/X vssd1 vssd1 vccd1 vccd1 _7384__144/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3978_/A vssd1 vssd1 vccd1 vccd1 _8403_/D sky130_fd_sc_hd__clkbuf_1
X_6766_ _8419_/Q _6789_/B _8420_/Q vssd1 vssd1 vccd1 vccd1 _7471_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5717_ _4144_/X _7876_/Q _5719_/S vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _5648_/A vssd1 vssd1 vccd1 vccd1 _7907_/D sky130_fd_sc_hd__clkbuf_1
X_8436_ _8441_/CLK _8436_/D vssd1 vssd1 vccd1 vccd1 _8436_/Q sky130_fd_sc_hd__dfxtp_1
X_5579_ _5579_/A vssd1 vssd1 vccd1 vccd1 _7937_/D sky130_fd_sc_hd__clkbuf_1
X_8367_ _8367_/CLK _8367_/D vssd1 vssd1 vccd1 vccd1 _8367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3377_ _6838_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3377_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8298_ _8315_/CLK _8298_/D vssd1 vssd1 vccd1 vccd1 _8298_/Q sky130_fd_sc_hd__dfxtp_1
X_7318_ _7247_/A _7316_/Y _7320_/D _7321_/B vssd1 vssd1 vccd1 vccd1 _7318_/X sky130_fd_sc_hd__a31o_1
XFILLER_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7249_ _7320_/B _7228_/C _7247_/X _7248_/X vssd1 vssd1 vccd1 vccd1 _8288_/D sky130_fd_sc_hd__o211a_1
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919__427 _6922__430/A vssd1 vssd1 vccd1 vccd1 _8105_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3059_ clkbuf_0__3059_/X vssd1 vssd1 vccd1 vccd1 _6263__199/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _8114_/Q _4244_/X _4952_/S vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__mux2_1
X_3901_ _3901_/A vssd1 vssd1 vccd1 vccd1 _8465_/D sky130_fd_sc_hd__clkbuf_1
X_4881_ _8289_/Q _4789_/A _8097_/Q _4814_/A _4715_/A vssd1 vssd1 vccd1 vccd1 _4881_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3401_ clkbuf_0__3401_/X vssd1 vssd1 vccd1 vccd1 _6918__426/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _3832_/A _5019_/B vssd1 vssd1 vccd1 vccd1 _3832_/Y sky130_fd_sc_hd__nor2_1
X_6620_ _7681_/A _7958_/Q _6622_/S vssd1 vssd1 vccd1 vccd1 _6621_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5502_ _5502_/A _5502_/B vssd1 vssd1 vccd1 vccd1 _5518_/S sky130_fd_sc_hd__nor2_2
X_6482_ _6482_/A vssd1 vssd1 vccd1 vccd1 _7722_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5433_ _5433_/A vssd1 vssd1 vccd1 vccd1 _8026_/D sky130_fd_sc_hd__clkbuf_1
X_8221_ _8221_/CLK _8221_/D vssd1 vssd1 vccd1 vccd1 _8221_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3231_ _6559_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3231_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_99_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5364_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__clkbuf_4
X_8152_ _8152_/CLK _8152_/D vssd1 vssd1 vccd1 vccd1 _8152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4315_ _4315_/A vssd1 vssd1 vccd1 vccd1 _8259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5295_ _5295_/A _5295_/B vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__or2_1
X_8083_ _8083_/CLK _8083_/D vssd1 vssd1 vccd1 vccd1 _8083_/Q sky130_fd_sc_hd__dfxtp_1
X_4246_ _4246_/A vssd1 vssd1 vccd1 vccd1 _8290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _8449_/Q vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__buf_2
XFILLER_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7936_ _7936_/CLK _7936_/D vssd1 vssd1 vccd1 vccd1 _7936_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7867_ _7867_/CLK _7867_/D vssd1 vssd1 vccd1 vccd1 _7867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6818_ _8433_/Q _8432_/Q _8431_/Q vssd1 vssd1 vccd1 vccd1 _6819_/A sky130_fd_sc_hd__and3_1
X_7798_ _7798_/CLK _7798_/D vssd1 vssd1 vccd1 vccd1 _7798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6749_ _6749_/A vssd1 vssd1 vccd1 vccd1 _6808_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8419_ _8425_/CLK _8419_/D vssd1 vssd1 vccd1 vccd1 _8419_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3429_ _7063_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3429_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6594__302 _6595__303/A vssd1 vssd1 vccd1 vccd1 _7942_/CLK sky130_fd_sc_hd__inv_2
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _5190_/S vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__clkbuf_2
X_4100_ _4100_/A vssd1 vssd1 vccd1 vccd1 _8357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4031_ _8387_/Q _3998_/X _4037_/S vssd1 vssd1 vccd1 vccd1 _4032_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5982_ _7961_/Q _5982_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__and2_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _4633_/X _4924_/X _4932_/Y _4900_/X vssd1 vssd1 vccd1 vccd1 _8123_/D sky130_fd_sc_hd__o211a_1
X_7721_ _7207_/A _7598_/C _7721_/S vssd1 vssd1 vccd1 vccd1 _7722_/B sky130_fd_sc_hd__mux2_1
X_7050__530 _7050__530/A vssd1 vssd1 vccd1 vccd1 _8211_/CLK sky130_fd_sc_hd__inv_2
X_4864_ _8106_/Q _4767_/A _4863_/X _4776_/A vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7652_ _7652_/A _7652_/B _7652_/C _7652_/D vssd1 vssd1 vccd1 vccd1 _7654_/C sky130_fd_sc_hd__or4_2
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _4801_/A vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__clkbuf_4
X_3815_ _3815_/A vssd1 vssd1 vccd1 vccd1 _5319_/A sky130_fd_sc_hd__clkbuf_2
X_7583_ _8436_/Q _7578_/X _7581_/X _7582_/X vssd1 vssd1 vccd1 vccd1 _8435_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6465_ _6465_/A vssd1 vssd1 vccd1 vccd1 _7849_/D sky130_fd_sc_hd__clkbuf_1
X_8204_ _8204_/CLK _8204_/D vssd1 vssd1 vccd1 vccd1 _8204_/Q sky130_fd_sc_hd__dfxtp_1
X_5416_ _3874_/X _8033_/Q _5422_/S vssd1 vssd1 vccd1 vccd1 _5417_/A sky130_fd_sc_hd__mux2_1
Xoutput120 _5948_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput142 _5905_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput131 _5955_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
X_6396_ _6412_/B vssd1 vssd1 vccd1 vccd1 _6408_/B sky130_fd_sc_hd__clkbuf_1
Xoutput153 _5927_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput175 _5863_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
Xoutput164 _5885_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5347_ _5347_/A vssd1 vssd1 vccd1 vccd1 _8059_/D sky130_fd_sc_hd__clkbuf_1
Xoutput186 _6087_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
X_8135_ _8135_/CLK _8135_/D vssd1 vssd1 vccd1 vccd1 _8135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5278_ _5278_/A _5278_/B _5278_/C vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__and3_1
Xoutput197 _6118_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
X_8066_ _8439_/CLK _8066_/D vssd1 vssd1 vccd1 vccd1 _8066_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _8066_/Q vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6582__294 _6583__295/A vssd1 vssd1 vccd1 vccd1 _7934_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7919_ _7919_/CLK _7919_/D vssd1 vssd1 vccd1 vccd1 _7919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8548__247 vssd1 vssd1 vccd1 vccd1 _8548__247/HI versionID[1] sky130_fd_sc_hd__conb_1
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _6115_/A sky130_fd_sc_hd__clkbuf_4
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _4419_/X _8154_/Q _4580_/S vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__mux2_1
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
Xinput55 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _3845_/B sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _3843_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _5960_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__clkbuf_2
Xinput88 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__buf_4
XFILLER_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput99 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _7615_/A sky130_fd_sc_hd__buf_4
X_5201_ _5305_/A _5199_/X _5200_/X vssd1 vssd1 vccd1 vccd1 _5202_/C sky130_fd_sc_hd__o21a_1
X_6181_ _6176_/X _7959_/Q _6178_/X _6180_/X _7748_/Q vssd1 vssd1 vccd1 vccd1 _7748_/D
+ sky130_fd_sc_hd__o32a_1
X_5132_ _5160_/A _5132_/B vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__and2_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5063_ _5190_/S vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4014_ _4359_/A vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _5965_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__and2_1
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5896_ _5896_/A vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7704_ _8016_/Q _7704_/B vssd1 vssd1 vccd1 vccd1 _7704_/Y sky130_fd_sc_hd__nand2_1
X_4916_ _4911_/X _4916_/B _6963_/C vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__and3b_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4847_ _7777_/Q _4765_/X _4845_/X _4846_/X vssd1 vssd1 vccd1 vccd1 _4847_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _4789_/A vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__clkbuf_2
X_7566_ _7563_/A _7562_/Y _7565_/X _7514_/X vssd1 vssd1 vccd1 vccd1 _8431_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7497_ _7497_/A _7497_/B _7497_/C _7497_/D vssd1 vssd1 vccd1 vccd1 _7500_/C sky130_fd_sc_hd__and4_1
Xclkbuf_1_1_0__3229_ clkbuf_0__3229_/X vssd1 vssd1 vccd1 vccd1 _6552__270/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6448_ _6448_/A vssd1 vssd1 vccd1 vccd1 _7841_/D sky130_fd_sc_hd__clkbuf_1
X_6379_ _7817_/Q _6343_/X _6371_/X _6376_/X _6378_/X vssd1 vssd1 vccd1 vccd1 _7817_/D
+ sky130_fd_sc_hd__a221o_1
X_8118_ _8118_/CLK _8118_/D vssd1 vssd1 vccd1 vccd1 _8118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6252__190 _6252__190/A vssd1 vssd1 vccd1 vccd1 _7782_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8049_ _8049_/CLK _8049_/D vssd1 vssd1 vccd1 vccd1 _8049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3059_ _6259_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3059_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3445_ clkbuf_0__3445_/X vssd1 vssd1 vccd1 vccd1 _7141__102/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3376_ clkbuf_0__3376_/X vssd1 vssd1 vccd1 vccd1 _6836__379/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8446_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5750_ _5750_/A vssd1 vssd1 vccd1 vccd1 _7862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5681_ _7892_/Q _4984_/X _5683_/S vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__mux2_1
X_4701_ _4673_/X _4696_/X _4700_/X _4746_/A vssd1 vssd1 vccd1 vccd1 _4701_/X sky130_fd_sc_hd__o211a_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4632_ _4670_/A vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__clkbuf_4
X_4563_ _4422_/X _8161_/Q _4567_/S vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__mux2_1
X_4494_ _5538_/B vssd1 vssd1 vccd1 vccd1 _4999_/C sky130_fd_sc_hd__buf_2
X_7282_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _8302_/D sky130_fd_sc_hd__nor2_1
X_6302_ _7832_/Q _6304_/C _6302_/C _6308_/B vssd1 vssd1 vccd1 vccd1 _6418_/B sky130_fd_sc_hd__or4_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6233_ _6233_/A vssd1 vssd1 vccd1 vccd1 _7774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6159_/X _7770_/Q _6161_/X _6163_/X _7738_/Q vssd1 vssd1 vccd1 vccd1 _7738_/D
+ sky130_fd_sc_hd__o32a_1
X_6906__418 _6906__418/A vssd1 vssd1 vccd1 vccd1 _8096_/CLK sky130_fd_sc_hd__inv_2
X_5115_ _5187_/A _5107_/X _5110_/X _5114_/X _5159_/A vssd1 vssd1 vccd1 vccd1 _5115_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5046_ _5054_/B _5046_/B vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__or2_2
Xclkbuf_1_0_0__3230_ clkbuf_0__3230_/X vssd1 vssd1 vccd1 vccd1 _6558__275/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5948_ _5948_/A vssd1 vssd1 vccd1 vccd1 _5948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6694__340 _6694__340/A vssd1 vssd1 vccd1 vccd1 _8004_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7549_ _8427_/Q _7510_/B _7544_/X _6754_/B vssd1 vssd1 vccd1 vccd1 _7550_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6846__387 _6846__387/A vssd1 vssd1 vccd1 vccd1 _8055_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6703__347 _6703__347/A vssd1 vssd1 vccd1 vccd1 _8011_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3428_ clkbuf_0__3428_/X vssd1 vssd1 vccd1 vccd1 _7059__537/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5802_ _5802_/A vssd1 vssd1 vccd1 vccd1 _7790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3994_ _4023_/S vssd1 vssd1 vccd1 vccd1 _4011_/S sky130_fd_sc_hd__buf_2
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6782_ _8418_/Q _6782_/B _6782_/C _7517_/A vssd1 vssd1 vccd1 vccd1 _7479_/B sky130_fd_sc_hd__nand4_2
X_5733_ _7869_/Q _5565_/A _5737_/S vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5664_ _5664_/A vssd1 vssd1 vccd1 vccd1 _7900_/D sky130_fd_sc_hd__clkbuf_1
X_8452_ _8452_/CLK _8452_/D vssd1 vssd1 vccd1 vccd1 _8452_/Q sky130_fd_sc_hd__dfxtp_1
X_5595_ _5574_/X _7930_/Q _5599_/S vssd1 vssd1 vccd1 vccd1 _5596_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4615_ _8124_/Q vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__inv_2
X_8383_ _8383_/CLK _8383_/D vssd1 vssd1 vccd1 vccd1 _8383_/Q sky130_fd_sc_hd__dfxtp_1
X_4546_ _4546_/A vssd1 vssd1 vccd1 vccd1 _8169_/D sky130_fd_sc_hd__clkbuf_1
X_7334_ _8081_/Q _7648_/B _7326_/X _7333_/X _7331_/X vssd1 vssd1 vccd1 vccd1 _8318_/D
+ sky130_fd_sc_hd__o311a_1
X_4477_ _4492_/S vssd1 vssd1 vccd1 vccd1 _4486_/S sky130_fd_sc_hd__buf_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7265_ _7208_/B _7270_/A _7264_/X vssd1 vssd1 vccd1 vccd1 _7265_/Y sky130_fd_sc_hd__o21bai_1
X_6216_ _6216_/A vssd1 vssd1 vccd1 vccd1 _7768_/D sky130_fd_sc_hd__clkbuf_1
X_7196_ _8301_/Q _7211_/C vssd1 vssd1 vccd1 vccd1 _7197_/B sky130_fd_sc_hd__xnor2_1
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6147_ _7773_/Q _7774_/Q vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__or2b_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_13 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_35 _6113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6078_ _7749_/Q _6082_/B vssd1 vssd1 vccd1 vccd1 _6078_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_46 _6119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_57 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_79 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _5029_/A vssd1 vssd1 vccd1 vccd1 _5084_/B sky130_fd_sc_hd__buf_2
XFILLER_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7382__142 _7384__144/A vssd1 vssd1 vccd1 vccd1 _8353_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _4362_/X _8224_/Q _4402_/S vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__mux2_1
X_5380_ _5349_/X _8050_/Q _5386_/S vssd1 vssd1 vccd1 vccd1 _5381_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4331_ _4331_/A vssd1 vssd1 vccd1 vccd1 _8252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4262_/A vssd1 vssd1 vccd1 vccd1 _8282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6001_ _6001_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6981__475 _6981__475/A vssd1 vssd1 vccd1 vccd1 _8156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4193_ _4193_/A vssd1 vssd1 vccd1 vccd1 _8336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2994_ clkbuf_0__2994_/X vssd1 vssd1 vccd1 vccd1 _6915_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7952_ _8490_/CLK _7952_/D vssd1 vssd1 vccd1 vccd1 _7952_/Q sky130_fd_sc_hd__dfxtp_1
X_6903_ _6909_/A vssd1 vssd1 vccd1 vccd1 _6903_/X sky130_fd_sc_hd__buf_1
X_7883_ _7883_/CLK _7883_/D vssd1 vssd1 vccd1 vccd1 _7883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3977_ _3925_/X _8403_/Q _3983_/S vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__mux2_1
X_6765_ _6786_/B _6789_/C vssd1 vssd1 vccd1 vccd1 _7471_/B sky130_fd_sc_hd__nand2_2
X_5716_ _5716_/A vssd1 vssd1 vccd1 vccd1 _7877_/D sky130_fd_sc_hd__clkbuf_1
X_8435_ _8441_/CLK _8435_/D vssd1 vssd1 vccd1 vccd1 _8435_/Q sky130_fd_sc_hd__dfxtp_1
X_5647_ _5571_/X _7907_/Q _5647_/S vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5578_ _5577_/X _7937_/Q _5581_/S vssd1 vssd1 vccd1 vccd1 _5579_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3445_ _7139_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3445_/X sky130_fd_sc_hd__clkbuf_16
X_8366_ _8366_/CLK _8366_/D vssd1 vssd1 vccd1 vccd1 _8366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3376_ _6832_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3376_/X sky130_fd_sc_hd__clkbuf_16
X_4529_ _4362_/X _8176_/Q _4531_/S vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__mux2_1
X_8297_ _8499_/CLK _8297_/D vssd1 vssd1 vccd1 vccd1 _8297_/Q sky130_fd_sc_hd__dfxtp_1
X_7317_ _8314_/Q _7317_/B vssd1 vssd1 vccd1 vccd1 _7320_/D sky130_fd_sc_hd__nand2_1
XFILLER_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7248_ _7345_/S vssd1 vssd1 vccd1 vccd1 _7248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7179_ _7217_/A _7217_/B _7193_/D vssd1 vssd1 vccd1 vccd1 _7181_/A sky130_fd_sc_hd__nand3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6546__265 _6546__265/A vssd1 vssd1 vccd1 vccd1 _7905_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3058_ clkbuf_0__3058_/X vssd1 vssd1 vccd1 vccd1 _6258__195/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7134__97 _7134__97/A vssd1 vssd1 vccd1 vccd1 _8278_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
X_7452__24 _7453__25/A vssd1 vssd1 vccd1 vccd1 _8410_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3900_ _8465_/Q _3812_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__mux2_1
X_4880_ _4753_/A _8052_/Q _7936_/Q _4796_/A vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__a22o_1
X_7389__148 _7389__148/A vssd1 vssd1 vccd1 vccd1 _8359_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3400_ clkbuf_0__3400_/X vssd1 vssd1 vccd1 vccd1 _6917_/A sky130_fd_sc_hd__clkbuf_4
X_3831_ _8071_/Q _8076_/Q vssd1 vssd1 vccd1 vccd1 _5019_/B sky130_fd_sc_hd__and2b_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5501_ _5501_/A vssd1 vssd1 vccd1 vccd1 _7992_/D sky130_fd_sc_hd__clkbuf_1
X_6481_ _6481_/A vssd1 vssd1 vccd1 vccd1 _7854_/D sky130_fd_sc_hd__clkbuf_1
X_5432_ _8026_/Q _4431_/X _5440_/S vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__mux2_1
X_8220_ _8220_/CLK _8220_/D vssd1 vssd1 vccd1 vccd1 _8220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3230_ _6553_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3230_/X sky130_fd_sc_hd__clkbuf_16
X_5363_ _5363_/A vssd1 vssd1 vccd1 vccd1 _8055_/D sky130_fd_sc_hd__clkbuf_1
X_8151_ _8151_/CLK _8151_/D vssd1 vssd1 vccd1 vccd1 _8151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _8259_/Q _4188_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__mux2_1
X_6489__219 _6490__220/A vssd1 vssd1 vccd1 vccd1 _7859_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5294_ _8279_/Q _8000_/Q _5294_/S vssd1 vssd1 vccd1 vccd1 _5295_/B sky130_fd_sc_hd__mux2_1
X_8082_ _8082_/CLK _8082_/D vssd1 vssd1 vccd1 vccd1 _8082_/Q sky130_fd_sc_hd__dfxtp_1
X_4245_ _8290_/Q _4244_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _4176_/A vssd1 vssd1 vccd1 vccd1 _8341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7935_ _7935_/CLK _7935_/D vssd1 vssd1 vccd1 vccd1 _7935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7866_ _7866_/CLK _7866_/D vssd1 vssd1 vccd1 vccd1 _7866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6817_ _7586_/A vssd1 vssd1 vccd1 vccd1 _7584_/B sky130_fd_sc_hd__clkbuf_2
X_7797_ _7797_/CLK _7797_/D vssd1 vssd1 vccd1 vccd1 _7797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6748_ _6751_/A vssd1 vssd1 vccd1 vccd1 _6808_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8418_ _8418_/CLK _8418_/D vssd1 vssd1 vccd1 vccd1 _8418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8349_ _8349_/CLK _8349_/D vssd1 vssd1 vccd1 vccd1 _8349_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3428_ _7057_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3428_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6925__432 _6926__433/A vssd1 vssd1 vccd1 vccd1 _8110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7395__152 _7396__153/A vssd1 vssd1 vccd1 vccd1 _8363_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4030_ _4030_/A vssd1 vssd1 vccd1 vccd1 _8388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _5981_/A vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7720_ _7720_/A vssd1 vssd1 vccd1 vccd1 _8498_/D sky130_fd_sc_hd__clkbuf_1
X_4932_ _4932_/A _4932_/B vssd1 vssd1 vccd1 vccd1 _4932_/Y sky130_fd_sc_hd__nand2_1
X_7651_ _7651_/A vssd1 vssd1 vccd1 vccd1 _8478_/D sky130_fd_sc_hd__clkbuf_1
X_4863_ _4770_/A _8037_/Q _7865_/Q _4769_/A vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4794_ _4794_/A vssd1 vssd1 vccd1 vccd1 _4932_/B sky130_fd_sc_hd__buf_2
X_7582_ _7582_/A vssd1 vssd1 vccd1 vccd1 _7582_/X sky130_fd_sc_hd__clkbuf_2
X_3814_ _8076_/Q vssd1 vssd1 vccd1 vccd1 _3815_/A sky130_fd_sc_hd__inv_2
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6464_ _7849_/Q _7964_/Q _6466_/S vssd1 vssd1 vccd1 vccd1 _6465_/A sky130_fd_sc_hd__mux2_1
Xoutput110 _5968_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
X_8203_ _8203_/CLK _8203_/D vssd1 vssd1 vccd1 vccd1 _8203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5415_ _5415_/A vssd1 vssd1 vccd1 vccd1 _8034_/D sky130_fd_sc_hd__clkbuf_1
Xoutput121 _5990_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput143 _5907_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput132 _5957_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
X_6395_ _6395_/A vssd1 vssd1 vccd1 vccd1 _7680_/A sky130_fd_sc_hd__clkbuf_4
Xoutput154 _5929_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput165 _5888_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
X_5346_ _5343_/X _8059_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__mux2_1
Xoutput176 _6127_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8134_ _8134_/CLK _8134_/D vssd1 vssd1 vccd1 vccd1 _8134_/Q sky130_fd_sc_hd__dfxtp_1
X_5277_ _5220_/A _5275_/X _5276_/X vssd1 vssd1 vccd1 vccd1 _5278_/C sky130_fd_sc_hd__o21ai_1
Xoutput187 _6090_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput198 _6120_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
X_8065_ _8439_/CLK _8065_/D vssd1 vssd1 vccd1 vccd1 _8065_/Q sky130_fd_sc_hd__dfxtp_2
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _8296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _5430_/B _4178_/B vssd1 vssd1 vccd1 vccd1 _4175_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_1_0_0__3392_ clkbuf_0__3392_/X vssd1 vssd1 vccd1 vccd1 _6891__410/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7918_ _7918_/CLK _7918_/D vssd1 vssd1 vccd1 vccd1 _7918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6994__485 _6994__485/A vssd1 vssd1 vccd1 vccd1 _8166_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7849_ _8060_/CLK _7849_/D vssd1 vssd1 vccd1 vccd1 _7849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7027__511 _7029__513/A vssd1 vssd1 vccd1 vccd1 _8192_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8531__230 vssd1 vssd1 vccd1 vccd1 _8531__230/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _6117_/A sky130_fd_sc_hd__clkbuf_4
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_4
Xinput45 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _3843_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_116_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput56 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _3845_/A sky130_fd_sc_hd__clkbuf_1
Xinput89 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__buf_4
Xinput67 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _5963_/A sky130_fd_sc_hd__buf_4
Xinput78 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5213_/A _8030_/Q _7795_/Q _5215_/A _5073_/A vssd1 vssd1 vccd1 vccd1 _5200_/X
+ sky130_fd_sc_hd__o221a_1
X_6180_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6180_/X sky130_fd_sc_hd__clkbuf_2
X_5131_ _8471_/Q _8212_/Q _8204_/Q _8236_/Q _5060_/A _5044_/A vssd1 vssd1 vccd1 vccd1
+ _5132_/B sky130_fd_sc_hd__mux4_1
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5062_ _5062_/A vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ _8444_/Q vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__buf_2
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5964_ _5964_/A vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6503__230 _6503__230/A vssd1 vssd1 vccd1 vccd1 _7870_/CLK sky130_fd_sc_hd__inv_2
X_7703_ _7703_/A vssd1 vssd1 vccd1 vccd1 _7707_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5895_ _7696_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5896_/A sky130_fd_sc_hd__or2_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4915_ _6854_/A vssd1 vssd1 vccd1 vccd1 _6963_/C sky130_fd_sc_hd__buf_2
X_4846_ _4796_/A _7905_/Q _7897_/Q _4753_/A _4757_/A vssd1 vssd1 vccd1 vccd1 _4846_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7565_ _7563_/Y _7504_/A _6820_/C _7564_/Y _7556_/X vssd1 vssd1 vccd1 vccd1 _7565_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4777_ _4753_/X _8055_/Q _7939_/Q _4749_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4777_/X
+ sky130_fd_sc_hd__a221o_1
X_6516_ _6522_/A vssd1 vssd1 vccd1 vccd1 _6516_/X sky130_fd_sc_hd__buf_1
X_7496_ _6791_/Y _6792_/X _6781_/X _6785_/X _6787_/X vssd1 vssd1 vccd1 vccd1 _7497_/D
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_1_1_0__3228_ clkbuf_0__3228_/X vssd1 vssd1 vccd1 vccd1 _6544__263/A sky130_fd_sc_hd__clkbuf_4
X_6447_ _7841_/Q _5971_/A _6455_/S vssd1 vssd1 vccd1 vccd1 _6448_/A sky130_fd_sc_hd__mux2_1
X_6378_ _6391_/A vssd1 vssd1 vccd1 vccd1 _6378_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _5329_/A _7604_/A _5329_/C vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__and3_1
X_8117_ _8117_/CLK _8117_/D vssd1 vssd1 vccd1 vccd1 _8117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8048_ _8048_/CLK _8048_/D vssd1 vssd1 vccd1 vccd1 _8048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3058_ _6253_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3058_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3375_ clkbuf_0__3375_/X vssd1 vssd1 vccd1 vccd1 _6873_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8515__214 vssd1 vssd1 vccd1 vccd1 _8515__214/HI core0Index[1] sky130_fd_sc_hd__conb_1
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7643__49 _7643__49/A vssd1 vssd1 vccd1 vccd1 _8472_/CLK sky130_fd_sc_hd__inv_2
X_7100__70 _7100__70/A vssd1 vssd1 vccd1 vccd1 _8251_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5680_ _5680_/A vssd1 vssd1 vccd1 vccd1 _7893_/D sky130_fd_sc_hd__clkbuf_1
X_4700_ _4663_/X _4697_/X _4699_/X vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__a21o_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4631_ _8123_/Q vssd1 vssd1 vccd1 vccd1 _4670_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _4562_/A vssd1 vssd1 vccd1 vccd1 _8162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4493_ _4493_/A vssd1 vssd1 vccd1 vccd1 _8191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7281_ _7211_/A _7280_/X _7272_/X _7241_/Y vssd1 vssd1 vccd1 vccd1 _7282_/B sky130_fd_sc_hd__o2bb2a_1
X_6301_ _7834_/Q _6301_/B _7833_/Q vssd1 vssd1 vccd1 vccd1 _6308_/B sky130_fd_sc_hd__or3b_1
X_6232_ _6231_/X _6232_/B vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6172_/A vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__clkbuf_2
X_5114_ _5038_/A _5112_/X _5113_/X vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6072_/A _6091_/X _6092_/X _6093_/X vssd1 vssd1 vccd1 vccd1 _6094_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5045_ _7799_/Q _8007_/Q _8286_/Q _8034_/Q _5269_/S _5044_/X vssd1 vssd1 vccd1 vccd1
+ _5045_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _5947_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__and2_1
XFILLER_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _7600_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__or2_1
X_4829_ _8153_/Q _4795_/X _4796_/X _8115_/Q vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__a22o_1
X_7548_ _7554_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _8426_/D sky130_fd_sc_hd__nor2_1
X_7479_ _8495_/Q _7479_/B _7479_/C vssd1 vssd1 vccd1 vccd1 _7479_/X sky130_fd_sc_hd__and3_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7086__58 _7088__60/A vssd1 vssd1 vccd1 vccd1 _8239_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3427_ clkbuf_0__3427_/X vssd1 vssd1 vccd1 vccd1 _7056__535/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3631_ clkbuf_0__3631_/X vssd1 vssd1 vccd1 vccd1 _7620__30/A sky130_fd_sc_hd__clkbuf_4
X_6850_ _6873_/A vssd1 vssd1 vccd1 vccd1 _6850_/X sky130_fd_sc_hd__buf_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5801_ _3874_/X _7790_/Q _5807_/S vssd1 vssd1 vccd1 vccd1 _5802_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6781_ _6774_/X _6775_/Y _6777_/Y _6779_/Y _6780_/X vssd1 vssd1 vccd1 vccd1 _6781_/X
+ sky130_fd_sc_hd__o2111a_1
X_5732_ _5732_/A vssd1 vssd1 vccd1 vccd1 _7870_/D sky130_fd_sc_hd__clkbuf_1
X_3993_ _4083_/A _5797_/B vssd1 vssd1 vccd1 vccd1 _4023_/S sky130_fd_sc_hd__nor2_2
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6719__355 _6719__355/A vssd1 vssd1 vccd1 vccd1 _8022_/CLK sky130_fd_sc_hd__inv_2
X_5663_ _5568_/X _7900_/Q _5665_/S vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__mux2_1
X_6912__423 _6914__425/A vssd1 vssd1 vccd1 vccd1 _8101_/CLK sky130_fd_sc_hd__inv_2
X_8451_ _8451_/CLK _8451_/D vssd1 vssd1 vccd1 vccd1 _8451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5594_ _5594_/A vssd1 vssd1 vccd1 vccd1 _7931_/D sky130_fd_sc_hd__clkbuf_1
X_8382_ _8382_/CLK _8382_/D vssd1 vssd1 vccd1 vccd1 _8382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4614_ _4745_/A vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4545_ _8169_/Q _4448_/X _4549_/S vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__mux2_1
X_7333_ _8318_/Q _7337_/B vssd1 vssd1 vccd1 vccd1 _7333_/X sky130_fd_sc_hd__or2_1
Xclkbuf_0__3392_ _6886_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3392_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4476_ _5815_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _4492_/S sky130_fd_sc_hd__nor2_2
X_7264_ _7295_/A vssd1 vssd1 vccd1 vccd1 _7264_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6215_ _7607_/A _7768_/Q _6217_/S vssd1 vssd1 vccd1 vccd1 _6216_/A sky130_fd_sc_hd__mux2_1
X_7195_ _7195_/A _7195_/B vssd1 vssd1 vccd1 vccd1 _7195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6146_ _6328_/A vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__buf_4
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_14 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_25 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_47 _6119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_36 _6113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_58 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6077_ _7824_/Q input10/X _6077_/S vssd1 vssd1 vccd1 vccd1 _6077_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_69 _5945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5054_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__and2_1
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _8252_/Q _4185_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ _8282_/Q _4191_/X _4261_/S vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6000_ _6000_/A _6105_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__and2_2
X_4192_ _8336_/Q _4191_/X _4192_/S vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7255__110 _7255__110/A vssd1 vssd1 vccd1 vccd1 _8293_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7951_ _7951_/CLK _7951_/D vssd1 vssd1 vccd1 vccd1 _7951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7882_ _7882_/CLK _7882_/D vssd1 vssd1 vccd1 vccd1 _7882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3614_ clkbuf_0__3614_/X vssd1 vssd1 vccd1 vccd1 _7373__135/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3976_ _3976_/A vssd1 vssd1 vccd1 vccd1 _8404_/D sky130_fd_sc_hd__clkbuf_1
X_6764_ _6359_/X _6763_/Y _7492_/B _7698_/A vssd1 vssd1 vccd1 vccd1 _6794_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6695_ _6701_/A vssd1 vssd1 vccd1 vccd1 _6695_/X sky130_fd_sc_hd__buf_1
X_5715_ _4141_/X _7877_/Q _5719_/S vssd1 vssd1 vccd1 vccd1 _5716_/A sky130_fd_sc_hd__mux2_1
X_5646_ _5646_/A vssd1 vssd1 vccd1 vccd1 _7908_/D sky130_fd_sc_hd__clkbuf_1
X_8434_ _8441_/CLK _8434_/D vssd1 vssd1 vccd1 vccd1 _8434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5577_ _5577_/A vssd1 vssd1 vccd1 vccd1 _5577_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3444_ _7138_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3444_/X sky130_fd_sc_hd__clkbuf_16
X_8365_ _8365_/CLK _8365_/D vssd1 vssd1 vccd1 vccd1 _8365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8296_ _8296_/CLK _8296_/D vssd1 vssd1 vccd1 vccd1 _8296_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3375_ _6831_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3375_/X sky130_fd_sc_hd__clkbuf_16
X_4528_ _4528_/A vssd1 vssd1 vccd1 vccd1 _8177_/D sky130_fd_sc_hd__clkbuf_1
X_7316_ _7320_/C vssd1 vssd1 vccd1 vccd1 _7316_/Y sky130_fd_sc_hd__inv_2
X_4459_ _4342_/X _8206_/Q _4467_/S vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__mux2_1
X_7247_ _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7247_/X sky130_fd_sc_hd__or2_1
XFILLER_104_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7178_ _8489_/Q _7178_/B vssd1 vssd1 vccd1 vccd1 _7183_/B sky130_fd_sc_hd__xor2_1
X_7021__506 _7024__509/A vssd1 vssd1 vccd1 vccd1 _8187_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6129_ _6480_/A _6473_/A _6129_/C vssd1 vssd1 vccd1 vccd1 _6130_/A sky130_fd_sc_hd__and3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3057_ clkbuf_0__3057_/X vssd1 vssd1 vccd1 vccd1 _6249__187/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7437__11 _7439__13/A vssd1 vssd1 vccd1 vccd1 _8397_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _8076_/Q _5054_/A vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__and2b_1
XFILLER_60_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5500_ _5373_/X _7992_/Q _5500_/S vssd1 vssd1 vccd1 vccd1 _5501_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ _6480_/A _6480_/B _6480_/C vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__and3_1
X_5431_ _5446_/S vssd1 vssd1 vccd1 vccd1 _5440_/S sky130_fd_sc_hd__clkbuf_4
X_8150_ _8150_/CLK _8150_/D vssd1 vssd1 vccd1 vccd1 _8150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5362_ _5361_/X _8055_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__mux2_1
X_4313_ _4313_/A vssd1 vssd1 vccd1 vccd1 _8260_/D sky130_fd_sc_hd__clkbuf_1
X_7101_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7101_/X sky130_fd_sc_hd__buf_1
X_8081_ _8081_/CLK _8081_/D vssd1 vssd1 vccd1 vccd1 _8081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7032_ _7038_/A vssd1 vssd1 vccd1 vccd1 _7032_/X sky130_fd_sc_hd__buf_1
X_5293_ _8450_/Q _5227_/X _5220_/A _5291_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5293_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4244_ _8061_/Q vssd1 vssd1 vccd1 vccd1 _4244_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4175_ _8341_/Q _4022_/X _4175_/S vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7934_ _7934_/CLK _7934_/D vssd1 vssd1 vccd1 vccd1 _7934_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7865_ _7865_/CLK _7865_/D vssd1 vssd1 vccd1 vccd1 _7865_/Q sky130_fd_sc_hd__dfxtp_1
X_7796_ _7796_/CLK _7796_/D vssd1 vssd1 vccd1 vccd1 _7796_/Q sky130_fd_sc_hd__dfxtp_1
X_6816_ _7500_/A _6816_/B _6816_/C _7572_/C vssd1 vssd1 vccd1 vccd1 _7586_/A sky130_fd_sc_hd__and4_1
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6747_ _8487_/Q vssd1 vssd1 vccd1 vccd1 _7459_/A sky130_fd_sc_hd__clkinv_4
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3959_ _3959_/A vssd1 vssd1 vccd1 vccd1 _8410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5629_ _7915_/Q _4987_/X _5629_/S vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__mux2_1
X_8417_ _8418_/CLK _8417_/D vssd1 vssd1 vccd1 vccd1 _8417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3427_ _7051_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3427_/X sky130_fd_sc_hd__clkbuf_16
X_8348_ _8348_/CLK _8348_/D vssd1 vssd1 vccd1 vccd1 _8348_/Q sky130_fd_sc_hd__dfxtp_1
X_6552__270 _6552__270/A vssd1 vssd1 vccd1 vccd1 _7910_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8279_ _8279_/CLK _8279_/D vssd1 vssd1 vccd1 vccd1 _8279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _7960_/Q _5982_/B vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__and2_1
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4760_/X _4924_/X _4930_/Y _4900_/X vssd1 vssd1 vccd1 vccd1 _8124_/D sky130_fd_sc_hd__o211a_1
X_4862_ _4789_/X _7857_/Q _4803_/X _8090_/Q _4663_/A vssd1 vssd1 vccd1 vccd1 _4862_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7650_ _8078_/Q _7662_/A vssd1 vssd1 vccd1 vccd1 _7651_/A sky130_fd_sc_hd__and2_1
X_3813_ _8077_/Q vssd1 vssd1 vccd1 vccd1 _4287_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4793_ _4793_/A vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__buf_2
X_6495__224 _6496__225/A vssd1 vssd1 vccd1 vccd1 _7864_/CLK sky130_fd_sc_hd__inv_2
X_7581_ _8435_/Q _7584_/B vssd1 vssd1 vccd1 vccd1 _7581_/X sky130_fd_sc_hd__or2_1
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6872__395 _6872__395/A vssd1 vssd1 vccd1 vccd1 _8071_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6463_ _6463_/A vssd1 vssd1 vccd1 vccd1 _7848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8202_ _8202_/CLK _8202_/D vssd1 vssd1 vccd1 vccd1 _8202_/Q sky130_fd_sc_hd__dfxtp_1
X_5414_ _3812_/X _8034_/Q _5422_/S vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__mux2_1
Xoutput122 _5992_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput111 _5970_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
Xoutput133 _5959_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
XFILLER_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6394_ _8485_/Q vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__clkbuf_4
X_8133_ _8133_/CLK _8133_/D vssd1 vssd1 vccd1 vccd1 _8133_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput144 _5910_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput155 _5932_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput166 _5890_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
X_5345_ _5374_/S vssd1 vssd1 vccd1 vccd1 _5362_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput177 _6019_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
X_5276_ _5213_/A _8028_/Q _7793_/Q _5292_/B _5098_/A vssd1 vssd1 vccd1 vccd1 _5276_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput199 _6026_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput188 _6022_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
X_8064_ _8439_/CLK _8064_/D vssd1 vssd1 vccd1 vccd1 _8064_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4227_ _8296_/Q _4223_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _4158_/A vssd1 vssd1 vccd1 vccd1 _8349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3391_ clkbuf_0__3391_/X vssd1 vssd1 vccd1 vccd1 _6885__405/A sky130_fd_sc_hd__clkbuf_4
X_4089_ _8362_/Q _4002_/X _4093_/S vssd1 vssd1 vccd1 vccd1 _4090_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7917_ _7917_/CLK _7917_/D vssd1 vssd1 vccd1 vccd1 _7917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7848_ _8141_/CLK _7848_/D vssd1 vssd1 vccd1 vccd1 _7848_/Q sky130_fd_sc_hd__dfxtp_1
X_7779_ _7779_/CLK _7779_/D vssd1 vssd1 vccd1 vccd1 _7779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6665__316 _6667__318/A vssd1 vssd1 vccd1 vccd1 _7980_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6264__200 _6264__200/A vssd1 vssd1 vccd1 vccd1 _7792_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _6119_/A sky130_fd_sc_hd__clkbuf_4
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _3842_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput68 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__buf_4
Xinput79 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__clkbuf_2
Xinput57 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
X_5130_ _5128_/X _5129_/X _5186_/S vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ _8364_/Q _8348_/Q _8340_/Q _8372_/Q _5060_/X _5052_/X vssd1 vssd1 vccd1 vccd1
+ _5061_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4012_ _4012_/A vssd1 vssd1 vccd1 vccd1 _8392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5963_ _5963_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__and2_1
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7702_ _7721_/S vssd1 vssd1 vccd1 vccd1 _7707_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4914_ _4903_/A _4911_/B _7645_/B _4999_/B vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__a31o_1
X_5894_ _5894_/A vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _7945_/Q _4653_/B _4767_/X vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__a21o_1
X_7633_ _7633_/A vssd1 vssd1 vccd1 vccd1 _7633_/X sky130_fd_sc_hd__buf_1
X_4776_ _4776_/A vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__clkbuf_2
X_7564_ _7577_/A _7577_/B vssd1 vssd1 vccd1 vccd1 _7564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3227_ clkbuf_0__3227_/X vssd1 vssd1 vccd1 vccd1 _6540__260/A sky130_fd_sc_hd__clkbuf_4
X_7495_ _8492_/Q _6763_/Y _6767_/Y _6768_/X vssd1 vssd1 vccd1 vccd1 _7497_/C sky130_fd_sc_hd__o2bb2a_1
X_6446_ _6468_/A vssd1 vssd1 vccd1 vccd1 _6455_/S sky130_fd_sc_hd__buf_2
X_6377_ _7654_/B _6353_/X _6355_/X _6482_/A vssd1 vssd1 vccd1 vccd1 _6391_/A sky130_fd_sc_hd__a31o_2
XFILLER_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8116_ _8116_/CLK _8116_/D vssd1 vssd1 vccd1 vccd1 _8116_/Q sky130_fd_sc_hd__dfxtp_1
X_5328_ _5328_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _5329_/C sky130_fd_sc_hd__or2_1
XFILLER_114_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8047_ _8047_/CLK _8047_/D vssd1 vssd1 vccd1 vccd1 _8047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5259_ _8224_/Q _5227_/X _5179_/X _8374_/Q _5062_/A vssd1 vssd1 vccd1 vccd1 _5259_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__3057_ _6247_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3057_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3443_ clkbuf_0__3443_/X vssd1 vssd1 vccd1 vccd1 _7136__99/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3374_ clkbuf_0__3374_/X vssd1 vssd1 vccd1 vccd1 _6827__372/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7628__36 _7629__37/A vssd1 vssd1 vccd1 vccd1 _8459_/CLK sky130_fd_sc_hd__inv_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6565__280 _6565__280/A vssd1 vssd1 vccd1 vccd1 _7920_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ _4630_/A vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ _7207_/A _6293_/X _6299_/X vssd1 vssd1 vccd1 vccd1 _6300_/X sky130_fd_sc_hd__a21o_1
X_4561_ _4419_/X _8162_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__mux2_1
X_4492_ _8191_/Q _4247_/X _4492_/S vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7280_ _7295_/A vssd1 vssd1 vccd1 vccd1 _7280_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6231_ _6231_/A _6231_/B _6231_/C vssd1 vssd1 vccd1 vccd1 _6231_/X sky130_fd_sc_hd__and3_1
XFILLER_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6159_/X _7769_/Q _6161_/X _6153_/X _7737_/Q vssd1 vssd1 vccd1 vccd1 _7737_/D
+ sky130_fd_sc_hd__o32a_1
X_5113_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__buf_2
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6093_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5044_ _5044_/A vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__buf_4
XFILLER_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8538__237 vssd1 vssd1 vccd1 vccd1 _8538__237/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
X_6995_ _7007_/A vssd1 vssd1 vccd1 vccd1 _6995_/X sky130_fd_sc_hd__buf_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5946_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5877_ _5877_/A vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__clkbuf_1
X_4828_ _4757_/X _4826_/X _4827_/X vssd1 vssd1 vccd1 vccd1 _4828_/X sky130_fd_sc_hd__o21a_1
X_7616_ _7616_/A vssd1 vssd1 vccd1 vccd1 _8449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _8124_/Q vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7547_ _8426_/Q _7530_/X _7544_/X _7494_/B vssd1 vssd1 vccd1 vccd1 _7548_/B sky130_fd_sc_hd__o2bb2a_1
X_7478_ _7478_/A _7478_/B vssd1 vssd1 vccd1 vccd1 _7478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6429_ _7833_/Q _5954_/A _6433_/S vssd1 vssd1 vccd1 vccd1 _6430_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8441_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3426_ clkbuf_0__3426_/X vssd1 vssd1 vccd1 vccd1 _7048__528/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7070__546 _7073__549/A vssd1 vssd1 vccd1 vccd1 _8227_/CLK sky130_fd_sc_hd__inv_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3630_ clkbuf_0__3630_/X vssd1 vssd1 vccd1 vccd1 _7639_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3992_ _4342_/A vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__buf_2
X_6678__326 _6682__330/A vssd1 vssd1 vccd1 vccd1 _7990_/CLK sky130_fd_sc_hd__inv_2
X_5800_ _5800_/A vssd1 vssd1 vccd1 vccd1 _7791_/D sky130_fd_sc_hd__clkbuf_1
X_6780_ _7207_/A _7517_/A vssd1 vssd1 vccd1 vccd1 _6780_/X sky130_fd_sc_hd__or2_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _7870_/Q _5562_/A _5737_/S vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__mux2_1
X_5662_ _5662_/A vssd1 vssd1 vccd1 vccd1 _7901_/D sky130_fd_sc_hd__clkbuf_1
X_8450_ _8450_/CLK _8450_/D vssd1 vssd1 vccd1 vccd1 _8450_/Q sky130_fd_sc_hd__dfxtp_1
X_5593_ _5571_/X _7931_/Q _5593_/S vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__mux2_1
X_6277__210 _6277__210/A vssd1 vssd1 vccd1 vccd1 _7802_/CLK sky130_fd_sc_hd__inv_2
X_8381_ _8381_/CLK _8381_/D vssd1 vssd1 vccd1 vccd1 _8381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4613_ _4613_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__nor2_1
X_4544_ _4544_/A vssd1 vssd1 vccd1 vccd1 _8170_/D sky130_fd_sc_hd__clkbuf_1
X_7332_ _8080_/Q _7648_/B _7326_/X _7330_/X _7331_/X vssd1 vssd1 vccd1 vccd1 _8317_/D
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_0__3391_ _6880_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3391_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7263_ _7247_/A _7247_/B _7262_/B vssd1 vssd1 vccd1 vccd1 _7295_/A sky130_fd_sc_hd__a21o_2
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _5538_/A _4475_/B _5538_/B vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__or3_2
X_6214_ _6214_/A vssd1 vssd1 vccd1 vccd1 _7767_/D sky130_fd_sc_hd__clkbuf_1
X_7194_ _7211_/C _7193_/C _7193_/D _8309_/Q vssd1 vssd1 vccd1 vccd1 _7195_/B sky130_fd_sc_hd__a31o_1
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6145_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6328_/A sky130_fd_sc_hd__buf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6076_ _6072_/X _6073_/X _6074_/X _6075_/X vssd1 vssd1 vccd1 vccd1 _6076_/X sky130_fd_sc_hd__o211a_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_48 _6119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_26 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5027_ _8070_/Q _8069_/Q _8068_/Q vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__and3_1
XINSDIODE2_37 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_59 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7091__62 _7094__65/A vssd1 vssd1 vccd1 vccd1 _8243_/CLK sky130_fd_sc_hd__inv_2
X_7416__170 _7416__170/A vssd1 vssd1 vccd1 vccd1 _8381_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5929_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3409_ clkbuf_0__3409_/X vssd1 vssd1 vccd1 vccd1 _6968__464/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _4260_/A vssd1 vssd1 vccd1 vccd1 _8283_/D sky130_fd_sc_hd__clkbuf_1
X_4191_ _8445_/Q vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__clkbuf_4
X_7359__124 _7360__125/A vssd1 vssd1 vccd1 vccd1 _8335_/CLK sky130_fd_sc_hd__inv_2
X_7950_ _7950_/CLK _7950_/D vssd1 vssd1 vccd1 vccd1 _7950_/Q sky130_fd_sc_hd__dfxtp_1
X_6725__360 _6725__360/A vssd1 vssd1 vccd1 vccd1 _8027_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7881_ _7881_/CLK _7881_/D vssd1 vssd1 vccd1 vccd1 _7881_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3613_ clkbuf_0__3613_/X vssd1 vssd1 vccd1 vccd1 _7366__129/A sky130_fd_sc_hd__clkbuf_4
X_6832_ _6844_/A vssd1 vssd1 vccd1 vccd1 _6832_/X sky130_fd_sc_hd__buf_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3975_ _3916_/X _8404_/Q _3983_/S vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__mux2_1
X_6763_ _7465_/B _7465_/C vssd1 vssd1 vccd1 vccd1 _6763_/Y sky130_fd_sc_hd__nand2_2
X_5714_ _5714_/A vssd1 vssd1 vccd1 vccd1 _7878_/D sky130_fd_sc_hd__clkbuf_1
X_5645_ _5568_/X _7908_/Q _5647_/S vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8433_ _8433_/CLK _8433_/D vssd1 vssd1 vccd1 vccd1 _8433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3443_ _7132_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3443_/X sky130_fd_sc_hd__clkbuf_16
X_5576_ _5576_/A vssd1 vssd1 vccd1 vccd1 _7938_/D sky130_fd_sc_hd__clkbuf_1
X_7425__1 _7426__2/A vssd1 vssd1 vccd1 vccd1 _8387_/CLK sky130_fd_sc_hd__inv_2
X_8364_ _8364_/CLK _8364_/D vssd1 vssd1 vccd1 vccd1 _8364_/Q sky130_fd_sc_hd__dfxtp_1
X_8295_ _8295_/CLK _8295_/D vssd1 vssd1 vccd1 vccd1 _8295_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3374_ _6825_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3374_/X sky130_fd_sc_hd__clkbuf_16
X_4527_ _4359_/X _8177_/Q _4531_/S vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__mux2_1
X_7315_ _7315_/A _7321_/B vssd1 vssd1 vccd1 vccd1 _7315_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4458_ _4473_/S vssd1 vssd1 vccd1 vccd1 _4467_/S sky130_fd_sc_hd__buf_2
X_7246_ _8287_/Q _7246_/B _7246_/C _7246_/D vssd1 vssd1 vccd1 vccd1 _7247_/B sky130_fd_sc_hd__and4_1
X_7177_ _8307_/Q _7216_/B vssd1 vssd1 vccd1 vccd1 _7178_/B sky130_fd_sc_hd__xnor2_2
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _8230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6128_ _6206_/A vssd1 vssd1 vccd1 vccd1 _6480_/A sky130_fd_sc_hd__clkinv_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6059_ _7744_/Q _6063_/B vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__or2_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7119__85 _7119__85/A vssd1 vssd1 vccd1 vccd1 _8266_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5430_ _5502_/A _5430_/B vssd1 vssd1 vccd1 vccd1 _5446_/S sky130_fd_sc_hd__nor2_2
X_5361_ _5571_/A vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4312_ _8260_/Q _4185_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5292_ _8458_/Q _5292_/B vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__or2_1
X_8080_ _8080_/CLK _8080_/D vssd1 vssd1 vccd1 vccd1 _8080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4243_ _4243_/A vssd1 vssd1 vccd1 vccd1 _8291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4174_/A vssd1 vssd1 vccd1 vccd1 _8342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7933_ _7933_/CLK _7933_/D vssd1 vssd1 vccd1 vccd1 _7933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7864_ _7864_/CLK _7864_/D vssd1 vssd1 vccd1 vccd1 _7864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7795_ _7795_/CLK _7795_/D vssd1 vssd1 vccd1 vccd1 _7795_/Q sky130_fd_sc_hd__dfxtp_1
X_6815_ _8413_/Q _7508_/A vssd1 vssd1 vccd1 vccd1 _7572_/C sky130_fd_sc_hd__and2b_2
X_6746_ _6746_/A vssd1 vssd1 vccd1 vccd1 _7498_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3958_ _8410_/Q _3877_/X _3962_/S vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__mux2_1
X_6677_ _6683_/A vssd1 vssd1 vccd1 vccd1 _6677_/X sky130_fd_sc_hd__buf_1
X_3889_ _8443_/Q vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__buf_2
X_5628_ _5628_/A vssd1 vssd1 vccd1 vccd1 _7916_/D sky130_fd_sc_hd__clkbuf_1
X_8416_ _8418_/CLK _8416_/D vssd1 vssd1 vccd1 vccd1 _8416_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3389_ clkbuf_0__3389_/X vssd1 vssd1 vccd1 vccd1 _6876__398/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5559_ _5581_/S vssd1 vssd1 vccd1 vccd1 _5572_/S sky130_fd_sc_hd__clkbuf_4
X_8347_ _8347_/CLK _8347_/D vssd1 vssd1 vccd1 vccd1 _8347_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3426_ _7045_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3426_/X sky130_fd_sc_hd__clkbuf_16
X_6884__404 _6885__405/A vssd1 vssd1 vccd1 vccd1 _8080_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8278_ _8278_/CLK _8278_/D vssd1 vssd1 vccd1 vccd1 _8278_/Q sky130_fd_sc_hd__dfxtp_1
X_7229_ _7229_/A vssd1 vssd1 vccd1 vccd1 _8287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6932__438 _6932__438/A vssd1 vssd1 vccd1 vccd1 _8116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _4932_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _4930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4861_ _4801_/X _7977_/Q _7881_/Q _4769_/X _4794_/A vssd1 vssd1 vccd1 vccd1 _4861_/X
+ sky130_fd_sc_hd__a221o_1
X_3812_ _8449_/Q vssd1 vssd1 vccd1 vccd1 _3812_/X sky130_fd_sc_hd__buf_2
X_4792_ _4757_/X _4788_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _4792_/X sky130_fd_sc_hd__o21a_1
X_7580_ _8435_/Q _7578_/X _7579_/X _7514_/X vssd1 vssd1 vccd1 vccd1 _8434_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6462_ _7848_/Q _7963_/Q _6466_/S vssd1 vssd1 vccd1 vccd1 _6463_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5413_ _5428_/S vssd1 vssd1 vccd1 vccd1 _5422_/S sky130_fd_sc_hd__clkbuf_2
X_8201_ _8201_/CLK _8201_/D vssd1 vssd1 vccd1 vccd1 _8201_/Q sky130_fd_sc_hd__dfxtp_1
X_6393_ _6393_/A vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__clkbuf_2
Xoutput123 _5994_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput112 _5972_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
Xoutput134 _5961_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
X_5344_ _5558_/A _5833_/A vssd1 vssd1 vccd1 vccd1 _5374_/S sky130_fd_sc_hd__or2_2
X_8132_ _8132_/CLK _8132_/D vssd1 vssd1 vccd1 vccd1 _8132_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput156 _5934_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput167 _5892_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
Xoutput145 _5912_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5275_ _8280_/Q _8001_/Q _5291_/S vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__mux2_1
Xoutput178 _6057_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput189 _6094_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
X_8063_ _8439_/CLK _8063_/D vssd1 vssd1 vccd1 vccd1 _8063_/Q sky130_fd_sc_hd__dfxtp_4
X_7014_ _7038_/A vssd1 vssd1 vccd1 vccd1 _7014_/X sky130_fd_sc_hd__buf_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _4248_/S vssd1 vssd1 vccd1 vccd1 _4239_/S sky130_fd_sc_hd__buf_2
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ _8349_/Q _4156_/X _4157_/S vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3390_ clkbuf_0__3390_/X vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__clkbuf_4
X_4088_ _4088_/A vssd1 vssd1 vccd1 vccd1 _8363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7916_ _7916_/CLK _7916_/D vssd1 vssd1 vccd1 vccd1 _7916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7847_ _8141_/CLK _7847_/D vssd1 vssd1 vccd1 vccd1 _7847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7778_ _7778_/CLK _7778_/D vssd1 vssd1 vccd1 vccd1 _7778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3409_ _6961_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3409_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7034__517 _7034__517/A vssd1 vssd1 vccd1 vccd1 _8198_/CLK sky130_fd_sc_hd__inv_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
Xinput36 wb_rst_i vssd1 vssd1 vccd1 vccd1 _6206_/A sky130_fd_sc_hd__buf_6
Xinput47 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__clkbuf_1
Xinput69 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_4
Xinput58 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6271__205 _6271__205/A vssd1 vssd1 vccd1 vccd1 _7797_/CLK sky130_fd_sc_hd__inv_2
X_5060_ _5060_/A vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__clkbuf_4
X_4011_ _8392_/Q _4010_/X _4011_/S vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5962_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5971_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7701_ _8016_/Q _7701_/B vssd1 vssd1 vccd1 vccd1 _7721_/S sky130_fd_sc_hd__and2_2
X_4913_ _5769_/S _4913_/B vssd1 vssd1 vccd1 vccd1 _8131_/D sky130_fd_sc_hd__nand2_1
X_5893_ _7699_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5894_/A sky130_fd_sc_hd__or2_1
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4844_ _4760_/X _7913_/Q _4814_/X _7921_/Q _4715_/X vssd1 vssd1 vccd1 vccd1 _4844_/X
+ sky130_fd_sc_hd__o221a_1
X_7410__165 _7410__165/A vssd1 vssd1 vccd1 vccd1 _8376_/CLK sky130_fd_sc_hd__inv_2
X_4775_ _4793_/A vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__clkbuf_2
X_7563_ _7563_/A vssd1 vssd1 vccd1 vccd1 _7563_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3226_ clkbuf_0__3226_/X vssd1 vssd1 vccd1 vccd1 _6534__255/A sky130_fd_sc_hd__clkbuf_4
X_7494_ _8488_/Q _7494_/B vssd1 vssd1 vccd1 vccd1 _7497_/B sky130_fd_sc_hd__xor2_1
X_6445_ _6445_/A vssd1 vssd1 vccd1 vccd1 _7840_/D sky130_fd_sc_hd__clkbuf_1
X_6376_ _8490_/Q _6390_/B _6387_/C vssd1 vssd1 vccd1 vccd1 _6376_/X sky130_fd_sc_hd__and3_1
X_8115_ _8115_/CLK _8115_/D vssd1 vssd1 vccd1 vccd1 _8115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5327_ _5327_/A vssd1 vssd1 vccd1 vccd1 _8074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8046_ _8046_/CLK _8046_/D vssd1 vssd1 vccd1 vccd1 _8046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7098__68 _7098__68/A vssd1 vssd1 vccd1 vccd1 _8249_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5258_ _8272_/Q _8009_/Q _5261_/S vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3442_ clkbuf_0__3442_/X vssd1 vssd1 vccd1 vccd1 _7128__92/A sky130_fd_sc_hd__clkbuf_4
X_5189_ _5292_/B vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__buf_2
X_4209_ _8331_/Q _4138_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6671__321 _6672__322/A vssd1 vssd1 vccd1 vccd1 _7985_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7353__119 _7354__120/A vssd1 vssd1 vccd1 vccd1 _8330_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6977__471 _6979__473/A vssd1 vssd1 vccd1 vccd1 _8152_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _8163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4491_ _4491_/A vssd1 vssd1 vccd1 vccd1 _8192_/D sky130_fd_sc_hd__clkbuf_1
X_6230_ _6230_/A vssd1 vssd1 vccd1 vccd1 _7773_/D sky130_fd_sc_hd__clkbuf_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6161_/A vssd1 vssd1 vccd1 vccd1 _6161_/X sky130_fd_sc_hd__clkbuf_2
X_6945__448 _6947__450/A vssd1 vssd1 vccd1 vccd1 _8127_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5112_ _8173_/Q _8149_/Q _8411_/Q _8181_/Q _5123_/A _5111_/X vssd1 vssd1 vccd1 vccd1
+ _5112_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _7753_/Q _6111_/A vssd1 vssd1 vccd1 vccd1 _6092_/X sky130_fd_sc_hd__or2_1
X_5043_ _5111_/A vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__buf_2
XFILLER_111_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5945_ _5945_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__and2_1
XFILLER_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5876_ _7597_/A _5884_/B vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__or2_1
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _8351_/Q _4619_/A _4790_/X _8327_/Q _4659_/A vssd1 vssd1 vccd1 vccd1 _4827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7615_ _7615_/A _7615_/B _7615_/C vssd1 vssd1 vccd1 vccd1 _7616_/A sky130_fd_sc_hd__and3_1
X_4758_ _4749_/X _7803_/Q _7728_/Q _4753_/X _4757_/X vssd1 vssd1 vccd1 vccd1 _4758_/X
+ sky130_fd_sc_hd__a221o_1
X_7546_ _7546_/A _7546_/B vssd1 vssd1 vccd1 vccd1 _8425_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7477_ _7477_/A _7477_/B _7477_/C _6777_/B vssd1 vssd1 vccd1 vccd1 _7477_/X sky130_fd_sc_hd__or4b_1
X_4689_ _8331_/Q _8221_/Q _7878_/Q _8355_/Q _4650_/X _4651_/X vssd1 vssd1 vccd1 vccd1
+ _4689_/X sky130_fd_sc_hd__mux4_1
X_6428_ _6428_/A vssd1 vssd1 vccd1 vccd1 _7832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _6359_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8029_ _8029_/CLK _8029_/D vssd1 vssd1 vccd1 vccd1 _8029_/Q sky130_fd_sc_hd__dfxtp_1
X_8521__220 vssd1 vssd1 vccd1 vccd1 _8521__220/HI core0Index[7] sky130_fd_sc_hd__conb_1
Xclkbuf_1_0_0__3425_ clkbuf_0__3425_/X vssd1 vssd1 vccd1 vccd1 _7057_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3287_ clkbuf_0__3287_/X vssd1 vssd1 vccd1 vccd1 _6824__370/A sky130_fd_sc_hd__clkbuf_4
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _8449_/Q vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__buf_2
XFILLER_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _5730_/A vssd1 vssd1 vccd1 vccd1 _7871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5661_ _5565_/X _7901_/Q _5665_/S vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__mux2_1
X_6951__452 _6954__455/A vssd1 vssd1 vccd1 vccd1 _8131_/CLK sky130_fd_sc_hd__inv_2
X_5592_ _5592_/A vssd1 vssd1 vccd1 vccd1 _7932_/D sky130_fd_sc_hd__clkbuf_1
X_8380_ _8380_/CLK _8380_/D vssd1 vssd1 vccd1 vccd1 _8380_/Q sky130_fd_sc_hd__dfxtp_1
X_4612_ _4613_/A vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__clkbuf_2
X_4543_ _8170_/Q _4445_/X _4543_/S vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3390_ _6879_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3390_/X sky130_fd_sc_hd__clkbuf_16
X_7331_ _7331_/A vssd1 vssd1 vccd1 vccd1 _7331_/X sky130_fd_sc_hd__clkbuf_2
X_7047__527 _7048__528/A vssd1 vssd1 vccd1 vccd1 _8208_/CLK sky130_fd_sc_hd__inv_2
X_7262_ _7262_/A _7262_/B vssd1 vssd1 vccd1 vccd1 _7262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ _4474_/A vssd1 vssd1 vccd1 vccd1 _8199_/D sky130_fd_sc_hd__clkbuf_1
X_6213_ _7603_/A _7767_/Q _6217_/S vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__mux2_1
X_7193_ _8309_/Q _7193_/B _7193_/C _7193_/D vssd1 vssd1 vccd1 vccd1 _7195_/A sky130_fd_sc_hd__nand4_1
XFILLER_97_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6144_ _6206_/A vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__clkbuf_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_16 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6075_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6075_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_38 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_49 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_27 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__clkbuf_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3758_ clkbuf_0__3758_/X vssd1 vssd1 vccd1 vccd1 _7643__49/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5928_ _5928_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__or2_4
XFILLER_110_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5859_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5866_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7529_ _7534_/A _7529_/B vssd1 vssd1 vccd1 vccd1 _8418_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7449__21 _7450__22/A vssd1 vssd1 vccd1 vccd1 _8407_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3408_ clkbuf_0__3408_/X vssd1 vssd1 vccd1 vccd1 _6957__457/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6523__246 _6524__247/A vssd1 vssd1 vccd1 vccd1 _7886_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6684__331 _6685__332/A vssd1 vssd1 vccd1 vccd1 _7995_/CLK sky130_fd_sc_hd__inv_2
X_4190_ _4190_/A vssd1 vssd1 vccd1 vccd1 _8337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6829__374 _6830__375/A vssd1 vssd1 vccd1 vccd1 _8042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7880_ _7880_/CLK _7880_/D vssd1 vssd1 vccd1 vccd1 _7880_/Q sky130_fd_sc_hd__dfxtp_1
X_6831_ _6879_/A vssd1 vssd1 vccd1 vccd1 _6831_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3612_ clkbuf_0__3612_/X vssd1 vssd1 vccd1 vccd1 _7380_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _3989_/S vssd1 vssd1 vccd1 vccd1 _3983_/S sky130_fd_sc_hd__buf_2
X_6762_ _6789_/A _6789_/B _6789_/C _8422_/Q vssd1 vssd1 vccd1 vccd1 _7465_/C sky130_fd_sc_hd__a31o_1
X_7366__129 _7366__129/A vssd1 vssd1 vccd1 vccd1 _8340_/CLK sky130_fd_sc_hd__inv_2
X_5713_ _4138_/X _7878_/Q _5719_/S vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__mux2_1
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _7909_/D sky130_fd_sc_hd__clkbuf_1
X_8432_ _8433_/CLK _8432_/D vssd1 vssd1 vccd1 vccd1 _8432_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3442_ _7126_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3442_/X sky130_fd_sc_hd__clkbuf_16
X_8363_ _8363_/CLK _8363_/D vssd1 vssd1 vccd1 vccd1 _8363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5575_ _5574_/X _7938_/Q _5581_/S vssd1 vssd1 vccd1 vccd1 _5576_/A sky130_fd_sc_hd__mux2_1
X_7314_ _7315_/A _7321_/B _7313_/X _7248_/X vssd1 vssd1 vccd1 vccd1 _8313_/D sky130_fd_sc_hd__o211a_1
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4526_ _4526_/A vssd1 vssd1 vccd1 vccd1 _8178_/D sky130_fd_sc_hd__clkbuf_1
X_8294_ _8294_/CLK _8294_/D vssd1 vssd1 vccd1 vccd1 _8294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ _4457_/A _5797_/A vssd1 vssd1 vccd1 vccd1 _4473_/S sky130_fd_sc_hd__or2_4
X_7245_ _7237_/X _7238_/Y _7240_/X _7243_/X _7244_/X vssd1 vssd1 vccd1 vccd1 _7246_/D
+ sky130_fd_sc_hd__o2111a_1
X_7176_ _7176_/A _7193_/C _7217_/C vssd1 vssd1 vccd1 vccd1 _7216_/B sky130_fd_sc_hd__and3_1
X_4388_ _4342_/X _8230_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__mux2_1
X_6127_ _6025_/B _7855_/Q _6125_/X _6126_/X _6037_/A vssd1 vssd1 vccd1 vccd1 _6127_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6058_ _7819_/Q input5/X _6058_/S vssd1 vssd1 vccd1 vccd1 _6058_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _8093_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6249__187 _6249__187/A vssd1 vssd1 vccd1 vccd1 _7779_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6958__458 _6960__460/A vssd1 vssd1 vccd1 vccd1 _8137_/CLK sky130_fd_sc_hd__inv_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5360_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _8261_/D sky130_fd_sc_hd__clkbuf_1
X_5291_ _7984_/Q _8019_/Q _5291_/S vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4242_ _8291_/Q _4241_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4243_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4173_ _8342_/Q _4018_/X _4175_/S vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__mux2_1
X_7443__16 _7445__18/A vssd1 vssd1 vccd1 vccd1 _8402_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7932_ _7932_/CLK _7932_/D vssd1 vssd1 vccd1 vccd1 _7932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7863_ _7863_/CLK _7863_/D vssd1 vssd1 vccd1 vccd1 _7863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7794_ _7794_/CLK _7794_/D vssd1 vssd1 vccd1 vccd1 _7794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6814_ _8414_/Q vssd1 vssd1 vccd1 vccd1 _7508_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3957_ _3957_/A vssd1 vssd1 vccd1 vccd1 _8411_/D sky130_fd_sc_hd__clkbuf_1
X_6745_ _8428_/Q _6745_/B vssd1 vssd1 vccd1 vccd1 _6746_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6676_ _6676_/A vssd1 vssd1 vccd1 vccd1 _6676_/X sky130_fd_sc_hd__buf_1
X_3888_ _3888_/A vssd1 vssd1 vccd1 vccd1 _8468_/D sky130_fd_sc_hd__clkbuf_1
X_8415_ _8418_/CLK _8415_/D vssd1 vssd1 vccd1 vccd1 _8415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5627_ _7916_/Q _4984_/X _5629_/S vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__mux2_1
X_5558_ _5558_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5581_/S sky130_fd_sc_hd__or2_2
X_8346_ _8346_/CLK _8346_/D vssd1 vssd1 vccd1 vccd1 _8346_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3425_ _7044_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3425_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8277_ _8277_/CLK _8277_/D vssd1 vssd1 vccd1 vccd1 _8277_/Q sky130_fd_sc_hd__dfxtp_1
X_4509_ _8185_/Q _4241_/X _4513_/S vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5489_ _5489_/A vssd1 vssd1 vccd1 vccd1 _7998_/D sky130_fd_sc_hd__clkbuf_1
X_7228_ _7331_/A _7228_/B _7228_/C vssd1 vssd1 vccd1 vccd1 _7229_/A sky130_fd_sc_hd__and3_1
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3287_ _6732_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3287_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7159_ _8486_/Q _7159_/B vssd1 vssd1 vccd1 vccd1 _7236_/C sky130_fd_sc_hd__xor2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6971__466 _6973__468/A vssd1 vssd1 vccd1 vccd1 _8147_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8501__251 vssd1 vssd1 vccd1 vccd1 partID[0] _8501__251/LO sky130_fd_sc_hd__conb_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4860_ _4932_/B _4858_/X _4859_/X vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4791_ _8186_/Q _4789_/X _4790_/X _8162_/Q _4663_/A vssd1 vssd1 vccd1 vccd1 _4791_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461_ _6461_/A vssd1 vssd1 vccd1 vccd1 _7847_/D sky130_fd_sc_hd__clkbuf_1
X_6536__256 _6539__259/A vssd1 vssd1 vccd1 vccd1 _7896_/CLK sky130_fd_sc_hd__inv_2
X_8200_ _8200_/CLK _8200_/D vssd1 vssd1 vccd1 vccd1 _8200_/Q sky130_fd_sc_hd__dfxtp_1
X_5412_ _5412_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5428_/S sky130_fd_sc_hd__or2_2
X_6392_ _7821_/Q _6383_/X _6371_/X _6390_/X _6391_/X vssd1 vssd1 vccd1 vccd1 _7821_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput124 _5996_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput113 _5975_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _5557_/A vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__buf_2
X_8131_ _8131_/CLK _8131_/D vssd1 vssd1 vccd1 vccd1 _8131_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput157 _5936_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput135 _5964_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
Xoutput146 _5914_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput168 _5894_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5274_ _5295_/A _5272_/X _5273_/X vssd1 vssd1 vccd1 vccd1 _5278_/B sky130_fd_sc_hd__o21ai_1
Xoutput179 _6060_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
X_8062_ _8439_/CLK _8062_/D vssd1 vssd1 vccd1 vccd1 _8062_/Q sky130_fd_sc_hd__dfxtp_4
X_7013_ _7013_/A vssd1 vssd1 vccd1 vccd1 _7013_/X sky130_fd_sc_hd__buf_1
X_4225_ _5539_/A _5558_/A vssd1 vssd1 vccd1 vccd1 _4248_/S sky130_fd_sc_hd__nor2_2
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _8060_/Q vssd1 vssd1 vccd1 vccd1 _4156_/X sky130_fd_sc_hd__buf_2
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4087_ _8363_/Q _3998_/X _4093_/S vssd1 vssd1 vccd1 vccd1 _4088_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7915_ _7915_/CLK _7915_/D vssd1 vssd1 vccd1 vccd1 _7915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7846_ _8483_/CLK _7846_/D vssd1 vssd1 vccd1 vccd1 _7846_/Q sky130_fd_sc_hd__dfxtp_1
X_7777_ _7777_/CLK _7777_/D vssd1 vssd1 vccd1 vccd1 _7777_/Q sky130_fd_sc_hd__dfxtp_1
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _8100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6659_ _6659_/A vssd1 vssd1 vccd1 vccd1 _7975_/D sky130_fd_sc_hd__clkbuf_1
X_8329_ _8329_/CLK _8329_/D vssd1 vssd1 vccd1 vccd1 _8329_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3408_ _6955_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3408_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__clkbuf_4
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
Xinput37 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _5945_/A sky130_fd_sc_hd__buf_4
XFILLER_116_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput48 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _5947_/A sky130_fd_sc_hd__buf_4
Xinput59 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__buf_4
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4010_ _4356_/A vssd1 vssd1 vccd1 vccd1 _4010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5961_ _5961_/A vssd1 vssd1 vccd1 vccd1 _5961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7700_ _7698_/Y _7699_/Y _6194_/X vssd1 vssd1 vccd1 vccd1 _8491_/D sky130_fd_sc_hd__a21oi_1
X_4912_ _4911_/X _6852_/B _4999_/A vssd1 vssd1 vccd1 vccd1 _4913_/B sky130_fd_sc_hd__nand3b_1
X_5892_ _5892_/A vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__clkbuf_1
X_4843_ _4749_/X _7801_/Q _7726_/Q _4795_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4843_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4774_ _4758_/X _4763_/X _4772_/X _4928_/B vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__a211o_1
X_7562_ _7584_/B _6820_/C _7556_/X vssd1 vssd1 vccd1 vccd1 _7562_/Y sky130_fd_sc_hd__a21oi_1
X_7493_ _6359_/X _6763_/Y _7492_/Y _6803_/A _6803_/B vssd1 vssd1 vccd1 vccd1 _7500_/B
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_1_1_0__3225_ clkbuf_0__3225_/X vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__clkbuf_4
X_6444_ _7840_/Q _5969_/A _6444_/S vssd1 vssd1 vccd1 vccd1 _6445_/A sky130_fd_sc_hd__mux2_1
X_6375_ _7672_/A vssd1 vssd1 vccd1 vccd1 _6387_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8114_ _8114_/CLK _8114_/D vssd1 vssd1 vccd1 vccd1 _8114_/Q sky130_fd_sc_hd__dfxtp_1
X_5326_ _5321_/B _5326_/B _7604_/A vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__and3b_1
X_8045_ _8045_/CLK _8045_/D vssd1 vssd1 vccd1 vccd1 _8045_/Q sky130_fd_sc_hd__dfxtp_1
X_5257_ _5220_/X _5255_/X _5256_/X vssd1 vssd1 vccd1 vccd1 _5257_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _8332_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3441_ clkbuf_0__3441_/X vssd1 vssd1 vccd1 vccd1 _7125__90/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5188_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5292_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _8355_/Q _4138_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4140_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7829_ _8489_/CLK _7829_/D vssd1 vssd1 vccd1 vccd1 _7829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7040__522 _7043__525/A vssd1 vssd1 vccd1 vccd1 _8203_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6823__369 _6824__370/A vssd1 vssd1 vccd1 vccd1 _8037_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4490_ _8192_/Q _4244_/X _4492_/S vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6159_/X _7768_/Q _6149_/X _6153_/X _7736_/Q vssd1 vssd1 vccd1 vccd1 _7736_/D
+ sky130_fd_sc_hd__o32a_1
X_6984__476 _6985__477/A vssd1 vssd1 vccd1 vccd1 _8157_/CLK sky130_fd_sc_hd__inv_2
X_5111_ _5111_/A vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _7828_/Q input15/X _6107_/A vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__mux2_1
X_5042_ _5164_/A vssd1 vssd1 vccd1 vccd1 _5111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5944_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5875_ _5943_/B vssd1 vssd1 vccd1 vccd1 _5884_/B sky130_fd_sc_hd__clkbuf_2
X_4826_ _8217_/Q _4770_/X _4787_/X _7874_/Q vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__a22o_1
X_7614_ _7614_/A vssd1 vssd1 vccd1 vccd1 _8448_/D sky130_fd_sc_hd__clkbuf_1
X_7545_ _8425_/Q _7530_/X _7544_/X _7461_/B vssd1 vssd1 vccd1 vccd1 _7546_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4757_/A vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__buf_2
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4688_ _8165_/Q _8157_/Q _8119_/Q _8189_/Q _4648_/X _4640_/X vssd1 vssd1 vccd1 vccd1
+ _4688_/X sky130_fd_sc_hd__mux4_2
X_7476_ _8496_/Q _7476_/B _7476_/C vssd1 vssd1 vccd1 vccd1 _7477_/C sky130_fd_sc_hd__and3b_1
X_6427_ _7832_/Q _5952_/A _6433_/S vssd1 vssd1 vccd1 vccd1 _6428_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6358_ _6289_/X _6356_/X _6357_/X vssd1 vssd1 vccd1 vccd1 _7814_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _5220_/A _5307_/X _5308_/X _5062_/A vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6289_ _6289_/A vssd1 vssd1 vccd1 vccd1 _6289_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8028_ _8028_/CLK _8028_/D vssd1 vssd1 vccd1 vccd1 _8028_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3424_ clkbuf_0__3424_/X vssd1 vssd1 vccd1 vccd1 _7041__523/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3286_ clkbuf_0__3286_/X vssd1 vssd1 vccd1 vccd1 _6728__362/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8017_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7005__494 _7006__495/A vssd1 vssd1 vccd1 vccd1 _8175_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _3990_/A vssd1 vssd1 vccd1 vccd1 _8397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _7902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _8142_/Q vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__inv_2
X_5591_ _5568_/X _7932_/Q _5593_/S vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__mux2_1
X_4542_ _4542_/A vssd1 vssd1 vccd1 vccd1 _8171_/D sky130_fd_sc_hd__clkbuf_1
X_7330_ _8317_/Q _7337_/B vssd1 vssd1 vccd1 vccd1 _7330_/X sky130_fd_sc_hd__or2_1
X_4473_ _4365_/X _8199_/Q _4473_/S vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__mux2_1
X_7261_ _8482_/Q _7261_/B vssd1 vssd1 vccd1 vccd1 _7262_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6212_ _6212_/A vssd1 vssd1 vccd1 vccd1 _7766_/D sky130_fd_sc_hd__clkbuf_1
X_7192_ _7471_/A _7192_/B vssd1 vssd1 vccd1 vccd1 _7192_/Y sky130_fd_sc_hd__xnor2_1
X_8544__243 vssd1 vssd1 vccd1 vccd1 _8544__243/HI partID[9] sky130_fd_sc_hd__conb_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _7748_/Q _6082_/B vssd1 vssd1 vccd1 vccd1 _6074_/X sky130_fd_sc_hd__or2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_39 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_28 _6096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_17 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _5025_/A _7323_/A vssd1 vssd1 vccd1 vccd1 _5139_/A sky130_fd_sc_hd__nor2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3757_ clkbuf_0__3757_/X vssd1 vssd1 vccd1 vccd1 _7635__42/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6976_ _6976_/A vssd1 vssd1 vccd1 vccd1 _6976_/X sky130_fd_sc_hd__buf_1
X_5927_ _5927_/A vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5858_ _5868_/A vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__buf_2
X_5789_ _7795_/Q _4356_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__mux2_1
X_4809_ _4721_/X _4792_/X _4800_/X _4808_/X _4622_/X vssd1 vssd1 vccd1 vccd1 _4809_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7528_ _8418_/Q _7522_/X _7527_/X _6785_/B vssd1 vssd1 vccd1 vccd1 _7529_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ _7459_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _7460_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3407_ clkbuf_0__3407_/X vssd1 vssd1 vccd1 vccd1 _6952__453/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8528__227 vssd1 vssd1 vccd1 vccd1 _8528__227/HI core1Index[7] sky130_fd_sc_hd__conb_1
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3611_ clkbuf_0__3611_/X vssd1 vssd1 vccd1 vccd1 _7356__121/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_110 _7597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7053__532 _7054__533/A vssd1 vssd1 vccd1 vccd1 _8213_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6761_ _8422_/Q _6789_/A _6786_/B _6789_/C vssd1 vssd1 vccd1 vccd1 _7465_/B sky130_fd_sc_hd__nand4_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3973_ _4515_/A _5797_/B vssd1 vssd1 vccd1 vccd1 _3989_/S sky130_fd_sc_hd__or2_2
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5712_ _5712_/A vssd1 vssd1 vccd1 vccd1 _7879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5643_ _5565_/X _7909_/Q _5647_/S vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__mux2_1
X_6836__379 _6836__379/A vssd1 vssd1 vccd1 vccd1 _8047_/CLK sky130_fd_sc_hd__inv_2
X_8431_ _8433_/CLK _8431_/D vssd1 vssd1 vccd1 vccd1 _8431_/Q sky130_fd_sc_hd__dfxtp_1
X_5574_ _5574_/A vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3441_ _7120_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3441_/X sky130_fd_sc_hd__clkbuf_16
X_8362_ _8362_/CLK _8362_/D vssd1 vssd1 vccd1 vccd1 _8362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4525_ _4356_/X _8178_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__mux2_1
X_7313_ _7247_/A _7262_/A _7311_/Y _7317_/B vssd1 vssd1 vccd1 vccd1 _7313_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8293_ _8293_/CLK _8293_/D vssd1 vssd1 vccd1 vccd1 _8293_/Q sky130_fd_sc_hd__dfxtp_1
X_4456_ _4456_/A vssd1 vssd1 vccd1 vccd1 _8207_/D sky130_fd_sc_hd__clkbuf_1
X_7244_ _7692_/A _7178_/B _7218_/X vssd1 vssd1 vccd1 vccd1 _7244_/X sky130_fd_sc_hd__o21a_1
X_4387_ _4402_/S vssd1 vssd1 vccd1 vccd1 _4396_/S sky130_fd_sc_hd__buf_2
X_7175_ _8306_/Q _7184_/A vssd1 vssd1 vccd1 vccd1 _7217_/C sky130_fd_sc_hd__and2_1
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6126_ _7830_/Q _6129_/C _6008_/A vssd1 vssd1 vccd1 vccd1 _6126_/X sky130_fd_sc_hd__a21o_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6585__296 _6588__299/A vssd1 vssd1 vccd1 vccd1 _7936_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6057_ _6053_/X _6054_/X _6055_/X _6056_/X vssd1 vssd1 vccd1 vccd1 _6057_/X sky130_fd_sc_hd__o211a_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _4416_/X _8093_/Q _5010_/S vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__mux2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6605__311 _6605__311/A vssd1 vssd1 vccd1 vccd1 _7951_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__3550_ clkbuf_0__3550_/X vssd1 vssd1 vccd1 vccd1 _7348__115/A sky130_fd_sc_hd__clkbuf_16
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4310_ _8261_/Q _4182_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__mux2_1
X_5290_ _5048_/X _5286_/X _5289_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__a211o_1
XFILLER_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4241_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _4241_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _8343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7931_ _7931_/CLK _7931_/D vssd1 vssd1 vccd1 vccd1 _7931_/Q sky130_fd_sc_hd__dfxtp_1
X_7372__134 _7373__135/A vssd1 vssd1 vccd1 vccd1 _8345_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7862_ _7862_/CLK _7862_/D vssd1 vssd1 vccd1 vccd1 _7862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7793_ _7793_/CLK _7793_/D vssd1 vssd1 vccd1 vccd1 _7793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6813_ _7499_/A _7499_/B _6813_/C _6813_/D vssd1 vssd1 vccd1 vccd1 _6816_/C sky130_fd_sc_hd__and4_1
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3956_ _8411_/Q _3874_/X _3962_/S vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__mux2_1
X_6744_ _8484_/Q _7557_/A vssd1 vssd1 vccd1 vccd1 _7500_/A sky130_fd_sc_hd__xor2_1
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5626_ _5626_/A vssd1 vssd1 vccd1 vccd1 _7917_/D sky130_fd_sc_hd__clkbuf_1
X_3887_ _8468_/Q _3886_/X _3893_/S vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__mux2_1
X_8414_ _8430_/CLK _8414_/D vssd1 vssd1 vccd1 vccd1 _8414_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3424_ _7038_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3424_/X sky130_fd_sc_hd__clkbuf_16
X_5557_ _5557_/A vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8345_ _8345_/CLK _8345_/D vssd1 vssd1 vccd1 vccd1 _8345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8276_ _8276_/CLK _8276_/D vssd1 vssd1 vccd1 vccd1 _8276_/Q sky130_fd_sc_hd__dfxtp_1
X_5488_ _5349_/X _7998_/Q _5494_/S vssd1 vssd1 vccd1 vccd1 _5489_/A sky130_fd_sc_hd__mux2_1
X_4508_ _4508_/A vssd1 vssd1 vccd1 vccd1 _8186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4439_ _8447_/Q vssd1 vssd1 vccd1 vccd1 _4439_/X sky130_fd_sc_hd__clkbuf_4
X_7227_ _7320_/C _7262_/A vssd1 vssd1 vccd1 vccd1 _7228_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3286_ _6726_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3286_/X sky130_fd_sc_hd__clkbuf_16
X_6255__192 _6258__195/A vssd1 vssd1 vccd1 vccd1 _7784_/CLK sky130_fd_sc_hd__inv_2
X_7158_ _8310_/Q _7158_/B vssd1 vssd1 vccd1 vccd1 _7159_/B sky130_fd_sc_hd__xnor2_1
X_7089_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7089_/X sky130_fd_sc_hd__buf_1
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6109_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4790_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3241_ clkbuf_0__3241_/X vssd1 vssd1 vccd1 vccd1 _6605__311/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _7847_/Q _7962_/Q _6466_/S vssd1 vssd1 vccd1 vccd1 _6461_/A sky130_fd_sc_hd__mux2_1
X_5411_ _5411_/A vssd1 vssd1 vccd1 vccd1 _8036_/D sky130_fd_sc_hd__clkbuf_1
X_6391_ _6391_/A vssd1 vssd1 vccd1 vccd1 _6391_/X sky130_fd_sc_hd__clkbuf_2
Xoutput125 _6001_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput114 _5977_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
X_5342_ _8067_/Q vssd1 vssd1 vccd1 vccd1 _5557_/A sky130_fd_sc_hd__buf_2
X_8130_ _8130_/CLK _8130_/D vssd1 vssd1 vccd1 vccd1 _8130_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput158 _5938_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput136 _5966_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput147 _5916_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
X_8061_ _8439_/CLK _8061_/D vssd1 vssd1 vccd1 vccd1 _8061_/Q sky130_fd_sc_hd__dfxtp_4
Xoutput169 _5896_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _8451_/Q _5227_/A _5292_/B _8459_/Q _5108_/A vssd1 vssd1 vccd1 vccd1 _5273_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ _5538_/A _4475_/B _5538_/B vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__or3b_2
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4155_ _4155_/A vssd1 vssd1 vccd1 vccd1 _8350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4086_/A vssd1 vssd1 vccd1 vccd1 _8364_/D sky130_fd_sc_hd__clkbuf_1
X_7914_ _7914_/CLK _7914_/D vssd1 vssd1 vccd1 vccd1 _7914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697__342 _6698__343/A vssd1 vssd1 vccd1 vccd1 _8006_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7845_ _8141_/CLK _7845_/D vssd1 vssd1 vccd1 vccd1 _7845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7776_ _7776_/CLK _7776_/D vssd1 vssd1 vccd1 vccd1 _7776_/Q sky130_fd_sc_hd__dfxtp_1
X_4988_ _8100_/Q _4987_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__mux2_1
X_3939_ _3939_/A vssd1 vssd1 vccd1 vccd1 _8452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3439_ clkbuf_0__3439_/X vssd1 vssd1 vccd1 vccd1 _7113__80/A sky130_fd_sc_hd__clkbuf_4
X_6658_ _7975_/Q _5943_/A _6658_/S vssd1 vssd1 vccd1 vccd1 _6659_/A sky130_fd_sc_hd__mux2_1
X_5609_ _5568_/X _7924_/Q _5611_/S vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__mux2_1
X_8328_ _8328_/CLK _8328_/D vssd1 vssd1 vccd1 vccd1 _8328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3407_ _6949_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3407_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8259_ _8259_/CLK _8259_/D vssd1 vssd1 vccd1 vccd1 _8259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _6123_/A sky130_fd_sc_hd__clkbuf_4
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _3842_/D sky130_fd_sc_hd__clkbuf_1
Xinput38 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__buf_4
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6908__420 _6908__420/A vssd1 vssd1 vccd1 vccd1 _8098_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _5960_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__and2_1
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _7615_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__or2_1
X_6542__261 _6544__263/A vssd1 vssd1 vccd1 vccd1 _7901_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4999_/B _4911_/B _4911_/C vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__and3_1
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ _4422_/X _4610_/A _4840_/X _4841_/X vssd1 vssd1 vccd1 vccd1 _8135_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _4773_/A vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__buf_2
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7561_ _8431_/Q vssd1 vssd1 vccd1 vccd1 _7563_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7492_ _7492_/A _7492_/B vssd1 vssd1 vccd1 vccd1 _7492_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3224_ clkbuf_0__3224_/X vssd1 vssd1 vccd1 vccd1 _6524__247/A sky130_fd_sc_hd__clkbuf_4
X_6443_ _6443_/A vssd1 vssd1 vccd1 vccd1 _7839_/D sky130_fd_sc_hd__clkbuf_1
X_6374_ _8017_/Q vssd1 vssd1 vccd1 vccd1 _7672_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8113_ _8113_/CLK _8113_/D vssd1 vssd1 vccd1 vccd1 _8113_/Q sky130_fd_sc_hd__dfxtp_1
X_5325_ _6892_/A vssd1 vssd1 vccd1 vccd1 _7604_/A sky130_fd_sc_hd__clkbuf_2
X_8508__258 vssd1 vssd1 vccd1 vccd1 partID[14] _8508__258/LO sky130_fd_sc_hd__conb_1
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8044_ _8044_/CLK _8044_/D vssd1 vssd1 vccd1 vccd1 _8044_/Q sky130_fd_sc_hd__dfxtp_1
X_5256_ _8176_/Q _5214_/X _5189_/X _8168_/Q _5038_/A vssd1 vssd1 vccd1 vccd1 _5256_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3440_ clkbuf_0__3440_/X vssd1 vssd1 vccd1 vccd1 _7118__84/A sky130_fd_sc_hd__clkbuf_4
X_4207_ _8332_/Q _4101_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__mux2_1
X_5187_ _5187_/A _5187_/B vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__or2_1
X_4138_ _8066_/Q vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4069_ _3925_/X _8371_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7828_ _8483_/CLK _7828_/D vssd1 vssd1 vccd1 vccd1 _7828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7759_ _8441_/CLK _7759_/D vssd1 vssd1 vccd1 vccd1 _7759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5110_ _5160_/A _5110_/B vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__and2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6072_/X _6088_/X _6089_/X _6075_/X vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__o211a_1
XFILLER_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5041_ _5291_/S vssd1 vssd1 vccd1 vccd1 _5269_/S sky130_fd_sc_hd__buf_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__or2_1
X_7017__503 _7019__505/A vssd1 vssd1 vccd1 vccd1 _8184_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5874_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4825_ _4820_/X _4821_/X _4824_/X _4673_/X vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__a211o_1
X_7613_ _7707_/A _7615_/B _7613_/C vssd1 vssd1 vccd1 vccd1 _7614_/A sky130_fd_sc_hd__and3_1
X_7544_ _7544_/A vssd1 vssd1 vccd1 vccd1 _7544_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4756_ _4793_/A vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__buf_2
X_4687_ _4930_/B _4684_/X _4686_/X vssd1 vssd1 vccd1 vccd1 _4687_/X sky130_fd_sc_hd__a21o_1
X_7475_ _7476_/B _7476_/C _7200_/A vssd1 vssd1 vccd1 vccd1 _7477_/B sky130_fd_sc_hd__a21boi_1
X_6426_ _6426_/A vssd1 vssd1 vccd1 vccd1 _7831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6357_ _7814_/Q _6401_/A _6192_/X vssd1 vssd1 vccd1 vccd1 _6357_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5308_ _8231_/Q _5227_/A _5215_/A _8466_/Q vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__o22a_1
XFILLER_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6288_ _7654_/B vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6549__267 _6549__267/A vssd1 vssd1 vccd1 vccd1 _7907_/CLK sky130_fd_sc_hd__inv_2
X_8027_ _8027_/CLK _8027_/D vssd1 vssd1 vccd1 vccd1 _8027_/Q sky130_fd_sc_hd__dfxtp_1
X_5239_ _8391_/Q _5239_/B vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__or2_1
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3423_ clkbuf_0__3423_/X vssd1 vssd1 vccd1 vccd1 _7037__520/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3285_ clkbuf_0__3285_/X vssd1 vssd1 vccd1 vccd1 _6725__360/A sky130_fd_sc_hd__clkbuf_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6990__481 _6991__482/A vssd1 vssd1 vccd1 vccd1 _8162_/CLK sky130_fd_sc_hd__inv_2
X_4610_ _4610_/A vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__clkbuf_2
X_5590_ _5590_/A vssd1 vssd1 vccd1 vccd1 _7933_/D sky130_fd_sc_hd__clkbuf_1
X_4541_ _8171_/Q _4442_/X _4543_/S vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4472_ _4472_/A vssd1 vssd1 vccd1 vccd1 _8200_/D sky130_fd_sc_hd__clkbuf_1
X_7260_ _8288_/Q _8287_/Q vssd1 vssd1 vccd1 vccd1 _7261_/B sky130_fd_sc_hd__or2_2
X_6211_ _7600_/A _7766_/Q _6217_/S vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__mux2_1
X_7191_ _7191_/A _7191_/B vssd1 vssd1 vccd1 vccd1 _7192_/B sky130_fd_sc_hd__nand2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6073_ _7823_/Q input9/X _6077_/S vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__mux2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_29 _6108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_18 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5025_/A vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3756_ clkbuf_0__3756_/X vssd1 vssd1 vccd1 vccd1 _7632__40/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5926_ _5926_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__or2_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5857_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__inv_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5788_ _5788_/A vssd1 vssd1 vccd1 vccd1 _7796_/D sky130_fd_sc_hd__clkbuf_1
X_4808_ _4802_/X _4804_/X _4807_/X _4644_/X vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ _8101_/Q _8056_/Q _7940_/Q _8293_/Q _4669_/X _4670_/X vssd1 vssd1 vccd1 vccd1
+ _4739_/X sky130_fd_sc_hd__mux4_1
X_7527_ _7544_/A vssd1 vssd1 vccd1 vccd1 _7527_/X sky130_fd_sc_hd__clkbuf_2
X_7458_ _8484_/Q _7458_/B vssd1 vssd1 vccd1 vccd1 _7487_/A sky130_fd_sc_hd__xnor2_1
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6409_ _7826_/Q _6401_/X _6393_/X _6408_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _7826_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3406_ clkbuf_0__3406_/X vssd1 vssd1 vccd1 vccd1 _6976_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__3421_ clkbuf_0__3421_/X vssd1 vssd1 vccd1 vccd1 _7025__510/A sky130_fd_sc_hd__clkbuf_16
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6597__305 _6597__305/A vssd1 vssd1 vccd1 vccd1 _7945_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_100 _3931_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0__3610_ clkbuf_0__3610_/X vssd1 vssd1 vccd1 vccd1 _7354__120/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6760_ _8420_/Q _8419_/Q vssd1 vssd1 vccd1 vccd1 _6789_/C sky130_fd_sc_hd__and2_1
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3972_ _4287_/B _3972_/B _4287_/A vssd1 vssd1 vccd1 vccd1 _5797_/B sky130_fd_sc_hd__or3b_4
X_5711_ _4101_/X _7879_/Q _5719_/S vssd1 vssd1 vccd1 vccd1 _5712_/A sky130_fd_sc_hd__mux2_1
X_5642_ _5642_/A vssd1 vssd1 vccd1 vccd1 _7910_/D sky130_fd_sc_hd__clkbuf_1
X_6691__337 _6692__338/A vssd1 vssd1 vccd1 vccd1 _8001_/CLK sky130_fd_sc_hd__inv_2
X_8430_ _8430_/CLK _8430_/D vssd1 vssd1 vccd1 vccd1 _8430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5573_ _5573_/A vssd1 vssd1 vccd1 vccd1 _7939_/D sky130_fd_sc_hd__clkbuf_1
X_8511__210 vssd1 vssd1 vccd1 vccd1 _8511__210/HI caravel_irq[1] sky130_fd_sc_hd__conb_1
Xclkbuf_0__3440_ _7114_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3440_/X sky130_fd_sc_hd__clkbuf_16
X_8361_ _8361_/CLK _8361_/D vssd1 vssd1 vccd1 vccd1 _8361_/Q sky130_fd_sc_hd__dfxtp_1
X_4524_ _4524_/A vssd1 vssd1 vccd1 vccd1 _8179_/D sky130_fd_sc_hd__clkbuf_1
X_7312_ _6963_/A _7261_/B _7262_/A _7320_/B _7311_/Y vssd1 vssd1 vccd1 vccd1 _7321_/B
+ sky130_fd_sc_hd__o221ai_4
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8292_ _8292_/CLK _8292_/D vssd1 vssd1 vccd1 vccd1 _8292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4455_ _8207_/Q _4454_/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__mux2_1
X_7243_ _7478_/A _7241_/Y _7242_/X _7197_/X _7209_/X vssd1 vssd1 vccd1 vccd1 _7243_/X
+ sky130_fd_sc_hd__o2111a_1
X_4386_ _4515_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _4402_/S sky130_fd_sc_hd__or2_4
X_7174_ _8305_/Q vssd1 vssd1 vccd1 vccd1 _7184_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6125_ input35/X input2/X _6105_/B vssd1 vssd1 vccd1 vccd1 _6125_/X sky130_fd_sc_hd__o21a_4
XFILLER_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6056_/X sky130_fd_sc_hd__clkbuf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _8094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6997__487 _6999__489/A vssd1 vssd1 vccd1 vccd1 _8168_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5909_ _7677_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__or2_4
XFILLER_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267__201 _6268__202/A vssd1 vssd1 vccd1 vccd1 _7793_/CLK sky130_fd_sc_hd__inv_2
X_6902__415 _6902__415/A vssd1 vssd1 vccd1 vccd1 _8093_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7406__161 _7409__164/A vssd1 vssd1 vccd1 vccd1 _8372_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4240_ _4240_/A vssd1 vssd1 vccd1 vccd1 _8292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4171_ _8343_/Q _4014_/X _4175_/S vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ _7930_/CLK _7930_/D vssd1 vssd1 vccd1 vccd1 _7930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6842__384 _6843__385/A vssd1 vssd1 vccd1 vccd1 _8052_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _7861_/CLK _7861_/D vssd1 vssd1 vccd1 vccd1 _7861_/Q sky130_fd_sc_hd__dfxtp_1
X_6506__232 _6508__234/A vssd1 vssd1 vccd1 vccd1 _7872_/CLK sky130_fd_sc_hd__inv_2
X_6812_ _7683_/A _7498_/B _7494_/B _7689_/A vssd1 vssd1 vccd1 vccd1 _6813_/D sky130_fd_sc_hd__o2bb2a_1
X_7792_ _7792_/CLK _7792_/D vssd1 vssd1 vccd1 vccd1 _7792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3955_ _3955_/A vssd1 vssd1 vccd1 vccd1 _8412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6743_ _8430_/Q _7457_/A _6742_/X vssd1 vssd1 vccd1 vccd1 _7557_/A sky130_fd_sc_hd__a21oi_2
X_5625_ _7917_/Q _4981_/X _5629_/S vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__mux2_1
X_3886_ _8444_/Q vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__clkbuf_2
X_8413_ _8430_/CLK _8413_/D vssd1 vssd1 vccd1 vccd1 _8413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5556_ _5556_/A vssd1 vssd1 vccd1 vccd1 _7944_/D sky130_fd_sc_hd__clkbuf_1
X_8344_ _8344_/CLK _8344_/D vssd1 vssd1 vccd1 vccd1 _8344_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3423_ _7032_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3423_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8275_ _8275_/CLK _8275_/D vssd1 vssd1 vccd1 vccd1 _8275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5487_ _5487_/A vssd1 vssd1 vccd1 vccd1 _7999_/D sky130_fd_sc_hd__clkbuf_1
X_4507_ _8186_/Q _4238_/X _4507_/S vssd1 vssd1 vccd1 vccd1 _4508_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4438_ _4438_/A vssd1 vssd1 vccd1 vccd1 _8213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3285_ _6720_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3285_/X sky130_fd_sc_hd__clkbuf_16
X_7226_ _7311_/B _7262_/A _7343_/B _7320_/C vssd1 vssd1 vccd1 vccd1 _7228_/B sky130_fd_sc_hd__a211o_1
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ _4384_/S vssd1 vssd1 vccd1 vccd1 _4378_/S sky130_fd_sc_hd__buf_2
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7157_ _7153_/A _7305_/B _6395_/A vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__a21bo_1
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6108_/X sky130_fd_sc_hd__and2_1
X_6039_ _7814_/Q input31/X _6039_/S vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7130__94 _7131__95/A vssd1 vssd1 vccd1 vccd1 _8275_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3240_ clkbuf_0__3240_/X vssd1 vssd1 vccd1 vccd1 _6603__310/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5410_ _5373_/X _8036_/Q _5410_/S vssd1 vssd1 vccd1 vccd1 _5411_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6390_ _7683_/A _6390_/B _7672_/A vssd1 vssd1 vccd1 vccd1 _6390_/X sky130_fd_sc_hd__and3_1
Xoutput115 _5979_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
X_5341_ _5235_/S _5331_/X _5340_/Y vssd1 vssd1 vccd1 vccd1 _8068_/D sky130_fd_sc_hd__a21oi_1
Xoutput126 _6003_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput137 _5866_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
Xoutput159 _5940_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput148 _5918_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
X_8060_ _8060_/CLK _8060_/D vssd1 vssd1 vccd1 vccd1 _8060_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5272_ _7985_/Q _8020_/Q _5291_/S vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4223_ _8067_/Q vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__buf_2
X_4154_ _8350_/Q _4153_/X _4157_/S vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4085_ _8364_/Q _3992_/X _4093_/S vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__mux2_1
X_7913_ _7913_/CLK _7913_/D vssd1 vssd1 vccd1 vccd1 _7913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7844_ _8481_/CLK _7844_/D vssd1 vssd1 vccd1 vccd1 _7844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7775_ _8439_/CLK _7775_/D vssd1 vssd1 vccd1 vccd1 _7775_/Q sky130_fd_sc_hd__dfxtp_1
X_4987_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__buf_2
X_6726_ _6726_/A vssd1 vssd1 vccd1 vccd1 _6726_/X sky130_fd_sc_hd__buf_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3938_ _3937_/X _8452_/Q _3944_/S vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3438_ clkbuf_0__3438_/X vssd1 vssd1 vccd1 vccd1 _7132_/A sky130_fd_sc_hd__clkbuf_4
X_3869_ _5779_/A vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__clkbuf_4
X_6657_ _6657_/A vssd1 vssd1 vccd1 vccd1 _7974_/D sky130_fd_sc_hd__clkbuf_1
X_5608_ _5608_/A vssd1 vssd1 vccd1 vccd1 _7925_/D sky130_fd_sc_hd__clkbuf_1
X_5539_ _5539_/A _5815_/B vssd1 vssd1 vccd1 vccd1 _5555_/S sky130_fd_sc_hd__nor2_2
X_7066__543 _7068__545/A vssd1 vssd1 vccd1 vccd1 _8224_/CLK sky130_fd_sc_hd__inv_2
X_8327_ _8327_/CLK _8327_/D vssd1 vssd1 vccd1 vccd1 _8327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3406_ _6948_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3406_/X sky130_fd_sc_hd__clkbuf_16
X_8258_ _8258_/CLK _8258_/D vssd1 vssd1 vccd1 vccd1 _8258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8189_ _8189_/CLK _8189_/D vssd1 vssd1 vccd1 vccd1 _8189_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_15_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8418_/CLK sky130_fd_sc_hd__clkbuf_16
X_7209_ _7202_/X _7203_/Y _7206_/Y _7207_/Y _7208_/X vssd1 vssd1 vccd1 vccd1 _7209_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__buf_4
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7103__72 _7104__73/A vssd1 vssd1 vccd1 vccd1 _8253_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5890_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__clkbuf_1
X_4910_ _5777_/S vssd1 vssd1 vccd1 vccd1 _5769_/S sky130_fd_sc_hd__buf_4
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _6852_/B vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4772_ _7779_/Q _4765_/X _4768_/X _4771_/X vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__o211a_1
X_7560_ _7560_/A vssd1 vssd1 vccd1 vccd1 _8430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7491_ _7508_/A _8413_/Q vssd1 vssd1 vccd1 vccd1 _7491_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3223_ clkbuf_0__3223_/X vssd1 vssd1 vccd1 vccd1 _6521__245/A sky130_fd_sc_hd__clkbuf_4
X_6442_ _7839_/Q _5967_/A _6444_/S vssd1 vssd1 vccd1 vccd1 _6443_/A sky130_fd_sc_hd__mux2_1
X_8112_ _8112_/CLK _8112_/D vssd1 vssd1 vccd1 vccd1 _8112_/Q sky130_fd_sc_hd__dfxtp_1
X_6373_ _6412_/B vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5324_ _5087_/A _5328_/A _7649_/B _3949_/A vssd1 vssd1 vccd1 vccd1 _5326_/B sky130_fd_sc_hd__a31o_1
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8043_ _8043_/CLK _8043_/D vssd1 vssd1 vccd1 vccd1 _8043_/Q sky130_fd_sc_hd__dfxtp_1
X_5255_ _8406_/Q _8144_/Q _5269_/S vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4206_ _4221_/S vssd1 vssd1 vccd1 vccd1 _4215_/S sky130_fd_sc_hd__buf_2
X_5186_ _5184_/X _5185_/X _5186_/S vssd1 vssd1 vccd1 vccd1 _5187_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4137_/A vssd1 vssd1 vccd1 vccd1 _8356_/D sky130_fd_sc_hd__clkbuf_1
X_4068_ _4068_/A vssd1 vssd1 vccd1 vccd1 _8372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7827_ _8483_/CLK _7827_/D vssd1 vssd1 vccd1 vccd1 _7827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7385__145 _7385__145/A vssd1 vssd1 vccd1 vccd1 _8356_/CLK sky130_fd_sc_hd__inv_2
X_7758_ _8441_/CLK _7758_/D vssd1 vssd1 vccd1 vccd1 _7758_/Q sky130_fd_sc_hd__dfxtp_1
X_7689_ _7689_/A _7692_/B vssd1 vssd1 vccd1 vccd1 _7689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7619__29 _7619__29/A vssd1 vssd1 vccd1 vccd1 _8452_/CLK sky130_fd_sc_hd__inv_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5291_/S sky130_fd_sc_hd__buf_4
X_7088__60 _7088__60/A vssd1 vssd1 vccd1 vccd1 _8241_/CLK sky130_fd_sc_hd__inv_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7258__112 _7259__113/A vssd1 vssd1 vccd1 vccd1 _8295_/CLK sky130_fd_sc_hd__inv_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5942_ _5942_/A vssd1 vssd1 vccd1 vccd1 _5942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5873_ _5873_/A vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__clkbuf_1
X_4824_ _8193_/Q _4765_/X _4661_/A _4823_/X vssd1 vssd1 vccd1 vccd1 _4824_/X sky130_fd_sc_hd__o211a_1
X_7428__4 _7429__5/A vssd1 vssd1 vccd1 vccd1 _8390_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7612_ _7612_/A vssd1 vssd1 vccd1 vccd1 _8447_/D sky130_fd_sc_hd__clkbuf_1
X_4755_ _4755_/A _4803_/A vssd1 vssd1 vccd1 vccd1 _4793_/A sky130_fd_sc_hd__nand2_1
X_7543_ _7546_/A _7543_/B vssd1 vssd1 vccd1 vccd1 _8424_/D sky130_fd_sc_hd__nor2_1
X_4686_ _4637_/X _4685_/X _4644_/X vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__a21o_1
X_7474_ _8497_/Q _7474_/B vssd1 vssd1 vccd1 vccd1 _7477_/A sky130_fd_sc_hd__xor2_1
X_6425_ _7831_/Q _5949_/A _6433_/S vssd1 vssd1 vccd1 vccd1 _6426_/A sky130_fd_sc_hd__mux2_1
X_6356_ _6792_/A _6293_/X _6371_/A _6354_/X _6355_/X vssd1 vssd1 vccd1 vccd1 _6356_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5307_ _8199_/Q _8207_/Q _5307_/S vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8026_ _8026_/CLK _8026_/D vssd1 vssd1 vccd1 vccd1 _8026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6287_ _6287_/A vssd1 vssd1 vccd1 vccd1 _7654_/B sky130_fd_sc_hd__buf_2
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5238_ _7786_/Q _8383_/Q _5261_/S vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__mux2_1
X_5169_ _8202_/Q _8210_/Q _5294_/S vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3422_ clkbuf_0__3422_/X vssd1 vssd1 vccd1 vccd1 _7029__513/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7400__156 _7401__157/A vssd1 vssd1 vccd1 vccd1 _8367_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6500__227 _6500__227/A vssd1 vssd1 vccd1 vccd1 _7867_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4540_/A vssd1 vssd1 vccd1 vccd1 _8172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4471_ _4362_/X _8200_/Q _4473_/S vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6210_ _6210_/A vssd1 vssd1 vccd1 vccd1 _7765_/D sky130_fd_sc_hd__clkbuf_1
X_7190_ _7211_/A _7211_/B _7193_/B _8303_/Q vssd1 vssd1 vccd1 vccd1 _7191_/B sky130_fd_sc_hd__a31o_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_19 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5023_ _8088_/Q vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__inv_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3755_ clkbuf_0__3755_/X vssd1 vssd1 vccd1 vccd1 _7624__33/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5856_ _5856_/A _6129_/C vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__or2_4
X_4807_ _8047_/Q _4765_/A _4659_/A _4806_/X vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__o211a_1
X_5787_ _7796_/Q _4353_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5788_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _8195_/Q _7996_/Q _7932_/Q _7892_/Q _4669_/X _4670_/X vssd1 vssd1 vccd1 vccd1
+ _4738_/X sky130_fd_sc_hd__mux4_1
X_7526_ _7534_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _8417_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6555__272 _6558__275/A vssd1 vssd1 vccd1 vccd1 _7912_/CLK sky130_fd_sc_hd__inv_2
X_4669_ _8122_/Q vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__buf_2
X_7457_ _7457_/A _7457_/B vssd1 vssd1 vccd1 vccd1 _7458_/B sky130_fd_sc_hd__nand2_1
X_6408_ _8481_/Q _6408_/B _6410_/C vssd1 vssd1 vccd1 vccd1 _6408_/X sky130_fd_sc_hd__and3_1
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6928__435 _6928__435/A vssd1 vssd1 vccd1 vccd1 _8113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6339_ _8137_/Q _6318_/A _6319_/X vssd1 vssd1 vccd1 vccd1 _6339_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8009_ _8009_/CLK _8009_/D vssd1 vssd1 vccd1 vccd1 _8009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3405_ clkbuf_0__3405_/X vssd1 vssd1 vccd1 vccd1 _6947__450/A sky130_fd_sc_hd__clkbuf_4
X_7082__55 _7082__55/A vssd1 vssd1 vccd1 vccd1 _8236_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3420_ clkbuf_0__3420_/X vssd1 vssd1 vccd1 vccd1 _7015__501/A sky130_fd_sc_hd__clkbuf_16
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7398__155 _7398__155/A vssd1 vssd1 vccd1 vccd1 _8366_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_101 _3934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3971_ _8076_/Q vssd1 vssd1 vccd1 vccd1 _4287_/B sky130_fd_sc_hd__clkbuf_2
X_5710_ _5725_/S vssd1 vssd1 vccd1 vccd1 _5719_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6875__397 _6876__398/A vssd1 vssd1 vccd1 vccd1 _8073_/CLK sky130_fd_sc_hd__inv_2
X_5641_ _5562_/X _7910_/Q _5647_/S vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5572_ _5571_/X _7939_/Q _5572_/S vssd1 vssd1 vccd1 vccd1 _5573_/A sky130_fd_sc_hd__mux2_1
X_8360_ _8360_/CLK _8360_/D vssd1 vssd1 vccd1 vccd1 _8360_/Q sky130_fd_sc_hd__dfxtp_1
X_4523_ _4353_/X _8179_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__mux2_1
X_8291_ _8291_/CLK _8291_/D vssd1 vssd1 vccd1 vccd1 _8291_/Q sky130_fd_sc_hd__dfxtp_1
X_7311_ _8287_/Q _7311_/B vssd1 vssd1 vccd1 vccd1 _7311_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7242_ _7191_/A _7191_/B _7471_/A vssd1 vssd1 vccd1 vccd1 _7242_/X sky130_fd_sc_hd__a21o_1
X_4454_ _8442_/Q vssd1 vssd1 vccd1 vccd1 _4454_/X sky130_fd_sc_hd__clkbuf_4
X_4385_ _4385_/A vssd1 vssd1 vccd1 vccd1 _8231_/D sky130_fd_sc_hd__clkbuf_1
X_7173_ _7173_/A vssd1 vssd1 vccd1 vccd1 _7193_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6124_ _7764_/Q _6025_/B _6112_/A _6123_/X _6037_/A vssd1 vssd1 vccd1 vccd1 _6124_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7060__538 _7062__540/A vssd1 vssd1 vccd1 vccd1 _8219_/CLK sky130_fd_sc_hd__inv_2
X_6055_ _7743_/Q _6063_/B vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__or2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4413_/X _8094_/Q _5010_/S vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5908_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5917_/B sky130_fd_sc_hd__clkbuf_2
X_5839_ _4141_/X _7730_/Q _5843_/S vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__mux2_1
X_7509_ _7557_/B vssd1 vssd1 vccd1 vccd1 _7510_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8489_ _8489_/CLK _8489_/D vssd1 vssd1 vccd1 vccd1 _8489_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8534__233 vssd1 vssd1 vccd1 vccd1 _8534__233/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4170_/A vssd1 vssd1 vccd1 vccd1 _8344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _7860_/CLK _7860_/D vssd1 vssd1 vccd1 vccd1 _7860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6811_ _7689_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _6813_/C sky130_fd_sc_hd__nand2_1
X_7791_ _7791_/CLK _7791_/D vssd1 vssd1 vccd1 vccd1 _7791_/Q sky130_fd_sc_hd__dfxtp_1
X_3954_ _8412_/Q _3812_/X _3962_/S vssd1 vssd1 vccd1 vccd1 _3955_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6742_ _8430_/Q _8429_/Q _8428_/Q _6745_/B vssd1 vssd1 vccd1 vccd1 _6742_/X sky130_fd_sc_hd__and4b_1
X_3885_ _3885_/A vssd1 vssd1 vccd1 vccd1 _8469_/D sky130_fd_sc_hd__clkbuf_1
X_8412_ _8412_/CLK _8412_/D vssd1 vssd1 vccd1 vccd1 _8412_/Q sky130_fd_sc_hd__dfxtp_1
X_5624_ _5624_/A vssd1 vssd1 vccd1 vccd1 _7918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3422_ _7026_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3422_/X sky130_fd_sc_hd__clkbuf_16
X_8343_ _8343_/CLK _8343_/D vssd1 vssd1 vccd1 vccd1 _8343_/Q sky130_fd_sc_hd__dfxtp_1
X_5555_ _7944_/Q _4996_/X _5555_/S vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__mux2_1
X_8274_ _8274_/CLK _8274_/D vssd1 vssd1 vccd1 vccd1 _8274_/Q sky130_fd_sc_hd__dfxtp_1
X_5486_ _5343_/X _7999_/Q _5494_/S vssd1 vssd1 vccd1 vccd1 _5487_/A sky130_fd_sc_hd__mux2_1
X_4506_ _4506_/A vssd1 vssd1 vccd1 vccd1 _8187_/D sky130_fd_sc_hd__clkbuf_1
X_4437_ _8213_/Q _4436_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__mux2_1
X_7225_ _7323_/A _7325_/A vssd1 vssd1 vccd1 vccd1 _7343_/B sky130_fd_sc_hd__nor2_2
XFILLER_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7156_ _8310_/Q _7158_/B _8311_/Q vssd1 vssd1 vccd1 vccd1 _7305_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4368_ _4457_/A _5412_/A vssd1 vssd1 vccd1 vccd1 _4384_/S sky130_fd_sc_hd__or2_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6107_/A vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4299_ _4299_/A vssd1 vssd1 vccd1 vccd1 _8266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6038_ _6034_/X _6035_/X _6036_/X _6037_/X vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__o211a_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ _7989_/CLK _7989_/D vssd1 vssd1 vccd1 vccd1 _7989_/Q sky130_fd_sc_hd__dfxtp_1
X_8518__217 vssd1 vssd1 vccd1 vccd1 _8518__217/HI core0Index[4] sky130_fd_sc_hd__conb_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6262__198 _6263__199/A vssd1 vssd1 vccd1 vccd1 _7790_/CLK sky130_fd_sc_hd__inv_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7115__81 _7119__85/A vssd1 vssd1 vccd1 vccd1 _8262_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6568__282 _6569__283/A vssd1 vssd1 vccd1 vccd1 _7922_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7252__107 _7252__107/A vssd1 vssd1 vccd1 vccd1 _8290_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput116 _5981_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _5235_/S _5331_/A _7598_/A vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__o21ai_1
Xoutput127 _6005_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput149 _5879_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput138 _5877_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
X_5271_ _5220_/X _5269_/X _5270_/X vssd1 vssd1 vccd1 vccd1 _5271_/Y sky130_fd_sc_hd__o21ai_1
X_4222_ _4222_/A vssd1 vssd1 vccd1 vccd1 _8325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6135__176 _6138__179/A vssd1 vssd1 vccd1 vccd1 _7725_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4153_ _8061_/Q vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__buf_2
XFILLER_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _4099_/S vssd1 vssd1 vccd1 vccd1 _4093_/S sky130_fd_sc_hd__buf_2
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7912_ _7912_/CLK _7912_/D vssd1 vssd1 vccd1 vccd1 _7912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7843_ _8447_/CLK _7843_/D vssd1 vssd1 vccd1 vccd1 _7843_/Q sky130_fd_sc_hd__dfxtp_1
X_4986_ _4986_/A vssd1 vssd1 vccd1 vccd1 _8101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7774_ _8308_/CLK _7774_/D vssd1 vssd1 vccd1 vccd1 _7774_/Q sky130_fd_sc_hd__dfxtp_1
X_3937_ _8444_/Q vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3437_ clkbuf_0__3437_/X vssd1 vssd1 vccd1 vccd1 _7104__73/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6656_ _7974_/Q _5941_/A _6658_/S vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__mux2_1
X_3868_ _3949_/A _5329_/A _3948_/A vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__or3b_4
X_5607_ _5565_/X _7925_/Q _5611_/S vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__mux2_1
X_5538_ _5538_/A _5538_/B _4475_/B vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__or3b_2
X_8326_ _8326_/CLK _8326_/D vssd1 vssd1 vccd1 vccd1 _8326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3405_ _6942_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3405_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8257_ _8257_/CLK _8257_/D vssd1 vssd1 vccd1 vccd1 _8257_/Q sky130_fd_sc_hd__dfxtp_2
X_5469_ _5469_/A vssd1 vssd1 vccd1 vccd1 _8007_/D sky130_fd_sc_hd__clkbuf_1
X_7208_ _8499_/Q _7208_/B vssd1 vssd1 vccd1 vccd1 _7208_/X sky130_fd_sc_hd__or2_1
X_8188_ _8188_/CLK _8188_/D vssd1 vssd1 vccd1 vccd1 _8188_/Q sky130_fd_sc_hd__dfxtp_1
X_7139_ _7355_/A vssd1 vssd1 vccd1 vccd1 _7139_/X sky130_fd_sc_hd__buf_1
XFILLER_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _6103_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _4613_/A _8135_/Q _4925_/A _4839_/X _4678_/A vssd1 vssd1 vccd1 vccd1 _4840_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ _4769_/X _7907_/Q _7899_/Q _4770_/X _4757_/A vssd1 vssd1 vccd1 vccd1 _4771_/X
+ sky130_fd_sc_hd__a221o_1
X_6510_ _6510_/A vssd1 vssd1 vccd1 vccd1 _6510_/X sky130_fd_sc_hd__buf_1
XFILLER_119_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7490_ _7490_/A _7504_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7490_/Y sky130_fd_sc_hd__nor3b_1
Xclkbuf_1_1_0__3222_ clkbuf_0__3222_/X vssd1 vssd1 vccd1 vccd1 _6515__240/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6441_ _6441_/A vssd1 vssd1 vccd1 vccd1 _7838_/D sky130_fd_sc_hd__clkbuf_1
X_6372_ _6415_/B vssd1 vssd1 vccd1 vccd1 _6412_/B sky130_fd_sc_hd__clkbuf_2
X_8111_ _8111_/CLK _8111_/D vssd1 vssd1 vccd1 vccd1 _8111_/Q sky130_fd_sc_hd__dfxtp_1
X_5323_ _5323_/A vssd1 vssd1 vccd1 vccd1 _8075_/D sky130_fd_sc_hd__clkbuf_1
X_8042_ _8042_/CLK _8042_/D vssd1 vssd1 vccd1 vccd1 _8042_/Q sky130_fd_sc_hd__dfxtp_1
X_5254_ _5338_/B _5252_/X _5253_/X vssd1 vssd1 vccd1 vccd1 _5254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185_ _8258_/Q _8250_/Q _8242_/Q _8266_/Q _5078_/X _5070_/X vssd1 vssd1 vccd1 vccd1
+ _5185_/X sky130_fd_sc_hd__mux4_1
X_4205_ _5709_/A _5815_/A vssd1 vssd1 vccd1 vccd1 _4221_/S sky130_fd_sc_hd__nor2_2
XFILLER_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4136_ _8356_/Q _4101_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4137_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7419__172 _7419__172/A vssd1 vssd1 vccd1 vccd1 _8383_/CLK sky130_fd_sc_hd__inv_2
X_4067_ _3916_/X _8372_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _8483_/CLK _7826_/D vssd1 vssd1 vccd1 vccd1 _7826_/Q sky130_fd_sc_hd__dfxtp_1
X_4969_ _8106_/Q _4244_/X _4971_/S vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__mux2_1
X_7757_ _8441_/CLK _7757_/D vssd1 vssd1 vccd1 vccd1 _7757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6708_ _6726_/A vssd1 vssd1 vccd1 vccd1 _6708_/X sky130_fd_sc_hd__buf_1
X_7688_ _7688_/A vssd1 vssd1 vccd1 vccd1 _8487_/D sky130_fd_sc_hd__clkbuf_1
X_6519__243 _6521__245/A vssd1 vssd1 vccd1 vccd1 _7883_/CLK sky130_fd_sc_hd__inv_2
X_6639_ _6639_/A vssd1 vssd1 vccd1 vccd1 _7966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8309_ _8309_/CLK _8309_/D vssd1 vssd1 vccd1 vccd1 _8309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6728__362 _6728__362/A vssd1 vssd1 vccd1 vccd1 _8029_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _5941_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__or2_1
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _6642_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__and2_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8315_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4823_ _7890_/Q _4767_/X _4822_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7611_ _7611_/A _7615_/B _7613_/C vssd1 vssd1 vccd1 vccd1 _7612_/A sky130_fd_sc_hd__and3_1
X_4754_ _8123_/Q _8122_/Q vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__or2_2
X_7542_ _7462_/B _7527_/X _7517_/B _6800_/Y vssd1 vssd1 vccd1 vccd1 _7543_/B sky130_fd_sc_hd__o22a_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7473_ _8416_/Q _7473_/B vssd1 vssd1 vccd1 vccd1 _7474_/B sky130_fd_sc_hd__xor2_2
X_4685_ _8095_/Q _7982_/Q _7886_/Q _7862_/Q _4650_/X _4651_/X vssd1 vssd1 vccd1 vccd1
+ _4685_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6424_ _6468_/A vssd1 vssd1 vccd1 vccd1 _6433_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6355_ _6355_/A _6355_/B vssd1 vssd1 vccd1 vccd1 _6355_/X sky130_fd_sc_hd__and2_1
X_5306_ _8175_/Q _5178_/X _5285_/B _8167_/Q _5098_/A vssd1 vssd1 vccd1 vccd1 _5306_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6286_ _6401_/A vssd1 vssd1 vccd1 vccd1 _6286_/X sky130_fd_sc_hd__clkbuf_2
X_7024__509 _7024__509/A vssd1 vssd1 vccd1 vccd1 _8190_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8025_ _8025_/CLK _8025_/D vssd1 vssd1 vccd1 vccd1 _8025_/Q sky130_fd_sc_hd__dfxtp_1
X_5237_ _5338_/B _5235_/X _5236_/X vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _5305_/A vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__buf_2
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5099_ _5186_/S vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__clkbuf_2
X_7391__150 _7391__150/A vssd1 vssd1 vccd1 vccd1 _8361_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4119_ _4119_/A vssd1 vssd1 vccd1 vccd1 _4911_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7809_ _8497_/CLK _7809_/D vssd1 vssd1 vccd1 vccd1 _7809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2998_ clkbuf_0__2998_/X vssd1 vssd1 vccd1 vccd1 _6246__185/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7624__33 _7624__33/A vssd1 vssd1 vccd1 vccd1 _8456_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3619_ clkbuf_0__3619_/X vssd1 vssd1 vccd1 vccd1 _7398__155/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _4470_/A vssd1 vssd1 vccd1 vccd1 _8201_/D sky130_fd_sc_hd__clkbuf_1
X_6140_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6140_/X sky130_fd_sc_hd__buf_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _6053_/X _6069_/X _6070_/X _6056_/X vssd1 vssd1 vccd1 vccd1 _6071_/X sky130_fd_sc_hd__o211a_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6661__313 _6663__315/A vssd1 vssd1 vccd1 vccd1 _7977_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5924_ _5924_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__or2_4
XFILLER_110_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5855_ _6000_/A _5854_/X _7724_/Q vssd1 vssd1 vccd1 vccd1 _6129_/C sky130_fd_sc_hd__a21o_2
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _8108_/Q _4767_/A _4805_/X _4776_/A vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5786_ _5786_/A vssd1 vssd1 vccd1 vccd1 _7797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4737_ _4715_/X _4736_/X _4665_/A vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__a21o_1
X_7525_ _7476_/B _7476_/C _7516_/X _7522_/X _6782_/B vssd1 vssd1 vccd1 vccd1 _7526_/B
+ sky130_fd_sc_hd__a32oi_1
X_6887__406 _6887__406/A vssd1 vssd1 vccd1 vccd1 _8082_/CLK sky130_fd_sc_hd__inv_2
X_4668_ _8104_/Q _8059_/Q _7943_/Q _8296_/Q _4648_/A _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4668_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6967__463 _6968__464/A vssd1 vssd1 vccd1 vccd1 _8144_/CLK sky130_fd_sc_hd__inv_2
X_6407_ _7825_/Q _6401_/X _6393_/X _6406_/X _6391_/X vssd1 vssd1 vccd1 vccd1 _7825_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4599_ _4599_/A vssd1 vssd1 vccd1 vccd1 _8146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6338_ _7197_/A _6293_/A _6299_/X vssd1 vssd1 vccd1 vccd1 _6338_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8008_ _8008_/CLK _8008_/D vssd1 vssd1 vccd1 vccd1 _8008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3404_ clkbuf_0__3404_/X vssd1 vssd1 vccd1 vccd1 _6941__445/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6562__277 _6563__278/A vssd1 vssd1 vccd1 vccd1 _7917_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3281_ clkbuf_0__3281_/X vssd1 vssd1 vccd1 vccd1 _6719__355/A sky130_fd_sc_hd__clkbuf_16
XFILLER_25_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_102 _6037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3970_ _5412_/A vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__buf_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _5640_/A vssd1 vssd1 vccd1 vccd1 _7911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5571_ _5571_/A vssd1 vssd1 vccd1 vccd1 _5571_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4522_ _4522_/A vssd1 vssd1 vccd1 vccd1 _8180_/D sky130_fd_sc_hd__clkbuf_1
X_8290_ _8290_/CLK _8290_/D vssd1 vssd1 vccd1 vccd1 _8290_/Q sky130_fd_sc_hd__dfxtp_1
X_7310_ _7317_/B vssd1 vssd1 vccd1 vccd1 _7315_/A sky130_fd_sc_hd__inv_2
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4453_ _4453_/A vssd1 vssd1 vccd1 vccd1 _8208_/D sky130_fd_sc_hd__clkbuf_1
X_7241_ _7241_/A _7241_/B vssd1 vssd1 vccd1 vccd1 _7241_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ _4365_/X _8231_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__mux2_1
X_7172_ _7468_/A _7172_/B vssd1 vssd1 vccd1 vccd1 _7183_/A sky130_fd_sc_hd__xnor2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6123_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__and2_1
XFILLER_100_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6054_ _7818_/Q input4/X _6058_/S vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__mux2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _8095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5907_ _5907_/A vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5838_ _5838_/A vssd1 vssd1 vccd1 vccd1 _7731_/D sky130_fd_sc_hd__clkbuf_1
X_6934__440 _6934__440/A vssd1 vssd1 vccd1 vccd1 _8118_/CLK sky130_fd_sc_hd__inv_2
X_5769_ _4144_/X _7804_/Q _5769_/S vssd1 vssd1 vccd1 vccd1 _5770_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7508_ _7508_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7557_/B sky130_fd_sc_hd__and2_2
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8488_ _8489_/CLK _8488_/D vssd1 vssd1 vccd1 vccd1 _8488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6668__319 _6669__320/A vssd1 vssd1 vccd1 vccd1 _7983_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6274__207 _6275__208/A vssd1 vssd1 vccd1 vccd1 _7799_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6810_ _6810_/A _6810_/B vssd1 vssd1 vccd1 vccd1 _7494_/B sky130_fd_sc_hd__nand2_2
XFILLER_36_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7413__167 _7414__168/A vssd1 vssd1 vccd1 vccd1 _8378_/CLK sky130_fd_sc_hd__inv_2
X_7790_ _7790_/CLK _7790_/D vssd1 vssd1 vccd1 vccd1 _7790_/Q sky130_fd_sc_hd__dfxtp_1
X_3953_ _3968_/S vssd1 vssd1 vccd1 vccd1 _3962_/S sky130_fd_sc_hd__buf_2
X_6741_ _8429_/Q _8428_/Q _6745_/B vssd1 vssd1 vccd1 vccd1 _7457_/A sky130_fd_sc_hd__nand3_2
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3884_ _8469_/Q _3883_/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8411_ _8411_/CLK _8411_/D vssd1 vssd1 vccd1 vccd1 _8411_/Q sky130_fd_sc_hd__dfxtp_1
X_5623_ _7918_/Q _4978_/X _5629_/S vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3421_ _7020_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3421_/X sky130_fd_sc_hd__clkbuf_16
X_8342_ _8342_/CLK _8342_/D vssd1 vssd1 vccd1 vccd1 _8342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _7945_/D sky130_fd_sc_hd__clkbuf_1
X_8273_ _8273_/CLK _8273_/D vssd1 vssd1 vccd1 vccd1 _8273_/Q sky130_fd_sc_hd__dfxtp_1
X_5485_ _5500_/S vssd1 vssd1 vccd1 vccd1 _5494_/S sky130_fd_sc_hd__clkbuf_4
X_4505_ _8187_/Q _4235_/X _4507_/S vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4436_ _8448_/Q vssd1 vssd1 vccd1 vccd1 _4436_/X sky130_fd_sc_hd__buf_2
X_7224_ _8482_/Q _7270_/A vssd1 vssd1 vccd1 vccd1 _7325_/A sky130_fd_sc_hd__nand2_1
X_6513__238 _6514__239/A vssd1 vssd1 vccd1 vccd1 _7878_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4367_ _4367_/A vssd1 vssd1 vccd1 vccd1 _8239_/D sky130_fd_sc_hd__clkbuf_1
X_7155_ _8484_/Q _7155_/B vssd1 vssd1 vccd1 vccd1 _7246_/B sky130_fd_sc_hd__xor2_1
XFILLER_116_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _7757_/Q _6095_/X _6099_/X _6105_/X _6093_/X vssd1 vssd1 vccd1 vccd1 _6106_/X
+ sky130_fd_sc_hd__o221a_1
X_4298_ _3934_/X _8266_/Q _4298_/S vssd1 vssd1 vccd1 vccd1 _4299_/A sky130_fd_sc_hd__mux2_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6037_ _6037_/A vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ _7988_/CLK _7988_/D vssd1 vssd1 vccd1 vccd1 _7988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2998_ _6140_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2998_/X sky130_fd_sc_hd__clkbuf_16
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3619_ _7393_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3619_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7141__102 _7141__102/A vssd1 vssd1 vccd1 vccd1 _8283_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6722__357 _6723__358/A vssd1 vssd1 vccd1 vccd1 _8024_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput128 _6007_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput139 _5899_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput117 _5983_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
X_5270_ _8398_/Q _5227_/X _5189_/X _8390_/Q _5152_/A vssd1 vssd1 vccd1 vccd1 _5270_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _8325_/Q _4156_/X _4221_/S vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4152_ _4152_/A vssd1 vssd1 vccd1 vccd1 _8351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4083_ _4083_/A _4178_/B vssd1 vssd1 vccd1 vccd1 _4099_/S sky130_fd_sc_hd__nor2_2
X_7911_ _7911_/CLK _7911_/D vssd1 vssd1 vccd1 vccd1 _7911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7842_ _8478_/CLK _7842_/D vssd1 vssd1 vccd1 vccd1 _7842_/Q sky130_fd_sc_hd__dfxtp_1
X_4985_ _8101_/Q _4984_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7773_ _8308_/CLK _7773_/D vssd1 vssd1 vccd1 vccd1 _7773_/Q sky130_fd_sc_hd__dfxtp_1
X_3936_ _3936_/A vssd1 vssd1 vccd1 vccd1 _8453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3436_ clkbuf_0__3436_/X vssd1 vssd1 vccd1 vccd1 _7100__70/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6655_ _6655_/A vssd1 vssd1 vccd1 vccd1 _7973_/D sky130_fd_sc_hd__clkbuf_1
X_3867_ _7607_/A _6473_/A _3866_/X _6206_/A vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__a31oi_4
X_5606_ _5606_/A vssd1 vssd1 vccd1 vccd1 _7926_/D sky130_fd_sc_hd__clkbuf_1
X_5537_ _5537_/A vssd1 vssd1 vccd1 vccd1 _7976_/D sky130_fd_sc_hd__clkbuf_1
X_8325_ _8325_/CLK _8325_/D vssd1 vssd1 vccd1 vccd1 _8325_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3404_ _6935_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3404_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8256_ _8256_/CLK _8256_/D vssd1 vssd1 vccd1 vccd1 _8256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _8007_/Q _4342_/A _5476_/S vssd1 vssd1 vccd1 vccd1 _5469_/A sky130_fd_sc_hd__mux2_1
X_7207_ _7207_/A _7208_/B vssd1 vssd1 vccd1 vccd1 _7207_/Y sky130_fd_sc_hd__nand2_1
X_5399_ _5399_/A vssd1 vssd1 vccd1 vccd1 _8042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4419_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _4419_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8187_ _8187_/CLK _8187_/D vssd1 vssd1 vccd1 vccd1 _8187_/Q sky130_fd_sc_hd__dfxtp_1
X_7138_ _7392_/A vssd1 vssd1 vccd1 vccd1 _7138_/X sky130_fd_sc_hd__buf_1
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7069_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7069_/X sky130_fd_sc_hd__buf_1
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7073__549 _7073__549/A vssd1 vssd1 vccd1 vccd1 _8230_/CLK sky130_fd_sc_hd__inv_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8498_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _6105_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6947__450 _6947__450/A vssd1 vssd1 vccd1 vccd1 _8129_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4770_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__3444_ clkbuf_0__3444_/X vssd1 vssd1 vccd1 vccd1 _7355_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3221_ clkbuf_0__3221_/X vssd1 vssd1 vccd1 vccd1 _6509__235/A sky130_fd_sc_hd__clkbuf_4
X_6141__181 _6143__183/A vssd1 vssd1 vccd1 vccd1 _7730_/CLK sky130_fd_sc_hd__inv_2
X_6440_ _7838_/Q _5965_/A _6444_/S vssd1 vssd1 vccd1 vccd1 _6441_/A sky130_fd_sc_hd__mux2_1
X_6371_ _6371_/A vssd1 vssd1 vccd1 vccd1 _6371_/X sky130_fd_sc_hd__clkbuf_2
X_8110_ _8110_/CLK _8110_/D vssd1 vssd1 vccd1 vccd1 _8110_/Q sky130_fd_sc_hd__dfxtp_1
X_5322_ _7598_/A _5322_/B _5322_/C vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__and3_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8041_ _8041_/CLK _8041_/D vssd1 vssd1 vccd1 vccd1 _8041_/Q sky130_fd_sc_hd__dfxtp_1
X_5253_ _8232_/Q _5163_/X _5189_/X _8467_/Q _5160_/A vssd1 vssd1 vccd1 vccd1 _5253_/X
+ sky130_fd_sc_hd__o221a_1
X_5184_ _8376_/Q _8274_/Q _8011_/Q _8226_/Q _5064_/A _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5184_/X sky130_fd_sc_hd__mux4_1
X_4204_ _5601_/A vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4157_/S vssd1 vssd1 vccd1 vccd1 _4148_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4081_/S vssd1 vssd1 vccd1 vccd1 _4075_/S sky130_fd_sc_hd__buf_2
X_7825_ _8483_/CLK _7825_/D vssd1 vssd1 vccd1 vccd1 _7825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _4968_/A vssd1 vssd1 vccd1 vccd1 _8107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7756_ _8441_/CLK _7756_/D vssd1 vssd1 vccd1 vccd1 _7756_/Q sky130_fd_sc_hd__dfxtp_1
X_6707_ _6879_/A vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__buf_1
X_7687_ _7722_/A _7687_/B vssd1 vssd1 vccd1 vccd1 _7688_/A sky130_fd_sc_hd__or2_1
X_4899_ _4428_/X _4610_/A _4898_/X _4841_/X vssd1 vssd1 vccd1 vccd1 _8133_/D sky130_fd_sc_hd__o211a_1
X_3919_ _5087_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _4025_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__3419_ clkbuf_0__3419_/X vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__clkbuf_4
X_6638_ _5924_/A _7966_/Q _6640_/S vssd1 vssd1 vccd1 vccd1 _6639_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8308_ _8308_/CLK _8308_/D vssd1 vssd1 vccd1 vccd1 _8308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8239_ _8239_/CLK _8239_/D vssd1 vssd1 vccd1 vccd1 _8239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5940_ _5940_/A vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5871_ _5871_/A vssd1 vssd1 vccd1 vccd1 _5871_/X sky130_fd_sc_hd__clkbuf_1
X_7610_ _7610_/A vssd1 vssd1 vccd1 vccd1 _8446_/D sky130_fd_sc_hd__clkbuf_1
X_4822_ _4801_/A _7994_/Q _7930_/Q _4787_/A vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4753_/A vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__clkbuf_2
X_7541_ _7546_/A _7541_/B vssd1 vssd1 vccd1 vccd1 _8423_/D sky130_fd_sc_hd__nor2_1
X_7472_ _7472_/A _7472_/B _7472_/C _7472_/D vssd1 vssd1 vccd1 vccd1 _7486_/B sky130_fd_sc_hd__or4_1
XFILLER_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4684_ _8050_/Q _8042_/Q _7870_/Q _8111_/Q _4630_/X _4633_/X vssd1 vssd1 vccd1 vccd1
+ _4684_/X sky130_fd_sc_hd__mux4_1
X_6423_ _6423_/A _7652_/A _7724_/D vssd1 vssd1 vccd1 vccd1 _6468_/A sky130_fd_sc_hd__and3_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ _8139_/Q _6318_/X _6353_/X vssd1 vssd1 vccd1 vccd1 _6354_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5305_ _5305_/A _5305_/B vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__or2_1
X_6285_ _6343_/A vssd1 vssd1 vccd1 vccd1 _6401_/A sky130_fd_sc_hd__buf_2
X_8024_ _8024_/CLK _8024_/D vssd1 vssd1 vccd1 vccd1 _8024_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5214_/X _8029_/Q _7794_/Q _5216_/X _5099_/X vssd1 vssd1 vccd1 vccd1 _5236_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5305_/A sky130_fd_sc_hd__clkbuf_2
X_7094__65 _7094__65/A vssd1 vssd1 vccd1 vccd1 _8246_/CLK sky130_fd_sc_hd__inv_2
X_5098_ _5098_/A vssd1 vssd1 vccd1 vccd1 _5186_/S sky130_fd_sc_hd__buf_2
X_4118_ _8130_/Q _4120_/B _4119_/A vssd1 vssd1 vccd1 vccd1 _4118_/X sky130_fd_sc_hd__o21a_1
X_4049_ _4049_/A vssd1 vssd1 vccd1 vccd1 _8380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7808_ _8499_/CLK _7808_/D vssd1 vssd1 vccd1 vccd1 _7808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7739_ _8490_/CLK _7739_/D vssd1 vssd1 vccd1 vccd1 _7739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2997_ clkbuf_0__2997_/X vssd1 vssd1 vccd1 vccd1 _6138__179/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3618_ clkbuf_0__3618_/X vssd1 vssd1 vccd1 vccd1 _7417_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3549_ clkbuf_0__3549_/X vssd1 vssd1 vccd1 vccd1 _7252__107/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6070_ _7747_/Q _6082_/B vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__or2_1
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5021_ _5087_/A _7323_/A vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__nand2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5923_ _5923_/A vssd1 vssd1 vccd1 vccd1 _5923_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ _7969_/Q _7970_/Q _7971_/Q vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__and3_1
X_4805_ _4780_/A _8039_/Q _7867_/Q _4781_/A vssd1 vssd1 vccd1 vccd1 _4805_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5785_ _7797_/Q _4350_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__mux2_1
X_7030__514 _7031__515/A vssd1 vssd1 vccd1 vccd1 _8195_/CLK sky130_fd_sc_hd__inv_2
X_7524_ _7534_/A _7524_/B vssd1 vssd1 vccd1 vccd1 _8416_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4736_ _7924_/Q _7804_/Q _7729_/Q _7916_/Q _4640_/A _4638_/X vssd1 vssd1 vccd1 vccd1
+ _4736_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7455_ _7633_/A vssd1 vssd1 vccd1 vccd1 _7455_/X sky130_fd_sc_hd__buf_1
X_4667_ _4670_/A vssd1 vssd1 vccd1 vccd1 _4667_/X sky130_fd_sc_hd__buf_2
X_7386_ _7386_/A vssd1 vssd1 vccd1 vccd1 _7386_/X sky130_fd_sc_hd__buf_1
X_6406_ _6963_/A _6408_/B _6410_/C vssd1 vssd1 vccd1 vccd1 _6406_/X sky130_fd_sc_hd__and3_1
X_4598_ _8146_/Q _4445_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__mux2_1
X_6337_ _8495_/Q vssd1 vssd1 vccd1 vccd1 _7197_/A sky130_fd_sc_hd__buf_4
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5219_ _8273_/Q _8010_/Q _5241_/S vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__mux2_1
X_8007_ _8007_/CLK _8007_/D vssd1 vssd1 vccd1 vccd1 _8007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6199_ _7969_/Q _6197_/X _6195_/X _6198_/X _7758_/Q vssd1 vssd1 vccd1 vccd1 _7758_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3403_ clkbuf_0__3403_/X vssd1 vssd1 vccd1 vccd1 _6932__438/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_103 _6037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5570_ _5570_/A vssd1 vssd1 vccd1 vccd1 _7940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ _4350_/X _8180_/Q _4525_/S vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4452_ _8208_/Q _4451_/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__mux2_1
X_7240_ _6792_/A _7192_/B _7200_/X _7239_/X vssd1 vssd1 vccd1 vccd1 _7240_/X sky130_fd_sc_hd__o211a_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4383_ _4383_/A vssd1 vssd1 vccd1 vccd1 _8232_/D sky130_fd_sc_hd__clkbuf_1
X_7171_ _7232_/B _7232_/C vssd1 vssd1 vccd1 vccd1 _7172_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6122_ _7763_/Q _6111_/X _6112_/X _6121_/X _6037_/A vssd1 vssd1 vccd1 vccd1 _6122_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6053_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__clkbuf_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _4410_/X _8095_/Q _5010_/S vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6976_/A vssd1 vssd1 vccd1 vccd1 _6955_/X sky130_fd_sc_hd__buf_1
X_5906_ _7681_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__or2_1
XFILLER_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6886_ _6886_/A vssd1 vssd1 vccd1 vccd1 _6886_/X sky130_fd_sc_hd__buf_1
X_5837_ _4138_/X _7731_/Q _5843_/S vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5768_ _5768_/A vssd1 vssd1 vccd1 vccd1 _7805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4719_ _8102_/Q _8057_/Q _7941_/Q _8294_/Q _4669_/X _4670_/X vssd1 vssd1 vccd1 vccd1
+ _4719_/X sky130_fd_sc_hd__mux4_1
X_7507_ _7544_/A _7506_/X _7508_/B vssd1 vssd1 vccd1 vccd1 _7511_/C sky130_fd_sc_hd__a21o_1
X_8487_ _8498_/CLK _8487_/D vssd1 vssd1 vccd1 vccd1 _8487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_108_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5699_ _7884_/Q _4984_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__mux2_1
X_7127__91 _7128__92/A vssd1 vssd1 vccd1 vccd1 _8272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6941__445 _6941__445/A vssd1 vssd1 vccd1 vccd1 _8124_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6740_ _8427_/Q _6808_/A _6789_/B _6749_/A vssd1 vssd1 vccd1 vccd1 _6745_/B sky130_fd_sc_hd__and4_1
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _4588_/A _5502_/B vssd1 vssd1 vccd1 vccd1 _3968_/S sky130_fd_sc_hd__nor2_2
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3883_ _8445_/Q vssd1 vssd1 vccd1 vccd1 _3883_/X sky130_fd_sc_hd__clkbuf_2
X_8410_ _8410_/CLK _8410_/D vssd1 vssd1 vccd1 vccd1 _8410_/Q sky130_fd_sc_hd__dfxtp_1
X_5622_ _5622_/A vssd1 vssd1 vccd1 vccd1 _7919_/D sky130_fd_sc_hd__clkbuf_1
X_5553_ _7945_/Q _4993_/X _5555_/S vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3420_ _7014_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3420_/X sky130_fd_sc_hd__clkbuf_16
X_8341_ _8341_/CLK _8341_/D vssd1 vssd1 vccd1 vccd1 _8341_/Q sky130_fd_sc_hd__dfxtp_1
X_4504_ _4504_/A vssd1 vssd1 vccd1 vccd1 _8188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5484_ _5655_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5500_/S sky130_fd_sc_hd__or2_2
X_8272_ _8272_/CLK _8272_/D vssd1 vssd1 vccd1 vccd1 _8272_/Q sky130_fd_sc_hd__dfxtp_1
X_4435_ _4435_/A vssd1 vssd1 vccd1 vccd1 _8214_/D sky130_fd_sc_hd__clkbuf_1
X_7223_ _7270_/B vssd1 vssd1 vccd1 vccd1 _7262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _4365_/X _8239_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__mux2_1
X_7154_ _8312_/Q _7305_/A vssd1 vssd1 vccd1 vccd1 _7155_/B sky130_fd_sc_hd__xor2_1
X_6105_ _6105_/A _6105_/B vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__and2_4
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4297_ _4297_/A vssd1 vssd1 vccd1 vccd1 _8267_/D sky130_fd_sc_hd__clkbuf_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6036_ _7738_/Q _6044_/B vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__or2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ _7987_/CLK _7987_/D vssd1 vssd1 vccd1 vccd1 _7987_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2997_ _6134_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2997_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _7649_/A _6938_/B vssd1 vssd1 vccd1 vccd1 _8121_/D sky130_fd_sc_hd__nor2_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6674__324 _6675__325/A vssd1 vssd1 vccd1 vccd1 _7988_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3618_ _7392_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3618_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3549_ _7250_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3549_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6280__212 _6282__214/A vssd1 vssd1 vccd1 vccd1 _7804_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6575__288 _6577__290/A vssd1 vssd1 vccd1 vccd1 _7928_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput118 _5986_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput129 _5950_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
XFILLER_114_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4220_ _4220_/A vssd1 vssd1 vccd1 vccd1 _8326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7121__86 _7123__88/A vssd1 vssd1 vccd1 vccd1 _8267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _8351_/Q _4150_/X _4157_/S vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__mux2_1
X_4082_ _4082_/A vssd1 vssd1 vccd1 vccd1 _8365_/D sky130_fd_sc_hd__clkbuf_1
X_7910_ _7910_/CLK _7910_/D vssd1 vssd1 vccd1 vccd1 _7910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7841_ _8446_/CLK _7841_/D vssd1 vssd1 vccd1 vccd1 _7841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4984_ _8064_/Q vssd1 vssd1 vccd1 vccd1 _4984_/X sky130_fd_sc_hd__buf_2
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7772_ _8490_/CLK _7772_/D vssd1 vssd1 vccd1 vccd1 _7772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _3934_/X _8453_/Q _3935_/S vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3435_ clkbuf_0__3435_/X vssd1 vssd1 vccd1 vccd1 _7094__65/A sky130_fd_sc_hd__clkbuf_4
X_6654_ _7973_/Q _5939_/A _6658_/S vssd1 vssd1 vccd1 vccd1 _6655_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5605_ _5562_/X _7926_/Q _5611_/S vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__mux2_1
X_3866_ _7659_/A _7659_/B _4108_/D vssd1 vssd1 vccd1 vccd1 _3866_/X sky130_fd_sc_hd__and3_1
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5536_ _5373_/X _7976_/Q _5536_/S vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3403_ _6929_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3403_/X sky130_fd_sc_hd__clkbuf_16
X_8324_ _8442_/CLK _8324_/D vssd1 vssd1 vccd1 vccd1 _8324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5482_/S vssd1 vssd1 vccd1 vccd1 _5476_/S sky130_fd_sc_hd__buf_2
X_8255_ _8255_/CLK _8255_/D vssd1 vssd1 vccd1 vccd1 _8255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7206_ _8498_/Q _7206_/B vssd1 vssd1 vccd1 vccd1 _7206_/Y sky130_fd_sc_hd__xnor2_1
X_4418_ _4418_/A vssd1 vssd1 vccd1 vccd1 _8219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5398_ _5349_/X _8042_/Q _5404_/S vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8186_ _8186_/CLK _8186_/D vssd1 vssd1 vccd1 vccd1 _8186_/Q sky130_fd_sc_hd__dfxtp_1
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _8245_/D sky130_fd_sc_hd__clkbuf_1
X_8524__223 vssd1 vssd1 vccd1 vccd1 _8524__223/HI core1Index[3] sky130_fd_sc_hd__conb_1
XFILLER_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6019_ _6009_/X _6011_/X _6014_/X _6018_/X vssd1 vssd1 vccd1 vccd1 _6019_/X sky130_fd_sc_hd__o211a_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7008__496 _7009__497/A vssd1 vssd1 vccd1 vccd1 _8177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6954__455 _6954__455/A vssd1 vssd1 vccd1 vccd1 _8134_/CLK sky130_fd_sc_hd__inv_2
X_6245__184 _6246__185/A vssd1 vssd1 vccd1 vccd1 _7776_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3220_ clkbuf_0__3220_/X vssd1 vssd1 vccd1 vccd1 _6503__230/A sky130_fd_sc_hd__clkbuf_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6370_ _6370_/A vssd1 vssd1 vccd1 vccd1 _7816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5321_ _5321_/A _5321_/B vssd1 vssd1 vccd1 vccd1 _5322_/C sky130_fd_sc_hd__or2_1
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8040_ _8040_/CLK _8040_/D vssd1 vssd1 vccd1 vccd1 _8040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5252_ _8200_/Q _8208_/Q _5269_/S vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5183_ _5336_/B _5173_/X _5181_/X _5334_/B vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__a211o_1
X_4203_ _4405_/B _4904_/A _4903_/B vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__or3b_4
X_4134_ _5709_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _4157_/S sky130_fd_sc_hd__nor2_2
XFILLER_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4515_/A _4178_/B vssd1 vssd1 vccd1 vccd1 _4081_/S sky130_fd_sc_hd__or2_2
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7824_ _8483_/CLK _7824_/D vssd1 vssd1 vccd1 vccd1 _7824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _8107_/Q _4241_/X _4971_/S vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7755_ _8418_/CLK _7755_/D vssd1 vssd1 vccd1 vccd1 _7755_/Q sky130_fd_sc_hd__dfxtp_1
X_7686_ _8487_/Q _7698_/B _7699_/B _5902_/A vssd1 vssd1 vccd1 vccd1 _7687_/B sky130_fd_sc_hd__a22o_1
XFILLER_22_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4898_ _4613_/A _8133_/Q _4925_/A _4897_/X _4678_/A vssd1 vssd1 vccd1 vccd1 _4898_/X
+ sky130_fd_sc_hd__a221o_1
X_3918_ _3918_/A vssd1 vssd1 vccd1 vccd1 _7649_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0__3418_ clkbuf_0__3418_/X vssd1 vssd1 vccd1 vccd1 _7012__500/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6637_ _6637_/A vssd1 vssd1 vccd1 vccd1 _7965_/D sky130_fd_sc_hd__clkbuf_1
X_3849_ _5853_/B vssd1 vssd1 vccd1 vccd1 _6473_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5519_ _5519_/A vssd1 vssd1 vccd1 vccd1 _7984_/D sky130_fd_sc_hd__clkbuf_1
X_8307_ _8308_/CLK _8307_/D vssd1 vssd1 vccd1 vccd1 _8307_/Q sky130_fd_sc_hd__dfxtp_1
X_8238_ _8238_/CLK _8238_/D vssd1 vssd1 vccd1 vccd1 _8238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7636__43 _7638__45/A vssd1 vssd1 vccd1 vccd1 _8466_/CLK sky130_fd_sc_hd__inv_2
X_8169_ _8169_/CLK _8169_/D vssd1 vssd1 vccd1 vccd1 _8169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6526__249 _6527__250/A vssd1 vssd1 vccd1 vccd1 _7889_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6687__334 _6688__335/A vssd1 vssd1 vccd1 vccd1 _7998_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5870_ _6624_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__and2_1
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4821_ _8291_/Q _4778_/X _8099_/Q _4762_/X _4696_/S vssd1 vssd1 vccd1 vccd1 _4821_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__clkbuf_2
X_7540_ _8423_/Q _7530_/X _7527_/X _7492_/B vssd1 vssd1 vccd1 vccd1 _7541_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7471_ _7471_/A _7471_/B _7471_/C vssd1 vssd1 vccd1 vccd1 _7472_/D sky130_fd_sc_hd__and3_1
X_4683_ _4404_/X _4610_/X _4679_/X _4682_/X vssd1 vssd1 vccd1 vccd1 _8140_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6422_ _6343_/X _6415_/X _6419_/X _7830_/Q _6421_/X vssd1 vssd1 vccd1 vccd1 _7830_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6353_ _6353_/A vssd1 vssd1 vccd1 vccd1 _6353_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5304_ _8405_/Q _8143_/Q _5307_/S vssd1 vssd1 vccd1 vccd1 _5305_/B sky130_fd_sc_hd__mux2_1
X_6284_ _6415_/B _6294_/A vssd1 vssd1 vccd1 vccd1 _6343_/A sky130_fd_sc_hd__and2b_1
X_8023_ _8023_/CLK _8023_/D vssd1 vssd1 vccd1 vccd1 _8023_/Q sky130_fd_sc_hd__dfxtp_1
X_7079__52 _7079__52/A vssd1 vssd1 vccd1 vccd1 _8233_/CLK sky130_fd_sc_hd__inv_2
X_5235_ _8281_/Q _8002_/Q _5235_/S vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__mux2_1
X_5166_ _5166_/A _5188_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5097_ _5038_/X _5093_/X _5096_/X vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4117_ _8129_/Q _8128_/Q _8127_/Q vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__and3_1
X_4048_ _8380_/Q _3992_/X _4056_/S vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7807_ _7807_/CLK _7807_/D vssd1 vssd1 vccd1 vccd1 _7807_/Q sky130_fd_sc_hd__dfxtp_1
X_5999_ _6061_/A vssd1 vssd1 vccd1 vccd1 _6105_/B sky130_fd_sc_hd__buf_8
XFILLER_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7738_ _8498_/CLK _7738_/D vssd1 vssd1 vccd1 vccd1 _7738_/Q sky130_fd_sc_hd__dfxtp_1
X_7669_ _6963_/A _7656_/X _7668_/X _7662_/X vssd1 vssd1 vccd1 vccd1 _8482_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2996_ clkbuf_0__2996_/X vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__clkbuf_4
X_6532__253 _6534__255/A vssd1 vssd1 vccd1 vccd1 _7893_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3617_ clkbuf_0__3617_/X vssd1 vssd1 vccd1 vccd1 _7389__148/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5020_ _6895_/C vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__clkinv_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7375__136 _7376__137/A vssd1 vssd1 vccd1 vccd1 _8347_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7630__38 _7632__40/A vssd1 vssd1 vccd1 vccd1 _8461_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _5922_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__or2_4
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5853_ _7968_/Q _5853_/B _5853_/C vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__and3_1
XFILLER_34_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5784_ _5784_/A vssd1 vssd1 vccd1 vccd1 _7798_/D sky130_fd_sc_hd__clkbuf_1
X_4804_ _4778_/X _7859_/Q _4803_/X _8092_/Q _4740_/S vssd1 vssd1 vccd1 vccd1 _4804_/X
+ sky130_fd_sc_hd__o221a_1
X_4735_ _4735_/A _4735_/B vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__and2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7523_ _7474_/B _7516_/X _7522_/X _6782_/C vssd1 vssd1 vccd1 vccd1 _7524_/B sky130_fd_sc_hd__a22oi_1
XFILLER_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7454_ _7454_/A vssd1 vssd1 vccd1 vccd1 _7454_/X sky130_fd_sc_hd__buf_1
X_4666_ _4663_/X _4664_/X _4773_/A vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__a21o_1
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _8147_/D sky130_fd_sc_hd__clkbuf_1
X_6405_ _8482_/Q vssd1 vssd1 vccd1 vccd1 _6963_/A sky130_fd_sc_hd__buf_4
X_6336_ _7811_/Q _6286_/X _6335_/X vssd1 vssd1 vccd1 vccd1 _7811_/D sky130_fd_sc_hd__a21o_1
XFILLER_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8006_ _8006_/CLK _8006_/D vssd1 vssd1 vccd1 vccd1 _8006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5218_ _5338_/B _5212_/X _5217_/X vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__o21a_1
X_6198_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6198_/X sky130_fd_sc_hd__clkbuf_2
X_5149_ _8259_/Q _8251_/Q _8243_/Q _8267_/Q _5078_/X _5064_/A vssd1 vssd1 vccd1 vccd1
+ _5149_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0_0__3402_ clkbuf_0__3402_/X vssd1 vssd1 vccd1 vccd1 _6928__435/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6974__469 _6975__470/A vssd1 vssd1 vccd1 vccd1 _8150_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8504__254 vssd1 vssd1 vccd1 vccd1 partID[6] _8504__254/LO sky130_fd_sc_hd__conb_1
XFILLER_75_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3615_ clkbuf_0__3615_/X vssd1 vssd1 vccd1 vccd1 _7379__140/A sky130_fd_sc_hd__clkbuf_16
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_104 _6146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539__259 _6539__259/A vssd1 vssd1 vccd1 vccd1 _7899_/CLK sky130_fd_sc_hd__inv_2
X_4520_ _4520_/A vssd1 vssd1 vccd1 vccd1 _8181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ _8443_/Q vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__buf_2
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7170_ _8303_/Q _7211_/A _7211_/B _7193_/B _8304_/Q vssd1 vssd1 vccd1 vccd1 _7232_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4382_ _4362_/X _8232_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__mux2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6121_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6121_/X sky130_fd_sc_hd__and2_1
X_7446__19 _7447__20/A vssd1 vssd1 vccd1 vccd1 _8405_/CLK sky130_fd_sc_hd__inv_2
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6052_ _6034_/X _6050_/X _6051_/X _6037_/X vssd1 vssd1 vccd1 vccd1 _6052_/X sky130_fd_sc_hd__o211a_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _8096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5836_ _5836_/A vssd1 vssd1 vccd1 vccd1 _7732_/D sky130_fd_sc_hd__clkbuf_1
X_5767_ _4141_/X _7805_/Q _5769_/S vssd1 vssd1 vccd1 vccd1 _5768_/A sky130_fd_sc_hd__mux2_1
X_4718_ _8196_/Q _7997_/Q _7933_/Q _7893_/Q _4669_/X _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4718_/X sky130_fd_sc_hd__mux4_1
X_5698_ _5698_/A vssd1 vssd1 vccd1 vccd1 _7885_/D sky130_fd_sc_hd__clkbuf_1
X_7506_ _7577_/A _6819_/A _7510_/A _7517_/B _7505_/X vssd1 vssd1 vccd1 vccd1 _7506_/X
+ sky130_fd_sc_hd__o221a_1
X_8486_ _8496_/CLK _8486_/D vssd1 vssd1 vccd1 vccd1 _8486_/Q sky130_fd_sc_hd__dfxtp_4
X_4649_ _8166_/Q _8158_/Q _8120_/Q _8190_/Q _4648_/X _4640_/X vssd1 vssd1 vccd1 vccd1
+ _4649_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7368_ _7386_/A vssd1 vssd1 vccd1 vccd1 _7368_/X sky130_fd_sc_hd__buf_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7299_ _8308_/Q _7295_/X _7286_/X _7182_/B vssd1 vssd1 vccd1 vccd1 _7300_/B sky130_fd_sc_hd__o2bb2a_1
X_6319_ _6353_/A vssd1 vssd1 vccd1 vccd1 _6319_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _7964_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _5797_/A vssd1 vssd1 vccd1 vccd1 _5502_/B sky130_fd_sc_hd__clkbuf_4
X_6918__426 _6918__426/A vssd1 vssd1 vccd1 vccd1 _8104_/CLK sky130_fd_sc_hd__inv_2
X_3882_ _3882_/A vssd1 vssd1 vccd1 vccd1 _8470_/D sky130_fd_sc_hd__clkbuf_1
X_6670_ _6670_/A vssd1 vssd1 vccd1 vccd1 _6670_/X sky130_fd_sc_hd__buf_1
X_5621_ _7919_/Q _4973_/X _5629_/S vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__mux2_1
X_5552_ _5552_/A vssd1 vssd1 vccd1 vccd1 _7946_/D sky130_fd_sc_hd__clkbuf_1
X_8340_ _8340_/CLK _8340_/D vssd1 vssd1 vccd1 vccd1 _8340_/Q sky130_fd_sc_hd__dfxtp_1
X_8271_ _8271_/CLK _8271_/D vssd1 vssd1 vccd1 vccd1 _8271_/Q sky130_fd_sc_hd__dfxtp_1
X_4503_ _8188_/Q _4232_/X _4507_/S vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__mux2_1
X_5483_ _5483_/A vssd1 vssd1 vccd1 vccd1 _8000_/D sky130_fd_sc_hd__clkbuf_1
X_4434_ _8214_/Q _4431_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3281_ _6708_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3281_/X sky130_fd_sc_hd__clkbuf_16
X_7222_ _7246_/B _7222_/B _7222_/C _7222_/D vssd1 vssd1 vccd1 vccd1 _7270_/B sky130_fd_sc_hd__and4_1
XFILLER_116_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _4365_/X sky130_fd_sc_hd__clkbuf_2
X_7153_ _7153_/A vssd1 vssd1 vccd1 vccd1 _7305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _7756_/Q _6095_/X _6099_/X _6103_/X _6093_/X vssd1 vssd1 vccd1 vccd1 _6104_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4296_ _3931_/X _8267_/Q _4298_/S vssd1 vssd1 vccd1 vccd1 _4297_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _7813_/Q input30/X _6039_/S vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__mux2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7986_ _7986_/CLK _7986_/D vssd1 vssd1 vccd1 vccd1 _7986_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2996_ _6133_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2996_/X sky130_fd_sc_hd__clkbuf_16
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6868_ _6868_/A vssd1 vssd1 vccd1 vccd1 _8067_/D sky130_fd_sc_hd__clkbuf_1
X_5819_ _7782_/Q _5562_/A _5825_/S vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3617_ _7386_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3617_/X sky130_fd_sc_hd__clkbuf_16
X_6799_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__inv_2
XFILLER_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8469_ _8469_/CLK _8469_/D vssd1 vssd1 vccd1 vccd1 _8469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7043__525 _7043__525/A vssd1 vssd1 vccd1 vccd1 _8206_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6681__329 _6681__329/A vssd1 vssd1 vccd1 vccd1 _7993_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987__479 _6988__480/A vssd1 vssd1 vccd1 vccd1 _8160_/CLK sky130_fd_sc_hd__inv_2
Xoutput119 _5988_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput108 _7775_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
XFILLER_107_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _4150_/X sky130_fd_sc_hd__buf_2
XFILLER_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4081_ _3943_/X _8365_/Q _4081_/S vssd1 vssd1 vccd1 vccd1 _4082_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7840_ _8497_/CLK _7840_/D vssd1 vssd1 vccd1 vccd1 _7840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _4983_/A vssd1 vssd1 vccd1 vccd1 _8102_/D sky130_fd_sc_hd__clkbuf_1
X_7771_ _8490_/CLK _7771_/D vssd1 vssd1 vccd1 vccd1 _7771_/Q sky130_fd_sc_hd__dfxtp_1
X_3934_ _8445_/Q vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__buf_4
X_6593__301 _6595__303/A vssd1 vssd1 vccd1 vccd1 _7941_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3434_ clkbuf_0__3434_/X vssd1 vssd1 vccd1 vccd1 _7085__57/A sky130_fd_sc_hd__clkbuf_4
X_6653_ _6653_/A vssd1 vssd1 vccd1 vccd1 _7972_/D sky130_fd_sc_hd__clkbuf_1
X_3865_ _6310_/A _6302_/C vssd1 vssd1 vccd1 vccd1 _4108_/D sky130_fd_sc_hd__nor2_1
X_5604_ _5604_/A vssd1 vssd1 vccd1 vccd1 _7927_/D sky130_fd_sc_hd__clkbuf_1
X_6584_ _6584_/A vssd1 vssd1 vccd1 vccd1 _6584_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3402_ _6923_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3402_/X sky130_fd_sc_hd__clkbuf_16
X_5535_ _5535_/A vssd1 vssd1 vccd1 vccd1 _7977_/D sky130_fd_sc_hd__clkbuf_1
X_8323_ _8442_/CLK _8323_/D vssd1 vssd1 vccd1 vccd1 _8323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8254_ _8254_/CLK _8254_/D vssd1 vssd1 vccd1 vccd1 _8254_/Q sky130_fd_sc_hd__dfxtp_1
X_5466_ _5466_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5482_/S sky130_fd_sc_hd__nor2_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7205_ _8298_/Q _7208_/B vssd1 vssd1 vccd1 vccd1 _7206_/B sky130_fd_sc_hd__xor2_1
X_4417_ _4416_/X _8219_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5397_ _5397_/A vssd1 vssd1 vccd1 vccd1 _8043_/D sky130_fd_sc_hd__clkbuf_1
X_8185_ _8185_/CLK _8185_/D vssd1 vssd1 vccd1 vccd1 _8185_/Q sky130_fd_sc_hd__dfxtp_1
X_4348_ _4347_/X _8245_/Q _4357_/S vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4279_ _8274_/Q _4191_/X _4279_/S vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6037_/A vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _8441_/CLK _7969_/D vssd1 vssd1 vccd1 vccd1 _7969_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6581__293 _6583__295/A vssd1 vssd1 vccd1 vccd1 _7933_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5320_ _5319_/A _5322_/B _5319_/Y _5282_/X vssd1 vssd1 vccd1 vccd1 _8076_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8547__246 vssd1 vssd1 vccd1 vccd1 _8547__246/HI versionID[0] sky130_fd_sc_hd__conb_1
X_7433__8 _7434__9/A vssd1 vssd1 vccd1 vccd1 _8394_/CLK sky130_fd_sc_hd__inv_2
X_5251_ _5247_/Y _5248_/Y _5250_/Y vssd1 vssd1 vccd1 vccd1 _8081_/D sky130_fd_sc_hd__a21oi_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _8333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5182_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5334_/B sky130_fd_sc_hd__buf_2
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4133_ _5745_/A vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4064_ _4250_/A _5319_/A _5321_/A vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__nand3_4
XFILLER_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7823_ _7964_/CLK _7823_/D vssd1 vssd1 vccd1 vccd1 _7823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7754_ _8418_/CLK _7754_/D vssd1 vssd1 vccd1 vccd1 _7754_/Q sky130_fd_sc_hd__dfxtp_1
X_4966_ _4966_/A vssd1 vssd1 vccd1 vccd1 _8108_/D sky130_fd_sc_hd__clkbuf_1
X_4897_ _4926_/B _4876_/X _4883_/X _4896_/X vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__a31o_1
X_7685_ _7683_/Y _7684_/Y _7678_/X vssd1 vssd1 vccd1 vccd1 _8486_/D sky130_fd_sc_hd__a21oi_1
X_3917_ _8087_/Q vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__3417_ clkbuf_0__3417_/X vssd1 vssd1 vccd1 vccd1 _7004__493/A sky130_fd_sc_hd__clkbuf_4
X_3848_ _6008_/A _6015_/A _6015_/B vssd1 vssd1 vccd1 vccd1 _5853_/B sky130_fd_sc_hd__nor3_4
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6636_ _5922_/A _7965_/Q _6640_/S vssd1 vssd1 vccd1 vccd1 _6637_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3279_ clkbuf_0__3279_/X vssd1 vssd1 vccd1 vccd1 _6706__350/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5518_ _7984_/Q _4365_/A _5518_/S vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__mux2_1
X_8306_ _8309_/CLK _8306_/D vssd1 vssd1 vccd1 vccd1 _8306_/Q sky130_fd_sc_hd__dfxtp_1
X_6498_ _6510_/A vssd1 vssd1 vccd1 vccd1 _6498_/X sky130_fd_sc_hd__buf_1
X_8237_ _8237_/CLK _8237_/D vssd1 vssd1 vccd1 vccd1 _8237_/Q sky130_fd_sc_hd__dfxtp_1
X_5449_ _5464_/S vssd1 vssd1 vccd1 vccd1 _5458_/S sky130_fd_sc_hd__clkbuf_2
X_8168_ _8168_/CLK _8168_/D vssd1 vssd1 vccd1 vccd1 _8168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8099_ _8099_/CLK _8099_/D vssd1 vssd1 vccd1 vccd1 _8099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6960__460 _6960__460/A vssd1 vssd1 vccd1 vccd1 _8139_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7056__535 _7056__535/A vssd1 vssd1 vccd1 vccd1 _8216_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4820_ _4753_/X _8054_/Q _7938_/Q _4796_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4820_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4780_/A vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7470_ _7471_/B _7471_/C _7471_/A vssd1 vssd1 vccd1 vccd1 _7472_/C sky130_fd_sc_hd__a21oi_1
X_4682_ _6852_/B vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__clkbuf_2
X_6421_ _7662_/A vssd1 vssd1 vccd1 vccd1 _6421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6352_ _6352_/A vssd1 vssd1 vccd1 vccd1 _6371_/A sky130_fd_sc_hd__clkbuf_2
X_5303_ _5174_/X _5301_/X _5302_/X vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__o21a_1
X_8022_ _8022_/CLK _8022_/D vssd1 vssd1 vccd1 vccd1 _8022_/Q sky130_fd_sc_hd__dfxtp_1
X_5234_ _5338_/B _5232_/X _5233_/X _5336_/B vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__o211a_1
X_6588__299 _6588__299/A vssd1 vssd1 vccd1 vccd1 _7939_/CLK sky130_fd_sc_hd__inv_2
X_5165_ _8069_/Q _5196_/S vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__or2_1
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _8125_/Q vssd1 vssd1 vccd1 vccd1 _4120_/B sky130_fd_sc_hd__inv_2
X_5096_ _5048_/X _5094_/X _5278_/A vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3280_ clkbuf_0__3280_/X vssd1 vssd1 vccd1 vccd1 _6726_/A sky130_fd_sc_hd__clkbuf_4
X_4047_ _4062_/S vssd1 vssd1 vccd1 vccd1 _4056_/S sky130_fd_sc_hd__buf_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _7806_/CLK _7806_/D vssd1 vssd1 vccd1 vccd1 _7806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5998_ _6080_/A vssd1 vssd1 vccd1 vccd1 _6061_/A sky130_fd_sc_hd__buf_2
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4949_ _4949_/A vssd1 vssd1 vccd1 vccd1 _8115_/D sky130_fd_sc_hd__clkbuf_1
X_7737_ _8308_/CLK _7737_/D vssd1 vssd1 vccd1 vccd1 _7737_/Q sky130_fd_sc_hd__dfxtp_1
X_7668_ _5913_/A _7657_/X _7660_/Y vssd1 vssd1 vccd1 vccd1 _7668_/X sky130_fd_sc_hd__a21o_1
X_6619_ _6619_/A vssd1 vssd1 vccd1 vccd1 _7957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _7599_/A vssd1 vssd1 vccd1 vccd1 _8442_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2995_ clkbuf_0__2995_/X vssd1 vssd1 vccd1 vccd1 _6497_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3616_ clkbuf_0__3616_/X vssd1 vssd1 vccd1 vccd1 _7385__145/A sky130_fd_sc_hd__clkbuf_4
X_6905__417 _6906__418/A vssd1 vssd1 vccd1 vccd1 _8095_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6845__386 _6846__387/A vssd1 vssd1 vccd1 vccd1 _8054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970_ _6970_/A vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__buf_1
X_5921_ _5921_/A vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6702__346 _6703__347/A vssd1 vssd1 vccd1 vccd1 _8010_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ _6473_/A _5853_/C vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__nand2_1
X_5783_ _7798_/Q _4347_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__mux2_1
X_4803_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4734_ _7780_/Q _7900_/Q _7908_/Q _7948_/Q _4648_/A _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4735_/B sky130_fd_sc_hd__mux4_1
X_7522_ _7557_/B vssd1 vssd1 vccd1 vccd1 _7522_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _4665_/A vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__clkbuf_2
X_4596_ _8147_/Q _4442_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__mux2_1
X_6404_ _7824_/Q _6401_/X _6393_/X _6403_/X _6391_/X vssd1 vssd1 vccd1 vccd1 _7824_/D
+ sky130_fd_sc_hd__a221o_1
X_6258__195 _6258__195/A vssd1 vssd1 vccd1 vccd1 _7787_/CLK sky130_fd_sc_hd__inv_2
X_6335_ _6289_/A _6332_/X _6334_/X _6369_/A vssd1 vssd1 vccd1 vccd1 _6335_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8005_ _8005_/CLK _8005_/D vssd1 vssd1 vccd1 vccd1 _8005_/Q sky130_fd_sc_hd__dfxtp_1
X_6266_ _6278_/A vssd1 vssd1 vccd1 vccd1 _6266_/X sky130_fd_sc_hd__buf_1
X_5217_ _8265_/Q _5214_/X _5216_/X _8257_/Q _5038_/A vssd1 vssd1 vccd1 vccd1 _5217_/X
+ sky130_fd_sc_hd__o221a_1
X_6197_ _6328_/A vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__clkbuf_2
X_5148_ _8377_/Q _8275_/Q _8012_/Q _8227_/Q _5111_/A _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5148_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3401_ clkbuf_0__3401_/X vssd1 vssd1 vccd1 vccd1 _6922__430/A sky130_fd_sc_hd__clkbuf_4
X_5079_ _8262_/Q _8254_/Q _8246_/Q _8270_/Q _5078_/X _5070_/X vssd1 vssd1 vccd1 vccd1
+ _5079_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_105 _7680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A vssd1 vssd1 vccd1 vccd1 _8209_/D sky130_fd_sc_hd__clkbuf_1
X_7381__141 _7385__145/A vssd1 vssd1 vccd1 vccd1 _8352_/CLK sky130_fd_sc_hd__inv_2
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _8233_/D sky130_fd_sc_hd__clkbuf_1
X_6120_ _7762_/Q _6111_/X _6112_/X _6119_/X _6109_/X vssd1 vssd1 vccd1 vccd1 _6120_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6051_ _7742_/Q _6063_/B vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__or2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _4404_/X _8096_/Q _5010_/S vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5904_ _7684_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__or2_1
XFILLER_81_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5835_ _4101_/X _7732_/Q _5843_/S vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5766_ _5766_/A vssd1 vssd1 vccd1 vccd1 _7806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4717_ _4715_/X _4716_/X _4665_/A vssd1 vssd1 vccd1 vccd1 _4717_/X sky130_fd_sc_hd__a21o_1
X_5697_ _7885_/Q _4981_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__mux2_1
X_7505_ _7508_/A _8413_/Q _7510_/A vssd1 vssd1 vccd1 vccd1 _7505_/X sky130_fd_sc_hd__or3b_1
X_8485_ _8498_/CLK _8485_/D vssd1 vssd1 vccd1 vccd1 _8485_/Q sky130_fd_sc_hd__dfxtp_1
X_4648_ _4648_/A vssd1 vssd1 vccd1 vccd1 _4648_/X sky130_fd_sc_hd__clkbuf_4
X_7436_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7436_/X sky130_fd_sc_hd__buf_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _4579_/A vssd1 vssd1 vccd1 vccd1 _8155_/D sky130_fd_sc_hd__clkbuf_1
X_7298_ _7321_/A vssd1 vssd1 vccd1 vccd1 _7309_/A sky130_fd_sc_hd__clkbuf_2
X_6318_ _6318_/A vssd1 vssd1 vccd1 vccd1 _6318_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980__474 _6981__475/A vssd1 vssd1 vccd1 vccd1 _8155_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7133__96 _7134__97/A vssd1 vssd1 vccd1 vccd1 _8277_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7451__23 _7453__25/A vssd1 vssd1 vccd1 vccd1 _8409_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6545__264 _6546__265/A vssd1 vssd1 vccd1 vccd1 _7904_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _6892_/A _5321_/B vssd1 vssd1 vccd1 vccd1 _5797_/A sky130_fd_sc_hd__nand2_2
X_3881_ _8470_/Q _3880_/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__mux2_1
X_5620_ _5635_/S vssd1 vssd1 vccd1 vccd1 _5629_/S sky130_fd_sc_hd__buf_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5551_ _7946_/Q _4990_/X _5555_/S vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8270_ _8270_/CLK _8270_/D vssd1 vssd1 vccd1 vccd1 _8270_/Q sky130_fd_sc_hd__dfxtp_1
X_4502_ _4502_/A vssd1 vssd1 vccd1 vccd1 _8189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5482_ _8000_/Q _4365_/A _5482_/S vssd1 vssd1 vccd1 vccd1 _5483_/A sky130_fd_sc_hd__mux2_1
X_7221_ _7186_/X _7187_/Y _7192_/Y _7210_/X _7220_/X vssd1 vssd1 vccd1 vccd1 _7222_/D
+ sky130_fd_sc_hd__o2111a_1
X_4433_ _4455_/S vssd1 vssd1 vccd1 vccd1 _4446_/S sky130_fd_sc_hd__buf_2
Xclkbuf_0__3280_ _6707_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3280_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4364_ _4364_/A vssd1 vssd1 vccd1 vccd1 _8240_/D sky130_fd_sc_hd__clkbuf_1
X_7152_ _8311_/Q _8310_/Q _7158_/B vssd1 vssd1 vccd1 vccd1 _7153_/A sky130_fd_sc_hd__nand3_1
X_6103_ _6103_/A _6105_/B vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__and2_4
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4295_ _4295_/A vssd1 vssd1 vccd1 vccd1 _8268_/D sky130_fd_sc_hd__clkbuf_1
X_7083_ _7083_/A vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__buf_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6034_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7985_ _7985_/CLK _7985_/D vssd1 vssd1 vccd1 vccd1 _7985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2995_ _6132_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2995_/X sky130_fd_sc_hd__clkbuf_16
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7388__147 _7389__148/A vssd1 vssd1 vccd1 vccd1 _8358_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6867_ _8441_/Q _6963_/C vssd1 vssd1 vccd1 vccd1 _6868_/A sky130_fd_sc_hd__and2_1
X_5818_ _5818_/A vssd1 vssd1 vccd1 vccd1 _7783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6798_ _8489_/Q _7461_/B vssd1 vssd1 vccd1 vccd1 _6803_/A sky130_fd_sc_hd__xor2_1
X_5749_ _7862_/Q _5562_/A _5755_/S vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3616_ _7380_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3616_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8468_ _8468_/CLK _8468_/D vssd1 vssd1 vccd1 vccd1 _8468_/Q sky130_fd_sc_hd__dfxtp_1
X_8399_ _8399_/CLK _8399_/D vssd1 vssd1 vccd1 vccd1 _8399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6488__218 _6488__218/A vssd1 vssd1 vccd1 vccd1 _7858_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3229_ clkbuf_0__3229_/X vssd1 vssd1 vccd1 vccd1 _6549__267/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput109 _5946_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924__431 _6926__433/A vssd1 vssd1 vccd1 vccd1 _8109_/CLK sky130_fd_sc_hd__inv_2
X_4080_ _4080_/A vssd1 vssd1 vccd1 vccd1 _8366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _8102_/Q _4981_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__mux2_1
X_7770_ _8498_/CLK _7770_/D vssd1 vssd1 vccd1 vccd1 _7770_/Q sky130_fd_sc_hd__dfxtp_1
X_3933_ _3933_/A vssd1 vssd1 vccd1 vccd1 _8454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8478_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__3433_ clkbuf_0__3433_/X vssd1 vssd1 vccd1 vccd1 _7082__55/A sky130_fd_sc_hd__clkbuf_4
X_6652_ _7972_/Q _5937_/A _6652_/S vssd1 vssd1 vccd1 vccd1 _6653_/A sky130_fd_sc_hd__mux2_1
X_3864_ _7839_/Q _7840_/Q _7652_/A _7831_/Q vssd1 vssd1 vccd1 vccd1 _6302_/C sky130_fd_sc_hd__or4b_1
XFILLER_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5603_ _5557_/X _7927_/Q _5611_/S vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3401_ _6917_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3401_/X sky130_fd_sc_hd__clkbuf_16
X_8322_ _8442_/CLK _8322_/D vssd1 vssd1 vccd1 vccd1 _8322_/Q sky130_fd_sc_hd__dfxtp_1
X_5534_ _5369_/X _7977_/Q _5536_/S vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__mux2_1
X_8253_ _8253_/CLK _8253_/D vssd1 vssd1 vccd1 vccd1 _8253_/Q sky130_fd_sc_hd__dfxtp_1
X_5465_ _5465_/A vssd1 vssd1 vccd1 vccd1 _8008_/D sky130_fd_sc_hd__clkbuf_1
X_8184_ _8184_/CLK _8184_/D vssd1 vssd1 vccd1 vccd1 _8184_/Q sky130_fd_sc_hd__dfxtp_1
X_7204_ _8297_/Q vssd1 vssd1 vccd1 vccd1 _7208_/B sky130_fd_sc_hd__clkbuf_2
X_4416_ _8064_/Q vssd1 vssd1 vccd1 vccd1 _4416_/X sky130_fd_sc_hd__clkbuf_2
X_5396_ _5343_/X _8043_/Q _5404_/S vssd1 vssd1 vccd1 vccd1 _5397_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4347_ _4347_/A vssd1 vssd1 vccd1 vccd1 _4347_/X sky130_fd_sc_hd__buf_2
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4278_ _4278_/A vssd1 vssd1 vccd1 vccd1 _8275_/D sky130_fd_sc_hd__clkbuf_1
X_7394__151 _7396__153/A vssd1 vssd1 vccd1 vccd1 _8362_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6017_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6037_/A sky130_fd_sc_hd__buf_4
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6602__309 _6603__310/A vssd1 vssd1 vccd1 vccd1 _7949_/CLK sky130_fd_sc_hd__inv_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7968_ _8441_/CLK _7968_/D vssd1 vssd1 vccd1 vccd1 _7968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7899_ _7899_/CLK _7899_/D vssd1 vssd1 vccd1 vccd1 _7899_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6993__484 _6994__485/A vssd1 vssd1 vccd1 vccd1 _8165_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5250_ _3937_/X _5022_/A _5249_/X vssd1 vssd1 vccd1 vccd1 _5250_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ _8333_/Q _4200_/X _4201_/S vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5174_/X _5177_/X _5180_/X vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4132_ _4904_/A _4903_/B _4405_/B vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__or3_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _8373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7822_ _8496_/CLK _7822_/D vssd1 vssd1 vccd1 vccd1 _7822_/Q sky130_fd_sc_hd__dfxtp_1
X_4965_ _8108_/Q _4238_/X _4965_/S vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__mux2_1
X_7753_ _7964_/CLK _7753_/D vssd1 vssd1 vccd1 vccd1 _7753_/Q sky130_fd_sc_hd__dfxtp_1
X_3916_ _8449_/Q vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1_0__3416_ clkbuf_0__3416_/X vssd1 vssd1 vccd1 vccd1 _7000__490/A sky130_fd_sc_hd__clkbuf_4
X_4896_ _4883_/A _4886_/X _4889_/X _4895_/X _4622_/A vssd1 vssd1 vccd1 vccd1 _4896_/X
+ sky130_fd_sc_hd__o311a_1
X_7684_ _7684_/A _7693_/B vssd1 vssd1 vccd1 vccd1 _7684_/Y sky130_fd_sc_hd__nand2_1
X_3847_ _3847_/A _3847_/B _3847_/C vssd1 vssd1 vccd1 vccd1 _6015_/B sky130_fd_sc_hd__or3_4
X_6635_ _6635_/A vssd1 vssd1 vccd1 vccd1 _7964_/D sky130_fd_sc_hd__clkbuf_1
X_6566_ _6578_/A vssd1 vssd1 vccd1 vccd1 _6566_/X sky130_fd_sc_hd__buf_1
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3278_ clkbuf_0__3278_/X vssd1 vssd1 vccd1 vccd1 _6698__343/A sky130_fd_sc_hd__clkbuf_4
X_5517_ _5517_/A vssd1 vssd1 vccd1 vccd1 _7985_/D sky130_fd_sc_hd__clkbuf_1
X_8305_ _8309_/CLK _8305_/D vssd1 vssd1 vccd1 vccd1 _8305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8236_ _8236_/CLK _8236_/D vssd1 vssd1 vccd1 vccd1 _8236_/Q sky130_fd_sc_hd__dfxtp_1
X_6497_ _6497_/A vssd1 vssd1 vccd1 vccd1 _6497_/X sky130_fd_sc_hd__buf_1
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5448_ _5466_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5464_/S sky130_fd_sc_hd__nor2_4
X_5379_ _5379_/A vssd1 vssd1 vccd1 vccd1 _8051_/D sky130_fd_sc_hd__clkbuf_1
X_8167_ _8167_/CLK _8167_/D vssd1 vssd1 vccd1 vccd1 _8167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8098_ _8098_/CLK _8098_/D vssd1 vssd1 vccd1 vccd1 _8098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7642__48 _7643__49/A vssd1 vssd1 vccd1 vccd1 _8471_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _8123_/Q vssd1 vssd1 vccd1 vccd1 _4780_/A sky130_fd_sc_hd__inv_2
X_8514__213 vssd1 vssd1 vccd1 vccd1 _8514__213/HI core0Index[0] sky130_fd_sc_hd__conb_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4681_ _6854_/A vssd1 vssd1 vccd1 vccd1 _6852_/B sky130_fd_sc_hd__clkbuf_2
X_6420_ _6480_/A vssd1 vssd1 vccd1 vccd1 _7662_/A sky130_fd_sc_hd__clkbuf_2
X_6351_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _6792_/A sky130_fd_sc_hd__buf_4
X_5302_ _8223_/Q _5227_/X _5285_/B _8373_/Q _5062_/A vssd1 vssd1 vccd1 vccd1 _5302_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3063_ clkbuf_0__3063_/X vssd1 vssd1 vccd1 vccd1 _6282__214/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5233_ _8452_/Q _5163_/X _5216_/X _8460_/Q vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__o22a_1
X_8021_ _8021_/CLK _8021_/D vssd1 vssd1 vccd1 vccd1 _8021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5164_ _5164_/A _5175_/A vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ _4607_/A _4113_/Y _4114_/Y vssd1 vssd1 vccd1 vccd1 _4129_/A sky130_fd_sc_hd__a21oi_1
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5095_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4046_ _4083_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _4062_/S sky130_fd_sc_hd__nor2_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7805_ _7805_/CLK _7805_/D vssd1 vssd1 vccd1 vccd1 _7805_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _6000_/A _5854_/X _7724_/Q vssd1 vssd1 vccd1 vccd1 _6080_/A sky130_fd_sc_hd__a21oi_1
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4948_ _8115_/Q _4241_/X _4952_/S vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__mux2_1
X_7736_ _8308_/CLK _7736_/D vssd1 vssd1 vccd1 vccd1 _7736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4879_ _7888_/Q _4755_/A _4878_/X vssd1 vssd1 vccd1 vccd1 _4883_/B sky130_fd_sc_hd__o21a_1
X_7667_ _8481_/Q _7656_/X _7666_/X _7662_/X vssd1 vssd1 vccd1 vccd1 _8481_/D sky130_fd_sc_hd__o211a_1
X_6618_ _7684_/A _7957_/Q _6622_/S vssd1 vssd1 vccd1 vccd1 _6619_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7598_ _7598_/A _7604_/B _7598_/C vssd1 vssd1 vccd1 vccd1 _7599_/A sky130_fd_sc_hd__and3_1
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2994_ clkbuf_0__2994_/X vssd1 vssd1 vccd1 vccd1 _7454_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8219_ _8219_/CLK _8219_/D vssd1 vssd1 vccd1 vccd1 _8219_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3229_ _6547_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3229_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7085__57 _7085__57/A vssd1 vssd1 vccd1 vccd1 _8238_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7409__164 _7409__164/A vssd1 vssd1 vccd1 vccd1 _8375_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7062__540 _7062__540/A vssd1 vssd1 vccd1 vccd1 _8221_/CLK sky130_fd_sc_hd__inv_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6509__235 _6509__235/A vssd1 vssd1 vccd1 vccd1 _7875_/CLK sky130_fd_sc_hd__inv_2
X_5920_ _5920_/A _5928_/B vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__or2_4
XFILLER_80_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5851_ _7974_/Q _7975_/Q _7972_/Q _7973_/Q vssd1 vssd1 vccd1 vccd1 _5853_/C sky130_fd_sc_hd__and4bb_2
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5782_ _5782_/A vssd1 vssd1 vccd1 vccd1 _7799_/D sky130_fd_sc_hd__clkbuf_1
X_4802_ _4801_/X _7979_/Q _7883_/Q _4769_/X _4794_/A vssd1 vssd1 vccd1 vccd1 _4802_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _4627_/A _4730_/X _4732_/X vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__a21o_1
X_7521_ _7554_/A vssd1 vssd1 vccd1 vccd1 _7534_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ _7927_/Q _7807_/Q _7732_/Q _7919_/Q _4640_/A _4638_/X vssd1 vssd1 vccd1 vccd1
+ _4664_/X sky130_fd_sc_hd__mux4_1
X_6403_ _8483_/Q _6408_/B _6410_/C vssd1 vssd1 vccd1 vccd1 _6403_/X sky130_fd_sc_hd__and3_1
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _8148_/D sky130_fd_sc_hd__clkbuf_1
X_6334_ _8476_/Q _6311_/X _6333_/X _6306_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _6334_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _6497_/A vssd1 vssd1 vccd1 vccd1 _6265_/X sky130_fd_sc_hd__buf_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8004_ _8004_/CLK _8004_/D vssd1 vssd1 vccd1 vccd1 _8004_/Q sky130_fd_sc_hd__dfxtp_1
X_5216_ _5239_/B vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6196_ _7968_/Q _6194_/X _6195_/X _6188_/X _7757_/Q vssd1 vssd1 vccd1 vccd1 _7757_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5147_ _5099_/X _5144_/X _5146_/X vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3400_ clkbuf_0__3400_/X vssd1 vssd1 vccd1 vccd1 _6942_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5078_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__buf_2
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4029_ _8388_/Q _3992_/X _4037_/S vssd1 vssd1 vccd1 vccd1 _4030_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7719_ _7722_/A _7719_/B vssd1 vssd1 vccd1 vccd1 _7720_/A sky130_fd_sc_hd__or2_1
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6718__354 _6718__354/A vssd1 vssd1 vccd1 vccd1 _8021_/CLK sky130_fd_sc_hd__inv_2
X_6911__422 _6911__422/A vssd1 vssd1 vccd1 vccd1 _8100_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_106 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6851__391 _6851__391/A vssd1 vssd1 vccd1 vccd1 _8059_/CLK sky130_fd_sc_hd__inv_2
X_4380_ _4359_/X _8233_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6050_ _7817_/Q input34/X _6058_/S vssd1 vssd1 vccd1 vccd1 _6050_/X sky130_fd_sc_hd__mux2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5016_/S vssd1 vssd1 vccd1 vccd1 _5010_/S sky130_fd_sc_hd__buf_2
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5903_ _5903_/A vssd1 vssd1 vccd1 vccd1 _5903_/X sky130_fd_sc_hd__clkbuf_1
X_5834_ _5849_/S vssd1 vssd1 vccd1 vccd1 _5843_/S sky130_fd_sc_hd__buf_2
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5765_ _4138_/X _7806_/Q _5769_/S vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4716_ _7925_/Q _7805_/Q _7730_/Q _7917_/Q _4640_/A _4638_/X vssd1 vssd1 vccd1 vccd1
+ _4716_/X sky130_fd_sc_hd__mux4_1
X_5696_ _5696_/A vssd1 vssd1 vccd1 vccd1 _7886_/D sky130_fd_sc_hd__clkbuf_1
X_8484_ _8496_/CLK _8484_/D vssd1 vssd1 vccd1 vccd1 _8484_/Q sky130_fd_sc_hd__dfxtp_4
X_7504_ _7504_/A _7508_/B vssd1 vssd1 vccd1 vccd1 _7517_/B sky130_fd_sc_hd__nand2_2
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4647_ _4650_/A vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6317_ _8498_/Q _6293_/X _6299_/X vssd1 vssd1 vccd1 vccd1 _6317_/X sky130_fd_sc_hd__a21o_1
X_4578_ _4416_/X _8155_/Q _4580_/S vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7297_ _7297_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _8307_/D sky130_fd_sc_hd__nor2_1
X_6179_ _6176_/X _7958_/Q _6178_/X _6172_/X _7747_/Q vssd1 vssd1 vccd1 vccd1 _7747_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8499_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3880_ _8446_/Q vssd1 vssd1 vccd1 vccd1 _3880_/X sky130_fd_sc_hd__buf_2
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _5550_/A vssd1 vssd1 vccd1 vccd1 _7947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5481_ _5481_/A vssd1 vssd1 vccd1 vccd1 _8001_/D sky130_fd_sc_hd__clkbuf_1
X_4501_ _8189_/Q _4229_/X _4507_/S vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__mux2_1
X_4432_ _4457_/A _5430_/B vssd1 vssd1 vccd1 vccd1 _4455_/S sky130_fd_sc_hd__nor2_4
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7220_ _7213_/Y _7214_/X _7216_/X _7218_/X _7219_/X vssd1 vssd1 vccd1 vccd1 _7220_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_113_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4363_ _4362_/X _8240_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7151_ _8309_/Q _7176_/A _7173_/A _7193_/D vssd1 vssd1 vccd1 vccd1 _7158_/B sky130_fd_sc_hd__and4_1
X_4294_ _3928_/X _8268_/Q _4298_/S vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _7755_/Q _6095_/X _6099_/X _6101_/X _6093_/X vssd1 vssd1 vccd1 vccd1 _6102_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6033_ _6009_/X _6031_/X _6032_/X _6018_/X vssd1 vssd1 vccd1 vccd1 _6033_/X sky130_fd_sc_hd__o211a_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7984_ _7984_/CLK _7984_/D vssd1 vssd1 vccd1 vccd1 _7984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6935_ _6942_/A vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__buf_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2994_ _6131_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2994_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6866_ _6866_/A vssd1 vssd1 vccd1 vccd1 _8066_/D sky130_fd_sc_hd__clkbuf_1
X_5817_ _7783_/Q _5557_/A _5825_/S vssd1 vssd1 vccd1 vccd1 _5818_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6797_ _8425_/Q _6797_/B vssd1 vssd1 vccd1 vccd1 _7461_/B sky130_fd_sc_hd__xor2_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3615_ _7374_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3615_/X sky130_fd_sc_hd__clkbuf_16
X_5748_ _5748_/A vssd1 vssd1 vccd1 vccd1 _7863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5679_ _7893_/Q _4981_/X _5683_/S vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__mux2_1
X_8467_ _8467_/CLK _8467_/D vssd1 vssd1 vccd1 vccd1 _8467_/Q sky130_fd_sc_hd__dfxtp_1
X_8398_ _8398_/CLK _8398_/D vssd1 vssd1 vccd1 vccd1 _8398_/Q sky130_fd_sc_hd__dfxtp_1
X_7349_ _7349_/A vssd1 vssd1 vccd1 vccd1 _7349_/X sky130_fd_sc_hd__buf_1
XFILLER_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3228_ clkbuf_0__3228_/X vssd1 vssd1 vccd1 vccd1 _6546__265/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7106__75 _7106__75/A vssd1 vssd1 vccd1 vccd1 _8256_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _8065_/Q vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _3931_/X _8454_/Q _3935_/S vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__mux2_1
X_6720_ _6726_/A vssd1 vssd1 vccd1 vccd1 _6720_/X sky130_fd_sc_hd__buf_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3432_ clkbuf_0__3432_/X vssd1 vssd1 vccd1 vccd1 _7083_/A sky130_fd_sc_hd__clkbuf_4
X_6651_ _6651_/A vssd1 vssd1 vccd1 vccd1 _7971_/D sky130_fd_sc_hd__clkbuf_1
X_3863_ _8016_/Q _6291_/A vssd1 vssd1 vccd1 vccd1 _6310_/A sky130_fd_sc_hd__nand2_1
X_5602_ _5617_/S vssd1 vssd1 vccd1 vccd1 _5611_/S sky130_fd_sc_hd__buf_2
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533_ _5533_/A vssd1 vssd1 vccd1 vccd1 _7978_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3400_ _6916_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3400_/X sky130_fd_sc_hd__clkbuf_16
X_8321_ _8442_/CLK _8321_/D vssd1 vssd1 vccd1 vccd1 _8321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8252_ _8252_/CLK _8252_/D vssd1 vssd1 vccd1 vccd1 _8252_/Q sky130_fd_sc_hd__dfxtp_1
X_5464_ _8008_/Q _4454_/X _5464_/S vssd1 vssd1 vccd1 vccd1 _5465_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5395_ _5410_/S vssd1 vssd1 vccd1 vccd1 _5404_/S sky130_fd_sc_hd__clkbuf_4
X_8183_ _8183_/CLK _8183_/D vssd1 vssd1 vccd1 vccd1 _8183_/Q sky130_fd_sc_hd__dfxtp_1
X_7203_ _7273_/A _7273_/B _6774_/A vssd1 vssd1 vccd1 vccd1 _7203_/Y sky130_fd_sc_hd__a21oi_1
X_4415_ _4415_/A vssd1 vssd1 vccd1 vccd1 _8220_/D sky130_fd_sc_hd__clkbuf_1
X_4346_ _4346_/A vssd1 vssd1 vccd1 vccd1 _8246_/D sky130_fd_sc_hd__clkbuf_1
X_4277_ _8275_/Q _4188_/X _4279_/S vssd1 vssd1 vccd1 vccd1 _4278_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6016_ _6016_/A vssd1 vssd1 vccd1 vccd1 _6109_/A sky130_fd_sc_hd__buf_2
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7967_ _8060_/CLK _7967_/D vssd1 vssd1 vccd1 vccd1 _7967_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7898_ _7898_/CLK _7898_/D vssd1 vssd1 vccd1 vccd1 _7898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6494__223 _6494__223/A vssd1 vssd1 vccd1 vccd1 _7863_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6871__394 _6872__395/A vssd1 vssd1 vccd1 vccd1 _8070_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7403__159 _7404__160/A vssd1 vssd1 vccd1 vccd1 _8370_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _8442_/Q vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5180_ _8178_/Q _5178_/X _5179_/X _8170_/Q _5037_/A vssd1 vssd1 vccd1 vccd1 _5180_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4131_ _4680_/A _4911_/C vssd1 vssd1 vccd1 vccd1 _4405_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4062_ _8373_/Q _4022_/X _4062_/S vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7821_ _8496_/CLK _7821_/D vssd1 vssd1 vccd1 vccd1 _7821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4964_ _4964_/A vssd1 vssd1 vccd1 vccd1 _8109_/D sky130_fd_sc_hd__clkbuf_1
X_7752_ _7964_/CLK _7752_/D vssd1 vssd1 vccd1 vccd1 _7752_/Q sky130_fd_sc_hd__dfxtp_1
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _8458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4895_ _4890_/X _4891_/X _4773_/A _4894_/X vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__a211o_1
X_7683_ _7683_/A _7692_/B vssd1 vssd1 vccd1 vccd1 _7683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3415_ clkbuf_0__3415_/X vssd1 vssd1 vccd1 vccd1 _6994__485/A sky130_fd_sc_hd__clkbuf_4
X_6558__275 _6558__275/A vssd1 vssd1 vccd1 vccd1 _7915_/CLK sky130_fd_sc_hd__inv_2
X_3846_ _3846_/A _3846_/B _3846_/C _3846_/D vssd1 vssd1 vccd1 vccd1 _3847_/C sky130_fd_sc_hd__or4_1
XFILLER_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6634_ _5920_/A _7964_/Q _6634_/S vssd1 vssd1 vccd1 vccd1 _6635_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3277_ clkbuf_0__3277_/X vssd1 vssd1 vccd1 vccd1 _6694__340/A sky130_fd_sc_hd__clkbuf_4
X_5516_ _7985_/Q _4362_/A _5518_/S vssd1 vssd1 vccd1 vccd1 _5517_/A sky130_fd_sc_hd__mux2_1
X_8304_ _8309_/CLK _8304_/D vssd1 vssd1 vccd1 vccd1 _8304_/Q sky130_fd_sc_hd__dfxtp_1
X_8235_ _8235_/CLK _8235_/D vssd1 vssd1 vccd1 vccd1 _8235_/Q sky130_fd_sc_hd__dfxtp_1
X_5447_ _5447_/A vssd1 vssd1 vccd1 vccd1 _8019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3631_ clkbuf_0__3631_/X vssd1 vssd1 vccd1 vccd1 _7619__29/A sky130_fd_sc_hd__clkbuf_4
X_5378_ _5343_/X _8051_/Q _5386_/S vssd1 vssd1 vccd1 vccd1 _5379_/A sky130_fd_sc_hd__mux2_1
X_8166_ _8166_/CLK _8166_/D vssd1 vssd1 vccd1 vccd1 _8166_/Q sky130_fd_sc_hd__dfxtp_1
X_4329_ _4329_/A vssd1 vssd1 vccd1 vccd1 _8253_/D sky130_fd_sc_hd__clkbuf_1
X_8097_ _8097_/CLK _8097_/D vssd1 vssd1 vccd1 vccd1 _8097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _4680_/A vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__buf_2
X_6350_ _7813_/Q _6343_/X _6349_/X vssd1 vssd1 vccd1 vccd1 _7813_/D sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0__3062_ clkbuf_0__3062_/X vssd1 vssd1 vccd1 vccd1 _6277__210/A sky130_fd_sc_hd__clkbuf_4
X_5301_ _8271_/Q _8008_/Q _5301_/S vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8020_ _8020_/CLK _8020_/D vssd1 vssd1 vccd1 vccd1 _8020_/Q sky130_fd_sc_hd__dfxtp_1
X_5232_ _7986_/Q _8021_/Q _5235_/S vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _8128_/Q _8123_/Q vssd1 vssd1 vccd1 vccd1 _4114_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _8395_/Q _8387_/Q _7790_/Q _8403_/Q _5294_/S _5064_/X vssd1 vssd1 vccd1 vccd1
+ _5094_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4250_/A _4287_/B _5321_/A vssd1 vssd1 vccd1 vccd1 _5448_/B sky130_fd_sc_hd__or3_4
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7804_ _7804_/CLK _7804_/D vssd1 vssd1 vccd1 vccd1 _7804_/Q sky130_fd_sc_hd__dfxtp_1
X_5996_ _5996_/A vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__clkbuf_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937__442 _6937__442/A vssd1 vssd1 vccd1 vccd1 _8120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4947_ _4947_/A vssd1 vssd1 vccd1 vccd1 _8116_/D sky130_fd_sc_hd__clkbuf_1
X_7735_ _8308_/CLK _7735_/D vssd1 vssd1 vccd1 vccd1 _7735_/Q sky130_fd_sc_hd__dfxtp_1
X_4878_ _8191_/Q _4814_/A _4776_/A _4877_/X _4659_/A vssd1 vssd1 vccd1 vccd1 _4878_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7666_ _5915_/A _7657_/X _7660_/Y vssd1 vssd1 vccd1 vccd1 _7666_/X sky130_fd_sc_hd__a21o_1
X_6617_ _6617_/A vssd1 vssd1 vccd1 vccd1 _7956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3829_ _5019_/A _5316_/A vssd1 vssd1 vccd1 vccd1 _3838_/B sky130_fd_sc_hd__and2b_1
XFILLER_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7597_ _7597_/A _7675_/B vssd1 vssd1 vccd1 vccd1 _7598_/C sky130_fd_sc_hd__and2_1
XFILLER_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _6343_/A _6415_/X _6474_/Y _6419_/X vssd1 vssd1 vccd1 vccd1 _6480_/C sky130_fd_sc_hd__o31a_1
X_8218_ _8218_/CLK _8218_/D vssd1 vssd1 vccd1 vccd1 _8218_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3228_ _6541_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3228_/X sky130_fd_sc_hd__clkbuf_16
X_8149_ _8149_/CLK _8149_/D vssd1 vssd1 vccd1 vccd1 _8149_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3614_ clkbuf_0__3614_/X vssd1 vssd1 vccd1 vccd1 _7370__132/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_0 _7775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8537__236 vssd1 vssd1 vccd1 vccd1 _8537__236/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ _5850_/A vssd1 vssd1 vccd1 vccd1 _7725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5781_ _7799_/Q _4342_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__mux2_1
X_4801_ _4801_/A vssd1 vssd1 vccd1 vccd1 _4801_/X sky130_fd_sc_hd__clkbuf_2
X_4732_ _4663_/X _4731_/X _4644_/X vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7520_ _7535_/A vssd1 vssd1 vccd1 vccd1 _7554_/A sky130_fd_sc_hd__clkbuf_2
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _4663_/X sky130_fd_sc_hd__buf_2
X_6402_ _8018_/Q vssd1 vssd1 vccd1 vccd1 _6410_/C sky130_fd_sc_hd__clkbuf_1
X_4594_ _8148_/Q _4439_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6333_ _8136_/Q _6318_/X _6319_/X vssd1 vssd1 vccd1 vccd1 _6333_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8003_ _8003_/CLK _8003_/D vssd1 vssd1 vccd1 vccd1 _8003_/Q sky130_fd_sc_hd__dfxtp_1
X_5215_ _5215_/A vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__buf_2
X_6195_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5146_ _5160_/A _5145_/X _5113_/X vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _5074_/X _5076_/X _5202_/A vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7039__521 _7041__523/A vssd1 vssd1 vccd1 vccd1 _8202_/CLK sky130_fd_sc_hd__inv_2
X_4028_ _4043_/S vssd1 vssd1 vccd1 vccd1 _4037_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7137__100 _7136__99/A vssd1 vssd1 vccd1 vccd1 _8281_/CLK sky130_fd_sc_hd__inv_2
X_7090__61 _7092__63/A vssd1 vssd1 vccd1 vccd1 _8242_/CLK sky130_fd_sc_hd__inv_2
X_5979_ _5979_/A vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7718_ _8498_/Q _7601_/C _7721_/S vssd1 vssd1 vccd1 vccd1 _7719_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7649_ _7649_/A _7649_/B vssd1 vssd1 vccd1 vccd1 _8477_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7620__30 _7620__30/A vssd1 vssd1 vccd1 vccd1 _8453_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_107 _7503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6515__240 _6515__240/A vssd1 vssd1 vccd1 vccd1 _7880_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6138__179 _6138__179/A vssd1 vssd1 vccd1 vccd1 _7728_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5000_ _5601_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5016_/S sky130_fd_sc_hd__or2_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5902_ _5902_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__or2_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5833_ _5833_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5849_/S sky130_fd_sc_hd__or2_2
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3631_ _7455_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3631_/X sky130_fd_sc_hd__clkbuf_16
X_5764_ _5764_/A vssd1 vssd1 vccd1 vccd1 _7807_/D sky130_fd_sc_hd__clkbuf_1
X_7503_ _7503_/A input1/X vssd1 vssd1 vccd1 vccd1 _7510_/A sky130_fd_sc_hd__or2_1
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__clkbuf_2
X_5695_ _7886_/Q _4978_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5696_/A sky130_fd_sc_hd__mux2_1
X_8483_ _8483_/CLK _8483_/D vssd1 vssd1 vccd1 vccd1 _8483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4646_ _4930_/B _4634_/X _4645_/X vssd1 vssd1 vccd1 vccd1 _4646_/X sky130_fd_sc_hd__a21o_1
X_4577_ _4577_/A vssd1 vssd1 vccd1 vccd1 _8156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _7808_/Q _6286_/X _6315_/X vssd1 vssd1 vccd1 vccd1 _7808_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7296_ _8307_/Q _7295_/X _7286_/X _7178_/B vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6247_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__buf_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7358__123 _7360__125/A vssd1 vssd1 vccd1 vccd1 _8334_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6178_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__buf_2
X_5129_ _8260_/Q _8252_/Q _8244_/Q _8268_/Q _5078_/X _5070_/X vssd1 vssd1 vccd1 vccd1
+ _5129_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7118__84 _7118__84/A vssd1 vssd1 vccd1 vccd1 _8265_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480_ _8001_/Q _4362_/A _5482_/S vssd1 vssd1 vccd1 vccd1 _5481_/A sky130_fd_sc_hd__mux2_1
X_4500_ _4500_/A vssd1 vssd1 vccd1 vccd1 _8190_/D sky130_fd_sc_hd__clkbuf_1
X_4431_ _8449_/Q vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__buf_2
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4362_ _4362_/A vssd1 vssd1 vccd1 vccd1 _4362_/X sky130_fd_sc_hd__clkbuf_2
X_7150_ _8308_/Q _8307_/Q _8306_/Q _8305_/Q vssd1 vssd1 vccd1 vccd1 _7193_/D sky130_fd_sc_hd__and4_1
X_6101_ _6101_/A _6105_/B vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__and2_4
XFILLER_112_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4293_ _4293_/A vssd1 vssd1 vccd1 vccd1 _8269_/D sky130_fd_sc_hd__clkbuf_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _7737_/Q _6044_/B vssd1 vssd1 vccd1 vccd1 _6032_/X sky130_fd_sc_hd__or2_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7983_ _7983_/CLK _7983_/D vssd1 vssd1 vccd1 vccd1 _7983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6865_ _8440_/Q _6963_/C vssd1 vssd1 vccd1 vccd1 _6866_/A sky130_fd_sc_hd__and2_1
X_5816_ _5831_/S vssd1 vssd1 vccd1 vccd1 _5825_/S sky130_fd_sc_hd__buf_2
X_6796_ _6796_/A _6808_/B _6808_/C vssd1 vssd1 vccd1 vccd1 _6797_/B sky130_fd_sc_hd__nand3_1
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3614_ _7368_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3614_/X sky130_fd_sc_hd__clkbuf_16
X_5747_ _7863_/Q _5557_/A _5755_/S vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8466_ _8466_/CLK _8466_/D vssd1 vssd1 vccd1 vccd1 _8466_/Q sky130_fd_sc_hd__dfxtp_1
X_5678_ _5678_/A vssd1 vssd1 vccd1 vccd1 _7894_/D sky130_fd_sc_hd__clkbuf_1
X_7417_ _7417_/A vssd1 vssd1 vccd1 vccd1 _7417_/X sky130_fd_sc_hd__buf_1
X_4629_ _4650_/A vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__clkbuf_4
X_8397_ _8397_/CLK _8397_/D vssd1 vssd1 vccd1 vccd1 _8397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7279_ _7282_/A _7279_/B vssd1 vssd1 vccd1 vccd1 _8301_/D sky130_fd_sc_hd__nor2_1
XFILLER_104_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3227_ clkbuf_0__3227_/X vssd1 vssd1 vccd1 vccd1 _6539__259/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6883__403 _6885__405/A vssd1 vssd1 vccd1 vccd1 _8079_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _4980_/A vssd1 vssd1 vccd1 vccd1 _8103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _8446_/Q vssd1 vssd1 vccd1 vccd1 _3931_/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_1_1_0__3431_ clkbuf_0__3431_/X vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__clkbuf_4
X_3862_ _7854_/Q _7853_/Q vssd1 vssd1 vccd1 vccd1 _6291_/A sky130_fd_sc_hd__or2_1
X_6650_ _7971_/Q _5935_/A _6652_/S vssd1 vssd1 vccd1 vccd1 _6651_/A sky130_fd_sc_hd__mux2_1
X_5601_ _5601_/A _5833_/B vssd1 vssd1 vccd1 vccd1 _5617_/S sky130_fd_sc_hd__or2_4
X_5532_ _5365_/X _7978_/Q _5536_/S vssd1 vssd1 vccd1 vccd1 _5533_/A sky130_fd_sc_hd__mux2_1
X_6931__437 _6932__438/A vssd1 vssd1 vccd1 vccd1 _8115_/CLK sky130_fd_sc_hd__inv_2
X_8320_ _8442_/CLK _8320_/D vssd1 vssd1 vccd1 vccd1 _8320_/Q sky130_fd_sc_hd__dfxtp_1
X_8251_ _8251_/CLK _8251_/D vssd1 vssd1 vccd1 vccd1 _8251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5463_ _5463_/A vssd1 vssd1 vccd1 vccd1 _8009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8182_ _8182_/CLK _8182_/D vssd1 vssd1 vccd1 vccd1 _8182_/Q sky130_fd_sc_hd__dfxtp_1
X_5394_ _5655_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5410_/S sky130_fd_sc_hd__or2_2
X_7202_ _8497_/Q _7273_/A _7273_/B vssd1 vssd1 vccd1 vccd1 _7202_/X sky130_fd_sc_hd__and3_1
X_4414_ _4413_/X _8220_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__mux2_1
X_4345_ _4342_/X _8246_/Q _4357_/S vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7112__79 _7113__80/A vssd1 vssd1 vccd1 vccd1 _8260_/CLK sky130_fd_sc_hd__inv_2
X_4276_ _4276_/A vssd1 vssd1 vccd1 vccd1 _8276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6015_ _6015_/A _6015_/B vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__nor2_2
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _8060_/CLK _7966_/D vssd1 vssd1 vccd1 vccd1 _7966_/Q sky130_fd_sc_hd__dfxtp_1
X_7897_ _7897_/CLK _7897_/D vssd1 vssd1 vccd1 vccd1 _7897_/Q sky130_fd_sc_hd__dfxtp_1
X_6917_ _6917_/A vssd1 vssd1 vccd1 vccd1 _6917_/X sky130_fd_sc_hd__buf_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3629_ clkbuf_0__3629_/X vssd1 vssd1 vccd1 vccd1 _7453__25/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6779_ _7207_/A _7517_/A vssd1 vssd1 vccd1 vccd1 _6779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8449_ _8478_/CLK _8449_/D vssd1 vssd1 vccd1 vccd1 _8449_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_wb_clk_i _6131_/A vssd1 vssd1 vccd1 vccd1 _8439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _8141_/Q _7645_/B vssd1 vssd1 vccd1 vccd1 _4911_/C sky130_fd_sc_hd__and2_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4061_ _4061_/A vssd1 vssd1 vccd1 vccd1 _8374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7820_ _8489_/CLK _7820_/D vssd1 vssd1 vccd1 vccd1 _7820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4963_ _8109_/Q _4235_/X _4965_/S vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__mux2_1
X_7751_ _7964_/CLK _7751_/D vssd1 vssd1 vccd1 vccd1 _7751_/Q sky130_fd_sc_hd__dfxtp_1
X_7033__516 _7034__517/A vssd1 vssd1 vccd1 vccd1 _8197_/CLK sky130_fd_sc_hd__inv_2
X_3914_ _8458_/Q _3892_/X _3914_/S vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7682_ _7680_/Y _7681_/Y _7678_/X vssd1 vssd1 vccd1 vccd1 _8485_/D sky130_fd_sc_hd__a21oi_2
X_4894_ _8105_/Q _4755_/A _4798_/X _4893_/X vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6633_ _6633_/A vssd1 vssd1 vccd1 vccd1 _7963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3414_ clkbuf_0__3414_/X vssd1 vssd1 vccd1 vccd1 _6985__477/A sky130_fd_sc_hd__clkbuf_4
X_3845_ _3845_/A _3845_/B input57/X input58/X vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__or4bb_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3276_ clkbuf_0__3276_/X vssd1 vssd1 vccd1 vccd1 _6688__335/A sky130_fd_sc_hd__clkbuf_4
X_5515_ _5515_/A vssd1 vssd1 vccd1 vccd1 _7986_/D sky130_fd_sc_hd__clkbuf_1
X_8303_ _8309_/CLK _8303_/D vssd1 vssd1 vccd1 vccd1 _8303_/Q sky130_fd_sc_hd__dfxtp_1
X_8234_ _8234_/CLK _8234_/D vssd1 vssd1 vccd1 vccd1 _8234_/Q sky130_fd_sc_hd__dfxtp_1
X_5446_ _8019_/Q _4454_/X _5446_/S vssd1 vssd1 vccd1 vccd1 _5447_/A sky130_fd_sc_hd__mux2_1
X_6270__204 _6271__205/A vssd1 vssd1 vccd1 vccd1 _7796_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3630_ clkbuf_0__3630_/X vssd1 vssd1 vccd1 vccd1 _7633_/A sky130_fd_sc_hd__clkbuf_4
X_5377_ _5392_/S vssd1 vssd1 vccd1 vccd1 _5386_/S sky130_fd_sc_hd__clkbuf_4
X_8165_ _8165_/CLK _8165_/D vssd1 vssd1 vccd1 vccd1 _8165_/Q sky130_fd_sc_hd__dfxtp_1
X_4328_ _8253_/Q _4182_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__mux2_1
X_7097__67 _7098__68/A vssd1 vssd1 vccd1 vccd1 _8248_/CLK sky130_fd_sc_hd__inv_2
X_8096_ _8096_/CLK _8096_/D vssd1 vssd1 vccd1 vccd1 _8096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4259_ _8283_/Q _4188_/X _4261_/S vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7949_ _7949_/CLK _7949_/D vssd1 vssd1 vccd1 vccd1 _7949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__3061_ clkbuf_0__3061_/X vssd1 vssd1 vccd1 vccd1 _6271__205/A sky130_fd_sc_hd__clkbuf_4
X_5300_ _5295_/A _5298_/X _5299_/X vssd1 vssd1 vccd1 vccd1 _5300_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5231_ _5083_/X _5218_/X _5222_/X _5230_/X _5332_/B vssd1 vssd1 vccd1 vccd1 _5231_/X
+ sky130_fd_sc_hd__o311a_1
X_5162_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__inv_2
X_5093_ _8363_/Q _8347_/Q _8339_/Q _8371_/Q _5060_/X _5044_/X vssd1 vssd1 vccd1 vccd1
+ _5093_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4113_ _8128_/Q _4113_/B vssd1 vssd1 vccd1 vccd1 _4113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4044_/A vssd1 vssd1 vccd1 vccd1 _8381_/D sky130_fd_sc_hd__clkbuf_1
X_7352__118 _7354__120/A vssd1 vssd1 vccd1 vccd1 _8329_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7803_ _7803_/CLK _7803_/D vssd1 vssd1 vccd1 vccd1 _7803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5995_ _7967_/Q _6006_/B vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__and2_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7734_ _8308_/CLK _7734_/D vssd1 vssd1 vccd1 vccd1 _7734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4946_ _8116_/Q _4238_/X _4946_/S vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _4770_/A _7992_/Q _7928_/Q _4769_/A vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__a22o_1
X_7665_ _8480_/Q _7656_/X _7664_/X _7662_/X vssd1 vssd1 vccd1 vccd1 _8480_/D sky130_fd_sc_hd__o211a_1
X_6616_ _5902_/A _7956_/Q _6616_/S vssd1 vssd1 vccd1 vccd1 _6617_/A sky130_fd_sc_hd__mux2_1
X_7596_ _7510_/A _7578_/A _7595_/X _7582_/A vssd1 vssd1 vccd1 vccd1 _8441_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3828_ _8075_/Q _8074_/Q _8073_/Q vssd1 vssd1 vccd1 vccd1 _5316_/A sky130_fd_sc_hd__and3_1
X_6547_ _6547_/A vssd1 vssd1 vccd1 vccd1 _6547_/X sky130_fd_sc_hd__buf_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6478_ _6478_/A vssd1 vssd1 vccd1 vccd1 _7853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5429_ _5429_/A vssd1 vssd1 vccd1 vccd1 _8027_/D sky130_fd_sc_hd__clkbuf_1
X_8217_ _8217_/CLK _8217_/D vssd1 vssd1 vccd1 vccd1 _8217_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3227_ _6535_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3227_/X sky130_fd_sc_hd__clkbuf_16
X_8148_ _8148_/CLK _8148_/D vssd1 vssd1 vccd1 vccd1 _8148_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3613_ clkbuf_0__3613_/X vssd1 vssd1 vccd1 vccd1 _7367__130/A sky130_fd_sc_hd__clkbuf_4
X_6944__447 _6944__447/A vssd1 vssd1 vccd1 vccd1 _8126_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_1 _7775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8079_ _8079_/CLK _8079_/D vssd1 vssd1 vccd1 vccd1 _8079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4932_/B _4797_/X _4799_/X vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5780_ _5795_/S vssd1 vssd1 vccd1 vccd1 _5789_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _8093_/Q _7980_/Q _7884_/Q _7860_/Q _4630_/A _4633_/A vssd1 vssd1 vccd1 vccd1
+ _4731_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__clkbuf_2
X_6401_ _6401_/A vssd1 vssd1 vccd1 vccd1 _6401_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _8149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6332_ _7200_/A _6293_/A _6299_/X vssd1 vssd1 vccd1 vccd1 _6332_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__clkbuf_2
X_8002_ _8002_/CLK _8002_/D vssd1 vssd1 vccd1 vccd1 _8002_/Q sky130_fd_sc_hd__dfxtp_1
X_6194_ _7678_/A vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__buf_4
XFILLER_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5145_ _8462_/Q _8023_/Q _7988_/Q _8454_/Q _5291_/S _5111_/X vssd1 vssd1 vccd1 vccd1
+ _5145_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5076_ _8174_/Q _8150_/Q _8412_/Q _8182_/Q _5123_/A _5044_/A vssd1 vssd1 vccd1 vccd1
+ _5076_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _5797_/B _5430_/B vssd1 vssd1 vccd1 vccd1 _4043_/S sky130_fd_sc_hd__nor2_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _7959_/Q _5982_/B vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__and2_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7717_ _7717_/A vssd1 vssd1 vccd1 vccd1 _8497_/D sky130_fd_sc_hd__clkbuf_1
X_4929_ _4653_/A _4924_/X _4928_/Y _4841_/X vssd1 vssd1 vccd1 vccd1 _8125_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7648_ _7649_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _8476_/D sky130_fd_sc_hd__nor2_1
X_6950__451 _6952__453/A vssd1 vssd1 vccd1 vccd1 _8130_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7579_ _8434_/Q _7584_/B vssd1 vssd1 vccd1 vccd1 _7579_/X sky130_fd_sc_hd__or2_1
X_7144__105 _7144__105/A vssd1 vssd1 vccd1 vccd1 _8286_/CLK sky130_fd_sc_hd__inv_2
X_7046__526 _7048__528/A vssd1 vssd1 vccd1 vccd1 _8207_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_108 _8490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3389_ clkbuf_0__3389_/X vssd1 vssd1 vccd1 vccd1 _6878__400/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5901_ _5901_/A vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _5832_/A vssd1 vssd1 vccd1 vccd1 _7776_/D sky130_fd_sc_hd__clkbuf_1
X_5763_ _4101_/X _7807_/Q _5769_/S vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3630_ _7454_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3630_/X sky130_fd_sc_hd__clkbuf_16
X_4714_ _4735_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4714_/X sky130_fd_sc_hd__and2_1
X_7502_ _8413_/Q _7508_/A vssd1 vssd1 vccd1 vccd1 _7577_/A sky130_fd_sc_hd__or2b_1
X_5694_ _5694_/A vssd1 vssd1 vccd1 vccd1 _7887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8482_ _8483_/CLK _8482_/D vssd1 vssd1 vccd1 vccd1 _8482_/Q sky130_fd_sc_hd__dfxtp_2
X_4645_ _4637_/X _4641_/X _4644_/X vssd1 vssd1 vccd1 vccd1 _4645_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4576_ _4413_/X _8156_/Q _4580_/S vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6315_ _6289_/X _6300_/X _6314_/X _6192_/X vssd1 vssd1 vccd1 vccd1 _6315_/X sky130_fd_sc_hd__a31o_1
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7295_ _7295_/A vssd1 vssd1 vccd1 vccd1 _7295_/X sky130_fd_sc_hd__clkbuf_2
X_6828__373 _6830__375/A vssd1 vssd1 vccd1 vccd1 _8041_/CLK sky130_fd_sc_hd__inv_2
X_6177_ _6176_/X _7957_/Q _6170_/X _6172_/X _7746_/Q vssd1 vssd1 vccd1 vccd1 _7746_/D
+ sky130_fd_sc_hd__o32a_1
X_5128_ _8378_/Q _8276_/Q _8013_/Q _8228_/Q _5111_/A _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5128_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__buf_2
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6577__290 _6577__290/A vssd1 vssd1 vccd1 vccd1 _7930_/CLK sky130_fd_sc_hd__inv_2
X_7365__128 _7366__129/A vssd1 vssd1 vccd1 vccd1 _8339_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6248__186 _6249__187/A vssd1 vssd1 vccd1 vccd1 _7778_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6957__457 _6957__457/A vssd1 vssd1 vccd1 vccd1 _8136_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4430_ _4430_/A vssd1 vssd1 vccd1 vccd1 _8215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4361_ _4361_/A vssd1 vssd1 vccd1 vccd1 _8241_/D sky130_fd_sc_hd__clkbuf_1
X_6100_ _7754_/Q _6095_/X _6096_/X _6099_/X _6093_/X vssd1 vssd1 vccd1 vccd1 _6100_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4292_ _3925_/X _8269_/Q _4298_/S vssd1 vssd1 vccd1 vccd1 _4293_/A sky130_fd_sc_hd__mux2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _7812_/Q input29/X _6039_/S vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7982_ _7982_/CLK _7982_/D vssd1 vssd1 vccd1 vccd1 _7982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6864_ _6864_/A vssd1 vssd1 vccd1 vccd1 _8065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5815_ _5815_/A _5815_/B vssd1 vssd1 vccd1 vccd1 _5831_/S sky130_fd_sc_hd__nor2_2
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6795_ _8424_/Q _8423_/Q vssd1 vssd1 vccd1 vccd1 _6796_/A sky130_fd_sc_hd__and2_1
Xclkbuf_0__3613_ _7362_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3613_/X sky130_fd_sc_hd__clkbuf_16
X_5746_ _5761_/S vssd1 vssd1 vccd1 vccd1 _5755_/S sky130_fd_sc_hd__buf_2
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5677_ _7894_/Q _4978_/X _5683_/S vssd1 vssd1 vccd1 vccd1 _5678_/A sky130_fd_sc_hd__mux2_1
X_8465_ _8465_/CLK _8465_/D vssd1 vssd1 vccd1 vccd1 _8465_/Q sky130_fd_sc_hd__dfxtp_1
X_4628_ _8122_/Q vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8396_ _8396_/CLK _8396_/D vssd1 vssd1 vccd1 vccd1 _8396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4559_ _4416_/X _8163_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7278_ _7211_/B _7264_/X _7272_/X _7197_/B vssd1 vssd1 vccd1 vccd1 _7279_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6229_ _6232_/B _6229_/B _6231_/C vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__and3_1
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3226_ clkbuf_0__3226_/X vssd1 vssd1 vccd1 vccd1 _6531__252/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _3930_/A vssd1 vssd1 vccd1 vccd1 _8455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _7832_/Q _6304_/C vssd1 vssd1 vccd1 vccd1 _7659_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5600_ _5600_/A vssd1 vssd1 vccd1 vccd1 _7928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5531_ _5531_/A vssd1 vssd1 vccd1 vccd1 _7979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8250_ _8250_/CLK _8250_/D vssd1 vssd1 vccd1 vccd1 _8250_/Q sky130_fd_sc_hd__dfxtp_1
X_5462_ _8009_/Q _4451_/X _5464_/S vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__mux2_1
X_7201_ _8298_/Q _8297_/Q _8299_/Q vssd1 vssd1 vccd1 vccd1 _7273_/B sky130_fd_sc_hd__a21o_1
X_8181_ _8181_/CLK _8181_/D vssd1 vssd1 vccd1 vccd1 _8181_/Q sky130_fd_sc_hd__dfxtp_1
X_5393_ _5393_/A vssd1 vssd1 vccd1 vccd1 _8044_/D sky130_fd_sc_hd__clkbuf_1
X_4413_ _8065_/Q vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__clkbuf_2
X_4344_ _4366_/S vssd1 vssd1 vccd1 vccd1 _4357_/S sky130_fd_sc_hd__buf_2
X_7132_ _7132_/A vssd1 vssd1 vccd1 vccd1 _7132_/X sky130_fd_sc_hd__buf_1
XFILLER_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7063_/X sky130_fd_sc_hd__buf_1
X_4275_ _8276_/Q _4185_/X _4279_/S vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _7733_/Q _6025_/B vssd1 vssd1 vccd1 vccd1 _6014_/X sky130_fd_sc_hd__or2_1
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8500__250 vssd1 vssd1 vccd1 vccd1 core1Index[0] _8500__250/LO sky130_fd_sc_hd__conb_1
X_7965_ _8060_/CLK _7965_/D vssd1 vssd1 vccd1 vccd1 _7965_/Q sky130_fd_sc_hd__dfxtp_1
X_7896_ _7896_/CLK _7896_/D vssd1 vssd1 vccd1 vccd1 _7896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6916_ _7044_/A vssd1 vssd1 vccd1 vccd1 _6916_/X sky130_fd_sc_hd__buf_1
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6778_ _8415_/Q vssd1 vssd1 vccd1 vccd1 _7517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5729_ _7871_/Q _5557_/A _5737_/S vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8448_ _8478_/CLK _8448_/D vssd1 vssd1 vccd1 vccd1 _8448_/Q sky130_fd_sc_hd__dfxtp_2
X_8379_ _8379_/CLK _8379_/D vssd1 vssd1 vccd1 vccd1 _8379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3389_ _6873_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3389_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4060_ _8374_/Q _4018_/X _4062_/S vssd1 vssd1 vccd1 vccd1 _4061_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4962_ _4962_/A vssd1 vssd1 vccd1 vccd1 _8110_/D sky130_fd_sc_hd__clkbuf_1
X_7750_ _7964_/CLK _7750_/D vssd1 vssd1 vccd1 vccd1 _7750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6701_ _6701_/A vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__buf_1
X_4893_ _8044_/Q _4814_/A _4776_/A _4892_/X vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__o22a_1
X_3913_ _3913_/A vssd1 vssd1 vccd1 vccd1 _8459_/D sky130_fd_sc_hd__clkbuf_1
X_7681_ _7681_/A _7693_/B vssd1 vssd1 vccd1 vccd1 _7681_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__3413_ clkbuf_0__3413_/X vssd1 vssd1 vccd1 vccd1 _6989_/A sky130_fd_sc_hd__clkbuf_4
X_3844_ _3844_/A _3844_/B input69/X vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__or3b_1
X_6632_ _5917_/A _7963_/Q _6634_/S vssd1 vssd1 vccd1 vccd1 _6633_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6682__330/A sky130_fd_sc_hd__clkbuf_4
X_5514_ _7986_/Q _4359_/A _5518_/S vssd1 vssd1 vccd1 vccd1 _5515_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8302_ _8309_/CLK _8302_/D vssd1 vssd1 vccd1 vccd1 _8302_/Q sky130_fd_sc_hd__dfxtp_1
X_8233_ _8233_/CLK _8233_/D vssd1 vssd1 vccd1 vccd1 _8233_/Q sky130_fd_sc_hd__dfxtp_1
X_5445_ _5445_/A vssd1 vssd1 vccd1 vccd1 _8020_/D sky130_fd_sc_hd__clkbuf_1
X_8164_ _8164_/CLK _8164_/D vssd1 vssd1 vccd1 vccd1 _8164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5376_ _5601_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5392_/S sky130_fd_sc_hd__or2_2
X_4327_ _4327_/A vssd1 vssd1 vccd1 vccd1 _8254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8095_ _8095_/CLK _8095_/D vssd1 vssd1 vccd1 vccd1 _8095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4258_ _4258_/A vssd1 vssd1 vccd1 vccd1 _8284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4189_ _8337_/Q _4188_/X _4192_/S vssd1 vssd1 vccd1 vccd1 _4190_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7948_ _7948_/CLK _7948_/D vssd1 vssd1 vccd1 vccd1 _7948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7879_ _7879_/CLK _7879_/D vssd1 vssd1 vccd1 vccd1 _7879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3758_ clkbuf_0__3758_/X vssd1 vssd1 vccd1 vccd1 _7644__50/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3421_ clkbuf_0__3421_/X vssd1 vssd1 vccd1 vccd1 _7024__509/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3060_ clkbuf_0__3060_/X vssd1 vssd1 vccd1 vccd1 _6278_/A sky130_fd_sc_hd__clkbuf_4
X_5230_ _5224_/X _5225_/X _5334_/B _5229_/X vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__a211o_1
XFILLER_6_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5161_ _8070_/Q vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _3916_/X _5022_/X _5089_/X _5091_/X vssd1 vssd1 vccd1 vccd1 _8086_/D sky130_fd_sc_hd__o211a_1
X_4112_ _8129_/Q _8124_/Q vssd1 vssd1 vccd1 vccd1 _4113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4043_ _8381_/Q _4022_/X _4043_/S vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822__368 _6824__370/A vssd1 vssd1 vccd1 vccd1 _8036_/CLK sky130_fd_sc_hd__inv_2
X_5994_ _5994_/A vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__clkbuf_1
X_7802_ _7802_/CLK _7802_/D vssd1 vssd1 vccd1 vccd1 _7802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7733_ _8308_/CLK _7733_/D vssd1 vssd1 vccd1 vccd1 _7733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ _4945_/A vssd1 vssd1 vccd1 vccd1 _8117_/D sky130_fd_sc_hd__clkbuf_1
X_4876_ _4871_/X _4872_/X _4875_/X _4928_/B vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__a211o_1
X_7664_ _5917_/A _7657_/X _7660_/Y vssd1 vssd1 vccd1 vccd1 _7664_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3827_ _3815_/A _5054_/A _3826_/Y vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__a21bo_1
X_6615_ _6615_/A vssd1 vssd1 vccd1 vccd1 _7955_/D sky130_fd_sc_hd__clkbuf_1
X_7595_ _8441_/Q _7595_/B vssd1 vssd1 vccd1 vccd1 _7595_/X sky130_fd_sc_hd__or2_1
XFILLER_118_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6571__285 _6571__285/A vssd1 vssd1 vccd1 vccd1 _7925_/CLK sky130_fd_sc_hd__inv_2
X_6477_ _7662_/A _6477_/B _6480_/B vssd1 vssd1 vccd1 vccd1 _6478_/A sky130_fd_sc_hd__and3_1
X_5428_ _3892_/X _8027_/Q _5428_/S vssd1 vssd1 vccd1 vccd1 _5429_/A sky130_fd_sc_hd__mux2_1
X_8216_ _8216_/CLK _8216_/D vssd1 vssd1 vccd1 vccd1 _8216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8147_ _8147_/CLK _8147_/D vssd1 vssd1 vccd1 vccd1 _8147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3226_ _6529_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3226_/X sky130_fd_sc_hd__clkbuf_16
X_5359_ _5359_/A vssd1 vssd1 vccd1 vccd1 _8056_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3612_ clkbuf_0__3612_/X vssd1 vssd1 vccd1 vccd1 _7386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_2 _7775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _8078_/CLK _8078_/D vssd1 vssd1 vccd1 vccd1 _8078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7632__40 _7632__40/A vssd1 vssd1 vccd1 vccd1 _8463_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _8048_/Q _8040_/Q _7868_/Q _8109_/Q _4648_/X _4640_/X vssd1 vssd1 vccd1 vccd1
+ _4730_/X sky130_fd_sc_hd__mux4_1
X_4661_ _4661_/A _4661_/B vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__and2_1
XFILLER_119_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7380_ _7380_/A vssd1 vssd1 vccd1 vccd1 _7380_/X sky130_fd_sc_hd__buf_1
X_6400_ _7823_/Q _6383_/X _6393_/X _6399_/X _6391_/X vssd1 vssd1 vccd1 vccd1 _7823_/D
+ sky130_fd_sc_hd__a221o_1
X_4592_ _8149_/Q _4436_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__mux2_1
X_6331_ _8496_/Q vssd1 vssd1 vccd1 vccd1 _7200_/A sky130_fd_sc_hd__buf_4
X_5213_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__buf_2
X_8001_ _8001_/CLK _8001_/D vssd1 vssd1 vccd1 vccd1 _8001_/Q sky130_fd_sc_hd__dfxtp_1
X_6193_ _6192_/X _7967_/Q _6186_/X _6188_/X _7756_/Q vssd1 vssd1 vccd1 vccd1 _7756_/D
+ sky130_fd_sc_hd__o32a_1
X_5144_ _7796_/Q _8004_/Q _8283_/Q _8031_/Q _5241_/S _5052_/X vssd1 vssd1 vccd1 vccd1
+ _5144_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5075_ _5190_/S vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__buf_2
XFILLER_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7004__493 _7004__493/A vssd1 vssd1 vccd1 vccd1 _8174_/CLK sky130_fd_sc_hd__inv_2
X_4026_ _5466_/A vssd1 vssd1 vccd1 vccd1 _5430_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ _5977_/A vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7716_ _7722_/A _7716_/B vssd1 vssd1 vccd1 vccd1 _7717_/A sky130_fd_sc_hd__or2_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4928_ _4932_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7647_ _7647_/A vssd1 vssd1 vccd1 vccd1 _8475_/D sky130_fd_sc_hd__clkbuf_1
X_4859_ _8350_/Q _4619_/A _4803_/X _8326_/Q _4798_/X vssd1 vssd1 vccd1 vccd1 _4859_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7578_ _7578_/A vssd1 vssd1 vccd1 vccd1 _7578_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6529_ _6553_/A vssd1 vssd1 vccd1 vccd1 _6529_/X sky130_fd_sc_hd__buf_1
XFILLER_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8543__242 vssd1 vssd1 vccd1 vccd1 _8543__242/HI partID[7] sky130_fd_sc_hd__conb_1
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6283__215 _6283__215/A vssd1 vssd1 vccd1 vccd1 _7807_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_109 _6228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7422__175 _7422__175/A vssd1 vssd1 vccd1 vccd1 _8386_/CLK sky130_fd_sc_hd__inv_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _7690_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__or2_1
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6880_ _6886_/A vssd1 vssd1 vccd1 vccd1 _6880_/X sky130_fd_sc_hd__buf_1
X_5831_ _7776_/Q _5580_/A _5831_/S vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _5762_/A vssd1 vssd1 vccd1 vccd1 _7856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4713_ _7781_/Q _7901_/Q _7909_/Q _7949_/Q _4630_/A _4633_/A vssd1 vssd1 vccd1 vccd1
+ _4714_/B sky130_fd_sc_hd__mux4_1
X_7501_ _7491_/X _7490_/A _7577_/B _7572_/C vssd1 vssd1 vccd1 vccd1 _7544_/A sky130_fd_sc_hd__a22oi_4
X_5693_ _7887_/Q _4973_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__mux2_1
X_8481_ _8481_/CLK _8481_/D vssd1 vssd1 vccd1 vccd1 _8481_/Q sky130_fd_sc_hd__dfxtp_1
X_4644_ _4665_/A vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__clkbuf_2
X_4575_ _4575_/A vssd1 vssd1 vccd1 vccd1 _8157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7294_ _7297_/A _7294_/B vssd1 vssd1 vccd1 vccd1 _8306_/D sky130_fd_sc_hd__nor2_1
X_6314_ _6306_/X _6309_/X _6311_/X _8121_/Q _6393_/A vssd1 vssd1 vccd1 vccd1 _6314_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8527__226 vssd1 vssd1 vccd1 vccd1 _8527__226/HI core1Index[6] sky130_fd_sc_hd__conb_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6176_ _7678_/A vssd1 vssd1 vccd1 vccd1 _6176_/X sky130_fd_sc_hd__buf_2
X_5127_ _5099_/X _5124_/X _5126_/X vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5058_ _5038_/X _5045_/X _5057_/X vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__a21o_1
X_4009_ _8445_/Q vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7052__531 _7054__533/A vssd1 vssd1 vccd1 vccd1 _8212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3758_ _7639_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3758_/X sky130_fd_sc_hd__clkbuf_16
X_6835__378 _6836__379/A vssd1 vssd1 vccd1 vccd1 _8046_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6731__365 _6731__365/A vssd1 vssd1 vccd1 vccd1 _8032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4360_ _4359_/X _8241_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7124__89 _7125__90/A vssd1 vssd1 vccd1 vccd1 _8270_/CLK sky130_fd_sc_hd__inv_2
X_4291_ _4291_/A vssd1 vssd1 vccd1 vccd1 _8270_/D sky130_fd_sc_hd__clkbuf_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6030_ _6009_/X _6027_/X _6029_/X _6018_/X vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__o211a_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7981_ _7981_/CLK _7981_/D vssd1 vssd1 vccd1 vccd1 _7981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6863_ _8439_/Q _6863_/B vssd1 vssd1 vccd1 vccd1 _6864_/A sky130_fd_sc_hd__and2_1
X_5814_ _5814_/A vssd1 vssd1 vccd1 vccd1 _7784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6794_ _6794_/A _6794_/B _6794_/C _6794_/D vssd1 vssd1 vccd1 vccd1 _6794_/X sky130_fd_sc_hd__and4_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3612_ _7361_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3612_/X sky130_fd_sc_hd__clkbuf_16
X_5745_ _5745_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5761_/S sky130_fd_sc_hd__nor2_2
XFILLER_108_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5676_ _5676_/A vssd1 vssd1 vccd1 vccd1 _7895_/D sky130_fd_sc_hd__clkbuf_1
X_8464_ _8464_/CLK _8464_/D vssd1 vssd1 vccd1 vccd1 _8464_/Q sky130_fd_sc_hd__dfxtp_1
X_4627_ _4627_/A vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__buf_2
X_8395_ _8395_/CLK _8395_/D vssd1 vssd1 vccd1 vccd1 _8395_/Q sky130_fd_sc_hd__dfxtp_1
X_7346_ _7346_/A vssd1 vssd1 vccd1 vccd1 _8324_/D sky130_fd_sc_hd__clkbuf_1
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _8164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _8193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7277_ _7282_/A _7277_/B vssd1 vssd1 vccd1 vccd1 _8300_/D sky130_fd_sc_hd__nor2_1
X_6228_ _7774_/Q _7773_/Q _6228_/C vssd1 vssd1 vccd1 vccd1 _6231_/C sky130_fd_sc_hd__or3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _7678_/A vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7371__133 _7373__135/A vssd1 vssd1 vccd1 vccd1 _8344_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3225_ clkbuf_0__3225_/X vssd1 vssd1 vccd1 vccd1 _6553_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6254__191 _6254__191/A vssd1 vssd1 vccd1 vccd1 _7783_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7059__537 _7059__537/A vssd1 vssd1 vccd1 vccd1 _8218_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6890__409 _6891__410/A vssd1 vssd1 vccd1 vccd1 _8085_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _7652_/A _7652_/B _7652_/C _7652_/D vssd1 vssd1 vccd1 vccd1 _6304_/C sky130_fd_sc_hd__or4_2
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _5361_/X _7979_/Q _5530_/S vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5461_ _5461_/A vssd1 vssd1 vccd1 vccd1 _8010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7200_ _7200_/A _7200_/B vssd1 vssd1 vccd1 vccd1 _7200_/X sky130_fd_sc_hd__xor2_1
X_4412_ _4412_/A vssd1 vssd1 vccd1 vccd1 _8221_/D sky130_fd_sc_hd__clkbuf_1
X_8180_ _8180_/CLK _8180_/D vssd1 vssd1 vccd1 vccd1 _8180_/Q sky130_fd_sc_hd__dfxtp_1
X_5392_ _5373_/X _8044_/Q _5392_/S vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__mux2_1
X_4343_ _5797_/A _4343_/B vssd1 vssd1 vccd1 vccd1 _4366_/S sky130_fd_sc_hd__or2_4
X_4274_ _4274_/A vssd1 vssd1 vccd1 vccd1 _8277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6013_ _6085_/A vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__buf_4
XFILLER_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6899__412 _6900__413/A vssd1 vssd1 vccd1 vccd1 _8090_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7964_ _7964_/CLK _7964_/D vssd1 vssd1 vccd1 vccd1 _7964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6915_/A vssd1 vssd1 vccd1 vccd1 _6915_/X sky130_fd_sc_hd__buf_1
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7895_ _7895_/CLK _7895_/D vssd1 vssd1 vccd1 vccd1 _7895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3627_ clkbuf_0__3627_/X vssd1 vssd1 vccd1 vccd1 _7441__15/A sky130_fd_sc_hd__clkbuf_4
X_6777_ _6782_/C _6777_/B vssd1 vssd1 vccd1 vccd1 _6777_/Y sky130_fd_sc_hd__xnor2_1
X_5728_ _5743_/S vssd1 vssd1 vccd1 vccd1 _5737_/S sky130_fd_sc_hd__clkbuf_4
X_3989_ _3943_/X _8397_/Q _3989_/S vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5659_ _5562_/X _7902_/Q _5665_/S vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8447_ _8447_/CLK _8447_/D vssd1 vssd1 vccd1 vccd1 _8447_/Q sky130_fd_sc_hd__dfxtp_2
X_8378_ _8378_/CLK _8378_/D vssd1 vssd1 vccd1 vccd1 _8378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7329_ _8079_/Q _7648_/B _7326_/X _7328_/X _7248_/X vssd1 vssd1 vccd1 vccd1 _8316_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6696__341 _6698__343/A vssd1 vssd1 vccd1 vccd1 _8005_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7378__139 _7379__140/A vssd1 vssd1 vccd1 vccd1 _8350_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i _8447_/CLK vssd1 vssd1 vccd1 vccd1 _8481_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4961_ _8110_/Q _4232_/X _4965_/S vssd1 vssd1 vccd1 vccd1 _4962_/A sky130_fd_sc_hd__mux2_1
X_4892_ _4770_/A _8036_/Q _7864_/Q _4769_/A vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__a22o_1
X_3912_ _8459_/Q _3889_/X _3914_/S vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__mux2_1
X_7680_ _7680_/A _7692_/B vssd1 vssd1 vccd1 vccd1 _7680_/Y sky130_fd_sc_hd__nand2_1
X_3843_ _3843_/A _3843_/B _3843_/C vssd1 vssd1 vccd1 vccd1 _6015_/A sky130_fd_sc_hd__or3_2
X_6631_ _6631_/A vssd1 vssd1 vccd1 vccd1 _7962_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3412_ clkbuf_0__3412_/X vssd1 vssd1 vccd1 vccd1 _6981__475/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8301_ _8315_/CLK _8301_/D vssd1 vssd1 vccd1 vccd1 _8301_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6683_/A sky130_fd_sc_hd__clkbuf_4
X_5513_ _5513_/A vssd1 vssd1 vccd1 vccd1 _7987_/D sky130_fd_sc_hd__clkbuf_1
X_8232_ _8232_/CLK _8232_/D vssd1 vssd1 vccd1 vccd1 _8232_/Q sky130_fd_sc_hd__dfxtp_1
X_5444_ _8020_/Q _4451_/X _5446_/S vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8163_ _8163_/CLK _8163_/D vssd1 vssd1 vccd1 vccd1 _8163_/Q sky130_fd_sc_hd__dfxtp_1
X_7114_ _7120_/A vssd1 vssd1 vccd1 vccd1 _7114_/X sky130_fd_sc_hd__buf_1
X_5375_ _5375_/A vssd1 vssd1 vccd1 vccd1 _8052_/D sky130_fd_sc_hd__clkbuf_1
X_4326_ _8254_/Q _4177_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8094_ _8094_/CLK _8094_/D vssd1 vssd1 vccd1 vccd1 _8094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _8284_/Q _4185_/X _4261_/S vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7045_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7045_/X sky130_fd_sc_hd__buf_1
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4188_ _8446_/Q vssd1 vssd1 vccd1 vccd1 _4188_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7947_ _7947_/CLK _7947_/D vssd1 vssd1 vccd1 vccd1 _7947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _7878_/CLK _7878_/D vssd1 vssd1 vccd1 vccd1 _7878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3757_ clkbuf_0__3757_/X vssd1 vssd1 vccd1 vccd1 _7638__45/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8507__257 vssd1 vssd1 vccd1 vccd1 partID[11] _8507__257/LO sky130_fd_sc_hd__conb_1
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3420_ clkbuf_0__3420_/X vssd1 vssd1 vccd1 vccd1 _7019__505/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _5160_/A vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__buf_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4111_ _8127_/Q _4127_/A vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__and2_1
X_5091_ _7598_/A vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4042_ _4042_/A vssd1 vssd1 vccd1 vccd1 _8382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7801_ _7801_/CLK _7801_/D vssd1 vssd1 vccd1 vccd1 _7801_/Q sky130_fd_sc_hd__dfxtp_1
X_5993_ _7966_/Q _5993_/B vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__and2_2
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7732_ _7732_/CLK _7732_/D vssd1 vssd1 vccd1 vccd1 _7732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4944_ _8117_/Q _4235_/X _4946_/S vssd1 vssd1 vccd1 vccd1 _4945_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _7944_/Q _4755_/A _4661_/A _4874_/X vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__o211a_1
X_7663_ _8479_/Q _7656_/X _7661_/X _7662_/X vssd1 vssd1 vccd1 vccd1 _8479_/D sky130_fd_sc_hd__o211a_1
X_3826_ _8077_/Q _8072_/Q vssd1 vssd1 vccd1 vccd1 _3826_/Y sky130_fd_sc_hd__xnor2_1
X_6614_ _7690_/A _7955_/Q _6616_/S vssd1 vssd1 vccd1 vccd1 _6615_/A sky130_fd_sc_hd__mux2_1
X_7594_ _8441_/Q _7578_/A _7593_/X _7582_/A vssd1 vssd1 vccd1 vccd1 _8440_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8215_ _8215_/CLK _8215_/D vssd1 vssd1 vccd1 vccd1 _8215_/Q sky130_fd_sc_hd__dfxtp_1
X_6476_ _6423_/A _7703_/A _6129_/C _6292_/B vssd1 vssd1 vccd1 vccd1 _6480_/B sky130_fd_sc_hd__a31o_1
X_5427_ _5427_/A vssd1 vssd1 vccd1 vccd1 _8028_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3225_ _6528_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3225_/X sky130_fd_sc_hd__clkbuf_16
X_5358_ _5357_/X _8056_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__mux2_1
X_8146_ _8146_/CLK _8146_/D vssd1 vssd1 vccd1 vccd1 _8146_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3611_ clkbuf_0__3611_/X vssd1 vssd1 vccd1 vccd1 _7360__125/A sky130_fd_sc_hd__clkbuf_4
X_4309_ _4309_/A vssd1 vssd1 vccd1 vccd1 _8262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_3 _7775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8077_ _8077_/CLK _8077_/D vssd1 vssd1 vccd1 vccd1 _8077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5289_ _5174_/X _5287_/X _5288_/X vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7016__502 _7019__505/A vssd1 vssd1 vccd1 vccd1 _8183_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6548__266 _6549__267/A vssd1 vssd1 vccd1 vccd1 _7906_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4660_ _7783_/Q _7903_/Q _7911_/Q _7951_/Q _4630_/A _4633_/A vssd1 vssd1 vccd1 vccd1
+ _4661_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4591_ _4591_/A vssd1 vssd1 vccd1 vccd1 _8150_/D sky130_fd_sc_hd__clkbuf_1
X_6330_ _7810_/Q _6286_/X _6329_/X vssd1 vssd1 vccd1 vccd1 _7810_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8000_ _8000_/CLK _8000_/D vssd1 vssd1 vccd1 vccd1 _8000_/Q sky130_fd_sc_hd__dfxtp_1
X_5212_ _8241_/Q _8249_/Q _5235_/S vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__mux2_1
X_6192_ _6328_/A vssd1 vssd1 vccd1 vccd1 _6192_/X sky130_fd_sc_hd__buf_2
X_5143_ _5038_/X _5140_/X _5142_/X vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5074_ _5098_/A vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__buf_4
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _5328_/A _4025_/B _3948_/A _3949_/A vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__or4bb_4
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5976_ _5976_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5977_/A sky130_fd_sc_hd__and2_1
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7715_ _6774_/A _7604_/C _7721_/S vssd1 vssd1 vccd1 vccd1 _7716_/B sky130_fd_sc_hd__mux2_1
X_4927_ _8126_/Q _4924_/X _4926_/Y _4841_/X vssd1 vssd1 vccd1 vccd1 _8126_/D sky130_fd_sc_hd__o211a_1
X_4858_ _8216_/Q _4795_/X _4796_/X _7873_/Q vssd1 vssd1 vccd1 vccd1 _4858_/X sky130_fd_sc_hd__a22o_1
X_7646_ _8132_/Q _7662_/A vssd1 vssd1 vccd1 vccd1 _7647_/A sky130_fd_sc_hd__and2_1
X_4789_ _4789_/A vssd1 vssd1 vccd1 vccd1 _4789_/X sky130_fd_sc_hd__clkbuf_2
X_7577_ _7577_/A _7577_/B vssd1 vssd1 vccd1 vccd1 _7578_/A sky130_fd_sc_hd__or2_1
X_6528_ _6559_/A vssd1 vssd1 vccd1 vccd1 _6528_/X sky130_fd_sc_hd__buf_1
XFILLER_106_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6459_ _6459_/A vssd1 vssd1 vccd1 vccd1 _7846_/D sky130_fd_sc_hd__clkbuf_1
X_8129_ _8129_/CLK _8129_/D vssd1 vssd1 vccd1 vccd1 _8129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6589__300 _6589__300/A vssd1 vssd1 vccd1 vccd1 _7940_/CLK sky130_fd_sc_hd__inv_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _5830_/A vssd1 vssd1 vccd1 vccd1 _7777_/D sky130_fd_sc_hd__clkbuf_1
X_6596__304 _6597__305/A vssd1 vssd1 vccd1 vccd1 _7944_/CLK sky130_fd_sc_hd__inv_2
X_5761_ _7856_/Q _5580_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__mux2_1
X_4712_ _4627_/A _4709_/X _4711_/X vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__a21o_1
X_7500_ _7500_/A _7500_/B _7500_/C _7500_/D vssd1 vssd1 vccd1 vccd1 _7577_/B sky130_fd_sc_hd__nand4_4
X_8480_ _8483_/CLK _8480_/D vssd1 vssd1 vccd1 vccd1 _8480_/Q sky130_fd_sc_hd__dfxtp_1
X_5692_ _5707_/S vssd1 vssd1 vccd1 vccd1 _5701_/S sky130_fd_sc_hd__clkbuf_2
X_4643_ _4653_/A _4653_/B vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__xnor2_4
X_7362_ _7386_/A vssd1 vssd1 vccd1 vccd1 _7362_/X sky130_fd_sc_hd__buf_1
X_4574_ _4410_/X _8157_/Q _4580_/S vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__mux2_1
X_7293_ _8306_/Q _7280_/X _7286_/X _7292_/Y vssd1 vssd1 vccd1 vccd1 _7294_/B sky130_fd_sc_hd__o2bb2a_1
X_6313_ _6352_/A vssd1 vssd1 vccd1 vccd1 _6393_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6244_ _7247_/A _6240_/X _7270_/A _7321_/A vssd1 vssd1 vccd1 vccd1 _7775_/D sky130_fd_sc_hd__a211o_4
XFILLER_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6175_ _6167_/X _7956_/Q _6170_/X _6172_/X _7745_/Q vssd1 vssd1 vccd1 vccd1 _7745_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5126_ _5062_/X _5125_/X _5056_/X vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__a21o_1
X_5057_ _5048_/X _5053_/X _5056_/X vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4008_ _4008_/A vssd1 vssd1 vccd1 vccd1 _8393_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3241_ clkbuf_0__3241_/X vssd1 vssd1 vccd1 vccd1 _6663__315/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__clkbuf_1
X_6690__336 _6694__340/A vssd1 vssd1 vccd1 vccd1 _8000_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3757_ _7633_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3757_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3439_ clkbuf_0__3439_/X vssd1 vssd1 vccd1 vccd1 _7110__77/A sky130_fd_sc_hd__clkbuf_4
X_6996__486 _6999__489/A vssd1 vssd1 vccd1 vccd1 _8167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7109__76 _7110__77/A vssd1 vssd1 vccd1 vccd1 _8257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4290_ _3916_/X _8270_/Q _4298_/S vssd1 vssd1 vccd1 vccd1 _4291_/A sky130_fd_sc_hd__mux2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7980_ _7980_/CLK _7980_/D vssd1 vssd1 vccd1 vccd1 _7980_/Q sky130_fd_sc_hd__dfxtp_1
X_6901__414 _6902__415/A vssd1 vssd1 vccd1 vccd1 _8092_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6862_ _6862_/A vssd1 vssd1 vccd1 vccd1 _8064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5813_ _3892_/X _7784_/Q _5813_/S vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3611_ _7355_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3611_/X sky130_fd_sc_hd__clkbuf_16
X_6793_ _6359_/X _6763_/Y _6791_/Y _6792_/X vssd1 vssd1 vccd1 vccd1 _6794_/D sky130_fd_sc_hd__o22a_1
X_5744_ _5744_/A vssd1 vssd1 vccd1 vccd1 _7864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5675_ _7895_/Q _4973_/X _5683_/S vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__mux2_1
X_8463_ _8463_/CLK _8463_/D vssd1 vssd1 vccd1 vccd1 _8463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7426__2 _7426__2/A vssd1 vssd1 vccd1 vccd1 _8388_/CLK sky130_fd_sc_hd__inv_2
X_8394_ _8394_/CLK _8394_/D vssd1 vssd1 vccd1 vccd1 _8394_/Q sky130_fd_sc_hd__dfxtp_1
X_4626_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7345_ _8324_/Q _7326_/A _7345_/S vssd1 vssd1 vccd1 vccd1 _7346_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4557_ _4413_/X _8164_/Q _4561_/S vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4488_ _8193_/Q _4241_/X _4492_/S vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__mux2_1
X_7276_ _8300_/Q _7264_/X _7272_/X _7200_/B vssd1 vssd1 vccd1 vccd1 _7277_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6227_ _7774_/Q _7773_/Q vssd1 vssd1 vccd1 vccd1 _6229_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6482_/A vssd1 vssd1 vccd1 vccd1 _7678_/A sky130_fd_sc_hd__clkbuf_2
X_5109_ _8472_/Q _8213_/Q _8205_/Q _8237_/Q _5060_/A _5044_/A vssd1 vssd1 vccd1 vccd1
+ _5110_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _7752_/Q _6111_/A vssd1 vssd1 vccd1 vccd1 _6089_/X sky130_fd_sc_hd__or2_1
X_6841__383 _6841__383/A vssd1 vssd1 vccd1 vccd1 _8051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3224_ clkbuf_0__3224_/X vssd1 vssd1 vccd1 vccd1 _6527__250/A sky130_fd_sc_hd__clkbuf_4
X_6505__231 _6509__235/A vssd1 vssd1 vccd1 vccd1 _7871_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460_ _8010_/Q _4448_/X _5464_/S vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4411_ _4410_/X _8221_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _5391_/A vssd1 vssd1 vccd1 vccd1 _8045_/D sky130_fd_sc_hd__clkbuf_1
X_4342_ _4342_/A vssd1 vssd1 vccd1 vccd1 _4342_/X sky130_fd_sc_hd__buf_2
X_4273_ _8277_/Q _4182_/X _4279_/S vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6012_ _6012_/A vssd1 vssd1 vccd1 vccd1 _6085_/A sky130_fd_sc_hd__buf_2
.ends

