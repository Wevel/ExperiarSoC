magic
tech sky130A
magscale 1 2
timestamp 1653090679
<< obsli1 >>
rect 1104 2159 58880 37553
<< obsm1 >>
rect 198 1504 59694 37584
<< metal2 >>
rect 3698 39200 3754 40000
rect 11150 39200 11206 40000
rect 18694 39200 18750 40000
rect 26146 39200 26202 40000
rect 33690 39200 33746 40000
rect 41142 39200 41198 40000
rect 48686 39200 48742 40000
rect 56138 39200 56194 40000
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
<< obsm2 >>
rect 204 39144 3642 39817
rect 3810 39144 11094 39817
rect 11262 39144 18638 39817
rect 18806 39144 26090 39817
rect 26258 39144 33634 39817
rect 33802 39144 41086 39817
rect 41254 39144 48630 39817
rect 48798 39144 56082 39817
rect 56250 39144 59688 39817
rect 204 856 59688 39144
rect 314 167 606 856
rect 774 167 1066 856
rect 1234 167 1526 856
rect 1694 167 2078 856
rect 2246 167 2538 856
rect 2706 167 2998 856
rect 3166 167 3550 856
rect 3718 167 4010 856
rect 4178 167 4470 856
rect 4638 167 5022 856
rect 5190 167 5482 856
rect 5650 167 5942 856
rect 6110 167 6402 856
rect 6570 167 6954 856
rect 7122 167 7414 856
rect 7582 167 7874 856
rect 8042 167 8426 856
rect 8594 167 8886 856
rect 9054 167 9346 856
rect 9514 167 9898 856
rect 10066 167 10358 856
rect 10526 167 10818 856
rect 10986 167 11278 856
rect 11446 167 11830 856
rect 11998 167 12290 856
rect 12458 167 12750 856
rect 12918 167 13302 856
rect 13470 167 13762 856
rect 13930 167 14222 856
rect 14390 167 14774 856
rect 14942 167 15234 856
rect 15402 167 15694 856
rect 15862 167 16154 856
rect 16322 167 16706 856
rect 16874 167 17166 856
rect 17334 167 17626 856
rect 17794 167 18178 856
rect 18346 167 18638 856
rect 18806 167 19098 856
rect 19266 167 19650 856
rect 19818 167 20110 856
rect 20278 167 20570 856
rect 20738 167 21030 856
rect 21198 167 21582 856
rect 21750 167 22042 856
rect 22210 167 22502 856
rect 22670 167 23054 856
rect 23222 167 23514 856
rect 23682 167 23974 856
rect 24142 167 24526 856
rect 24694 167 24986 856
rect 25154 167 25446 856
rect 25614 167 25906 856
rect 26074 167 26458 856
rect 26626 167 26918 856
rect 27086 167 27378 856
rect 27546 167 27930 856
rect 28098 167 28390 856
rect 28558 167 28850 856
rect 29018 167 29402 856
rect 29570 167 29862 856
rect 30030 167 30322 856
rect 30490 167 30782 856
rect 30950 167 31334 856
rect 31502 167 31794 856
rect 31962 167 32254 856
rect 32422 167 32806 856
rect 32974 167 33266 856
rect 33434 167 33726 856
rect 33894 167 34278 856
rect 34446 167 34738 856
rect 34906 167 35198 856
rect 35366 167 35658 856
rect 35826 167 36210 856
rect 36378 167 36670 856
rect 36838 167 37130 856
rect 37298 167 37682 856
rect 37850 167 38142 856
rect 38310 167 38602 856
rect 38770 167 39154 856
rect 39322 167 39614 856
rect 39782 167 40074 856
rect 40242 167 40534 856
rect 40702 167 41086 856
rect 41254 167 41546 856
rect 41714 167 42006 856
rect 42174 167 42558 856
rect 42726 167 43018 856
rect 43186 167 43478 856
rect 43646 167 44030 856
rect 44198 167 44490 856
rect 44658 167 44950 856
rect 45118 167 45410 856
rect 45578 167 45962 856
rect 46130 167 46422 856
rect 46590 167 46882 856
rect 47050 167 47434 856
rect 47602 167 47894 856
rect 48062 167 48354 856
rect 48522 167 48906 856
rect 49074 167 49366 856
rect 49534 167 49826 856
rect 49994 167 50286 856
rect 50454 167 50838 856
rect 51006 167 51298 856
rect 51466 167 51758 856
rect 51926 167 52310 856
rect 52478 167 52770 856
rect 52938 167 53230 856
rect 53398 167 53782 856
rect 53950 167 54242 856
rect 54410 167 54702 856
rect 54870 167 55162 856
rect 55330 167 55714 856
rect 55882 167 56174 856
rect 56342 167 56634 856
rect 56802 167 57186 856
rect 57354 167 57646 856
rect 57814 167 58106 856
rect 58274 167 58658 856
rect 58826 167 59118 856
rect 59286 167 59578 856
<< metal3 >>
rect 0 39720 800 39840
rect 0 39312 800 39432
rect 0 38904 800 39024
rect 0 38496 800 38616
rect 0 38088 800 38208
rect 0 37680 800 37800
rect 0 37272 800 37392
rect 0 36864 800 36984
rect 0 36456 800 36576
rect 0 36048 800 36168
rect 0 35640 800 35760
rect 0 35232 800 35352
rect 0 34824 800 34944
rect 0 34416 800 34536
rect 0 34008 800 34128
rect 0 33600 800 33720
rect 0 33328 800 33448
rect 0 32920 800 33040
rect 0 32512 800 32632
rect 0 32104 800 32224
rect 0 31696 800 31816
rect 0 31288 800 31408
rect 0 30880 800 31000
rect 0 30472 800 30592
rect 0 30064 800 30184
rect 0 29656 800 29776
rect 0 29248 800 29368
rect 0 28840 800 28960
rect 0 28432 800 28552
rect 0 28024 800 28144
rect 0 27616 800 27736
rect 0 27208 800 27328
rect 0 26800 800 26920
rect 0 26528 800 26648
rect 0 26120 800 26240
rect 0 25712 800 25832
rect 0 25304 800 25424
rect 0 24896 800 25016
rect 0 24488 800 24608
rect 0 24080 800 24200
rect 0 23672 800 23792
rect 0 23264 800 23384
rect 0 22856 800 22976
rect 0 22448 800 22568
rect 0 22040 800 22160
rect 0 21632 800 21752
rect 0 21224 800 21344
rect 0 20816 800 20936
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19320 800 19440
rect 0 18912 800 19032
rect 0 18504 800 18624
rect 0 18096 800 18216
rect 0 17688 800 17808
rect 0 17280 800 17400
rect 0 16872 800 16992
rect 0 16464 800 16584
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 0 15240 800 15360
rect 0 14832 800 14952
rect 0 14424 800 14544
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 12112 800 12232
rect 0 11704 800 11824
rect 0 11296 800 11416
rect 0 10888 800 11008
rect 0 10480 800 10600
rect 0 10072 800 10192
rect 0 9664 800 9784
rect 0 9256 800 9376
rect 0 8848 800 8968
rect 0 8440 800 8560
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6808 800 6928
rect 0 6536 800 6656
rect 0 6128 800 6248
rect 0 5720 800 5840
rect 0 5312 800 5432
rect 0 4904 800 5024
rect 0 4496 800 4616
rect 0 4088 800 4208
rect 0 3680 800 3800
rect 0 3272 800 3392
rect 0 2864 800 2984
rect 0 2456 800 2576
rect 0 2048 800 2168
rect 0 1640 800 1760
rect 0 1232 800 1352
rect 0 824 800 944
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 39640 55923 39813
rect 800 39512 55923 39640
rect 880 39232 55923 39512
rect 800 39104 55923 39232
rect 880 38824 55923 39104
rect 800 38696 55923 38824
rect 880 38416 55923 38696
rect 800 38288 55923 38416
rect 880 38008 55923 38288
rect 800 37880 55923 38008
rect 880 37600 55923 37880
rect 800 37472 55923 37600
rect 880 37192 55923 37472
rect 800 37064 55923 37192
rect 880 36784 55923 37064
rect 800 36656 55923 36784
rect 880 36376 55923 36656
rect 800 36248 55923 36376
rect 880 35968 55923 36248
rect 800 35840 55923 35968
rect 880 35560 55923 35840
rect 800 35432 55923 35560
rect 880 35152 55923 35432
rect 800 35024 55923 35152
rect 880 34744 55923 35024
rect 800 34616 55923 34744
rect 880 34336 55923 34616
rect 800 34208 55923 34336
rect 880 33928 55923 34208
rect 800 33800 55923 33928
rect 880 33248 55923 33800
rect 800 33120 55923 33248
rect 880 32840 55923 33120
rect 800 32712 55923 32840
rect 880 32432 55923 32712
rect 800 32304 55923 32432
rect 880 32024 55923 32304
rect 800 31896 55923 32024
rect 880 31616 55923 31896
rect 800 31488 55923 31616
rect 880 31208 55923 31488
rect 800 31080 55923 31208
rect 880 30800 55923 31080
rect 800 30672 55923 30800
rect 880 30392 55923 30672
rect 800 30264 55923 30392
rect 880 29984 55923 30264
rect 800 29856 55923 29984
rect 880 29576 55923 29856
rect 800 29448 55923 29576
rect 880 29168 55923 29448
rect 800 29040 55923 29168
rect 880 28760 55923 29040
rect 800 28632 55923 28760
rect 880 28352 55923 28632
rect 800 28224 55923 28352
rect 880 27944 55923 28224
rect 800 27816 55923 27944
rect 880 27536 55923 27816
rect 800 27408 55923 27536
rect 880 27128 55923 27408
rect 800 27000 55923 27128
rect 880 26448 55923 27000
rect 800 26320 55923 26448
rect 880 26040 55923 26320
rect 800 25912 55923 26040
rect 880 25632 55923 25912
rect 800 25504 55923 25632
rect 880 25224 55923 25504
rect 800 25096 55923 25224
rect 880 24816 55923 25096
rect 800 24688 55923 24816
rect 880 24408 55923 24688
rect 800 24280 55923 24408
rect 880 24000 55923 24280
rect 800 23872 55923 24000
rect 880 23592 55923 23872
rect 800 23464 55923 23592
rect 880 23184 55923 23464
rect 800 23056 55923 23184
rect 880 22776 55923 23056
rect 800 22648 55923 22776
rect 880 22368 55923 22648
rect 800 22240 55923 22368
rect 880 21960 55923 22240
rect 800 21832 55923 21960
rect 880 21552 55923 21832
rect 800 21424 55923 21552
rect 880 21144 55923 21424
rect 800 21016 55923 21144
rect 880 20736 55923 21016
rect 800 20608 55923 20736
rect 880 20056 55923 20608
rect 800 19928 55923 20056
rect 880 19648 55923 19928
rect 800 19520 55923 19648
rect 880 19240 55923 19520
rect 800 19112 55923 19240
rect 880 18832 55923 19112
rect 800 18704 55923 18832
rect 880 18424 55923 18704
rect 800 18296 55923 18424
rect 880 18016 55923 18296
rect 800 17888 55923 18016
rect 880 17608 55923 17888
rect 800 17480 55923 17608
rect 880 17200 55923 17480
rect 800 17072 55923 17200
rect 880 16792 55923 17072
rect 800 16664 55923 16792
rect 880 16384 55923 16664
rect 800 16256 55923 16384
rect 880 15976 55923 16256
rect 800 15848 55923 15976
rect 880 15568 55923 15848
rect 800 15440 55923 15568
rect 880 15160 55923 15440
rect 800 15032 55923 15160
rect 880 14752 55923 15032
rect 800 14624 55923 14752
rect 880 14344 55923 14624
rect 800 14216 55923 14344
rect 880 13936 55923 14216
rect 800 13808 55923 13936
rect 880 13256 55923 13808
rect 800 13128 55923 13256
rect 880 12848 55923 13128
rect 800 12720 55923 12848
rect 880 12440 55923 12720
rect 800 12312 55923 12440
rect 880 12032 55923 12312
rect 800 11904 55923 12032
rect 880 11624 55923 11904
rect 800 11496 55923 11624
rect 880 11216 55923 11496
rect 800 11088 55923 11216
rect 880 10808 55923 11088
rect 800 10680 55923 10808
rect 880 10400 55923 10680
rect 800 10272 55923 10400
rect 880 9992 55923 10272
rect 800 9864 55923 9992
rect 880 9584 55923 9864
rect 800 9456 55923 9584
rect 880 9176 55923 9456
rect 800 9048 55923 9176
rect 880 8768 55923 9048
rect 800 8640 55923 8768
rect 880 8360 55923 8640
rect 800 8232 55923 8360
rect 880 7952 55923 8232
rect 800 7824 55923 7952
rect 880 7544 55923 7824
rect 800 7416 55923 7544
rect 880 7136 55923 7416
rect 800 7008 55923 7136
rect 880 6456 55923 7008
rect 800 6328 55923 6456
rect 880 6048 55923 6328
rect 800 5920 55923 6048
rect 880 5640 55923 5920
rect 800 5512 55923 5640
rect 880 5232 55923 5512
rect 800 5104 55923 5232
rect 880 4824 55923 5104
rect 800 4696 55923 4824
rect 880 4416 55923 4696
rect 800 4288 55923 4416
rect 880 4008 55923 4288
rect 800 3880 55923 4008
rect 880 3600 55923 3880
rect 800 3472 55923 3600
rect 880 3192 55923 3472
rect 800 3064 55923 3192
rect 880 2784 55923 3064
rect 800 2656 55923 2784
rect 880 2376 55923 2656
rect 800 2248 55923 2376
rect 880 1968 55923 2248
rect 800 1840 55923 1968
rect 880 1560 55923 1840
rect 800 1432 55923 1560
rect 880 1152 55923 1432
rect 800 1024 55923 1152
rect 880 744 55923 1024
rect 800 616 55923 744
rect 880 171 55923 616
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
<< labels >>
rlabel metal2 s 3698 39200 3754 40000 6 flash_csb
port 1 nsew signal output
rlabel metal2 s 11150 39200 11206 40000 6 flash_io0_read
port 2 nsew signal input
rlabel metal2 s 18694 39200 18750 40000 6 flash_io0_we
port 3 nsew signal output
rlabel metal2 s 26146 39200 26202 40000 6 flash_io0_write
port 4 nsew signal output
rlabel metal2 s 33690 39200 33746 40000 6 flash_io1_read
port 5 nsew signal input
rlabel metal2 s 41142 39200 41198 40000 6 flash_io1_we
port 6 nsew signal output
rlabel metal2 s 48686 39200 48742 40000 6 flash_io1_write
port 7 nsew signal output
rlabel metal2 s 56138 39200 56194 40000 6 flash_sck
port 8 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 sram_addr0[0]
port 9 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 sram_addr0[1]
port 10 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 sram_addr0[2]
port 11 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 sram_addr0[3]
port 12 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[4]
port 13 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 sram_addr0[5]
port 14 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 sram_addr0[6]
port 15 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 sram_addr0[7]
port 16 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 sram_addr0[8]
port 17 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 sram_addr1[0]
port 18 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 sram_addr1[1]
port 19 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 sram_addr1[2]
port 20 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 sram_addr1[3]
port 21 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 sram_addr1[4]
port 22 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 sram_addr1[5]
port 23 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 sram_addr1[6]
port 24 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 sram_addr1[7]
port 25 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 sram_addr1[8]
port 26 nsew signal output
rlabel metal2 s 202 0 258 800 6 sram_clk0
port 27 nsew signal output
rlabel metal2 s 662 0 718 800 6 sram_clk1
port 28 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 sram_csb0
port 29 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 sram_csb1
port 30 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 sram_din0[0]
port 31 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 sram_din0[10]
port 32 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 33 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 34 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 sram_din0[13]
port 35 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 sram_din0[14]
port 36 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 sram_din0[15]
port 37 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 sram_din0[16]
port 38 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 sram_din0[17]
port 39 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 sram_din0[18]
port 40 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 sram_din0[19]
port 41 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 sram_din0[1]
port 42 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 sram_din0[20]
port 43 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 sram_din0[21]
port 44 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 sram_din0[22]
port 45 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 sram_din0[23]
port 46 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 sram_din0[24]
port 47 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 sram_din0[25]
port 48 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 sram_din0[26]
port 49 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 sram_din0[27]
port 50 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 sram_din0[28]
port 51 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 sram_din0[29]
port 52 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 sram_din0[2]
port 53 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 sram_din0[30]
port 54 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 sram_din0[31]
port 55 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 sram_din0[3]
port 56 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 sram_din0[4]
port 57 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 sram_din0[5]
port 58 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 sram_din0[6]
port 59 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 sram_din0[7]
port 60 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 sram_din0[8]
port 61 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 sram_din0[9]
port 62 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 sram_dout0[0]
port 63 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 sram_dout0[10]
port 64 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 65 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 sram_dout0[12]
port 66 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sram_dout0[13]
port 67 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 sram_dout0[14]
port 68 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout0[15]
port 69 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 sram_dout0[16]
port 70 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout0[17]
port 71 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 sram_dout0[18]
port 72 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 sram_dout0[19]
port 73 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 sram_dout0[1]
port 74 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[20]
port 75 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 sram_dout0[21]
port 76 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 sram_dout0[22]
port 77 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout0[23]
port 78 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 sram_dout0[24]
port 79 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 sram_dout0[25]
port 80 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 sram_dout0[26]
port 81 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 sram_dout0[27]
port 82 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[28]
port 83 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout0[29]
port 84 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 sram_dout0[2]
port 85 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 sram_dout0[30]
port 86 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 sram_dout0[31]
port 87 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 sram_dout0[3]
port 88 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 sram_dout0[4]
port 89 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 sram_dout0[5]
port 90 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 sram_dout0[6]
port 91 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 sram_dout0[7]
port 92 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 sram_dout0[8]
port 93 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 sram_dout0[9]
port 94 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 sram_dout1[0]
port 95 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 sram_dout1[10]
port 96 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 97 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 sram_dout1[12]
port 98 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 sram_dout1[13]
port 99 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 sram_dout1[14]
port 100 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 sram_dout1[15]
port 101 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 sram_dout1[16]
port 102 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 sram_dout1[17]
port 103 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 sram_dout1[18]
port 104 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 sram_dout1[19]
port 105 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 sram_dout1[1]
port 106 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 sram_dout1[20]
port 107 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 sram_dout1[21]
port 108 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout1[22]
port 109 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 sram_dout1[23]
port 110 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 sram_dout1[24]
port 111 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 sram_dout1[25]
port 112 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[26]
port 113 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[27]
port 114 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[28]
port 115 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 sram_dout1[29]
port 116 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 sram_dout1[2]
port 117 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 sram_dout1[30]
port 118 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 sram_dout1[31]
port 119 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 sram_dout1[3]
port 120 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 sram_dout1[4]
port 121 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 sram_dout1[5]
port 122 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 sram_dout1[6]
port 123 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 sram_dout1[7]
port 124 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout1[8]
port 125 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[9]
port 126 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 sram_web0
port 127 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 sram_wmask0[0]
port 128 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 sram_wmask0[1]
port 129 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 sram_wmask0[2]
port 130 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 sram_wmask0[3]
port 131 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 134 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 wb_adr_i[0]
port 135 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wb_adr_i[10]
port 136 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_adr_i[11]
port 137 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 wb_adr_i[12]
port 138 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 wb_adr_i[13]
port 139 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wb_adr_i[14]
port 140 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 wb_adr_i[15]
port 141 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wb_adr_i[16]
port 142 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wb_adr_i[17]
port 143 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wb_adr_i[18]
port 144 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 wb_adr_i[19]
port 145 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 wb_adr_i[1]
port 146 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 wb_adr_i[20]
port 147 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 wb_adr_i[21]
port 148 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wb_adr_i[22]
port 149 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 wb_adr_i[23]
port 150 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 wb_adr_i[2]
port 151 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 wb_adr_i[3]
port 152 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 wb_adr_i[4]
port 153 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wb_adr_i[5]
port 154 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 wb_adr_i[6]
port 155 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 wb_adr_i[7]
port 156 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wb_adr_i[8]
port 157 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wb_adr_i[9]
port 158 nsew signal input
rlabel metal3 s 0 416 800 536 6 wb_clk_i
port 159 nsew signal input
rlabel metal3 s 0 824 800 944 6 wb_cyc_i
port 160 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 wb_data_i[0]
port 161 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 wb_data_i[10]
port 162 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wb_data_i[11]
port 163 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 wb_data_i[12]
port 164 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 wb_data_i[13]
port 165 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 wb_data_i[14]
port 166 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 wb_data_i[15]
port 167 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[16]
port 168 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[17]
port 169 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wb_data_i[18]
port 170 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 wb_data_i[19]
port 171 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 wb_data_i[1]
port 172 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wb_data_i[20]
port 173 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 wb_data_i[21]
port 174 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 wb_data_i[22]
port 175 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_data_i[23]
port 176 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 wb_data_i[24]
port 177 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 wb_data_i[25]
port 178 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 wb_data_i[26]
port 179 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 wb_data_i[27]
port 180 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 wb_data_i[28]
port 181 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 wb_data_i[29]
port 182 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_data_i[2]
port 183 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 wb_data_i[30]
port 184 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 wb_data_i[31]
port 185 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_data_i[3]
port 186 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 wb_data_i[4]
port 187 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 wb_data_i[5]
port 188 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 wb_data_i[6]
port 189 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wb_data_i[7]
port 190 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 wb_data_i[8]
port 191 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wb_data_i[9]
port 192 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wb_data_o[0]
port 193 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 wb_data_o[10]
port 194 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 wb_data_o[11]
port 195 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 wb_data_o[12]
port 196 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 wb_data_o[13]
port 197 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 wb_data_o[14]
port 198 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 wb_data_o[15]
port 199 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 wb_data_o[16]
port 200 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 wb_data_o[17]
port 201 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 wb_data_o[18]
port 202 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 wb_data_o[19]
port 203 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 wb_data_o[1]
port 204 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 wb_data_o[20]
port 205 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 wb_data_o[21]
port 206 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 wb_data_o[22]
port 207 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 wb_data_o[23]
port 208 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 wb_data_o[24]
port 209 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 wb_data_o[25]
port 210 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 wb_data_o[26]
port 211 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 wb_data_o[27]
port 212 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 wb_data_o[28]
port 213 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 wb_data_o[29]
port 214 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 wb_data_o[2]
port 215 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 wb_data_o[30]
port 216 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 wb_data_o[31]
port 217 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 wb_data_o[3]
port 218 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 wb_data_o[4]
port 219 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 wb_data_o[5]
port 220 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 wb_data_o[6]
port 221 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 wb_data_o[7]
port 222 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 wb_data_o[8]
port 223 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 wb_data_o[9]
port 224 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 wb_error_o
port 225 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 wb_rst_i
port 226 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 wb_sel_i[0]
port 227 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wb_sel_i[1]
port 228 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wb_sel_i[2]
port 229 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 wb_sel_i[3]
port 230 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 wb_stall_o
port 231 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 wb_stb_i
port 232 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 wb_we_i
port 233 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1272638
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Flash/runs/Flash/results/signoff/Flash.magic.gds
string GDS_START 156742
<< end >>

