magic
tech sky130A
magscale 1 2
timestamp 1651273041
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 1104 2128 68816 67504
<< metal2 >>
rect 17498 0 17554 800
rect 52458 0 52514 800
<< obsm2 >>
rect 1398 856 68154 67504
rect 1398 575 17442 856
rect 17610 575 52402 856
rect 52570 575 68154 856
<< metal3 >>
rect 0 69368 800 69488
rect 0 68144 800 68264
rect 0 66920 800 67040
rect 69200 67056 70000 67176
rect 0 65832 800 65952
rect 0 64608 800 64728
rect 0 63384 800 63504
rect 0 62160 800 62280
rect 0 61072 800 61192
rect 69200 61208 70000 61328
rect 0 59848 800 59968
rect 0 58624 800 58744
rect 0 57400 800 57520
rect 0 56312 800 56432
rect 69200 55360 70000 55480
rect 0 55088 800 55208
rect 0 53864 800 53984
rect 0 52776 800 52896
rect 0 51552 800 51672
rect 0 50328 800 50448
rect 69200 49512 70000 49632
rect 0 49104 800 49224
rect 0 48016 800 48136
rect 0 46792 800 46912
rect 0 45568 800 45688
rect 0 44344 800 44464
rect 69200 43664 70000 43784
rect 0 43256 800 43376
rect 0 42032 800 42152
rect 0 40808 800 40928
rect 0 39720 800 39840
rect 0 38496 800 38616
rect 69200 37816 70000 37936
rect 0 37272 800 37392
rect 0 36048 800 36168
rect 0 34960 800 35080
rect 0 33736 800 33856
rect 0 32512 800 32632
rect 69200 31968 70000 32088
rect 0 31288 800 31408
rect 0 30200 800 30320
rect 0 28976 800 29096
rect 0 27752 800 27872
rect 0 26664 800 26784
rect 69200 26120 70000 26240
rect 0 25440 800 25560
rect 0 24216 800 24336
rect 0 22992 800 23112
rect 0 21904 800 22024
rect 0 20680 800 20800
rect 69200 20272 70000 20392
rect 0 19456 800 19576
rect 0 18232 800 18352
rect 0 17144 800 17264
rect 0 15920 800 16040
rect 0 14696 800 14816
rect 69200 14424 70000 14544
rect 0 13608 800 13728
rect 0 12384 800 12504
rect 0 11160 800 11280
rect 0 9936 800 10056
rect 0 8848 800 8968
rect 69200 8576 70000 8696
rect 0 7624 800 7744
rect 0 6400 800 6520
rect 0 5176 800 5296
rect 0 4088 800 4208
rect 0 2864 800 2984
rect 69200 2864 70000 2984
rect 0 1640 800 1760
rect 0 552 800 672
<< obsm3 >>
rect 800 67256 69200 67489
rect 800 67120 69120 67256
rect 880 66976 69120 67120
rect 880 66840 69200 66976
rect 800 66032 69200 66840
rect 880 65752 69200 66032
rect 800 64808 69200 65752
rect 880 64528 69200 64808
rect 800 63584 69200 64528
rect 880 63304 69200 63584
rect 800 62360 69200 63304
rect 880 62080 69200 62360
rect 800 61408 69200 62080
rect 800 61272 69120 61408
rect 880 61128 69120 61272
rect 880 60992 69200 61128
rect 800 60048 69200 60992
rect 880 59768 69200 60048
rect 800 58824 69200 59768
rect 880 58544 69200 58824
rect 800 57600 69200 58544
rect 880 57320 69200 57600
rect 800 56512 69200 57320
rect 880 56232 69200 56512
rect 800 55560 69200 56232
rect 800 55288 69120 55560
rect 880 55280 69120 55288
rect 880 55008 69200 55280
rect 800 54064 69200 55008
rect 880 53784 69200 54064
rect 800 52976 69200 53784
rect 880 52696 69200 52976
rect 800 51752 69200 52696
rect 880 51472 69200 51752
rect 800 50528 69200 51472
rect 880 50248 69200 50528
rect 800 49712 69200 50248
rect 800 49432 69120 49712
rect 800 49304 69200 49432
rect 880 49024 69200 49304
rect 800 48216 69200 49024
rect 880 47936 69200 48216
rect 800 46992 69200 47936
rect 880 46712 69200 46992
rect 800 45768 69200 46712
rect 880 45488 69200 45768
rect 800 44544 69200 45488
rect 880 44264 69200 44544
rect 800 43864 69200 44264
rect 800 43584 69120 43864
rect 800 43456 69200 43584
rect 880 43176 69200 43456
rect 800 42232 69200 43176
rect 880 41952 69200 42232
rect 800 41008 69200 41952
rect 880 40728 69200 41008
rect 800 39920 69200 40728
rect 880 39640 69200 39920
rect 800 38696 69200 39640
rect 880 38416 69200 38696
rect 800 38016 69200 38416
rect 800 37736 69120 38016
rect 800 37472 69200 37736
rect 880 37192 69200 37472
rect 800 36248 69200 37192
rect 880 35968 69200 36248
rect 800 35160 69200 35968
rect 880 34880 69200 35160
rect 800 33936 69200 34880
rect 880 33656 69200 33936
rect 800 32712 69200 33656
rect 880 32432 69200 32712
rect 800 32168 69200 32432
rect 800 31888 69120 32168
rect 800 31488 69200 31888
rect 880 31208 69200 31488
rect 800 30400 69200 31208
rect 880 30120 69200 30400
rect 800 29176 69200 30120
rect 880 28896 69200 29176
rect 800 27952 69200 28896
rect 880 27672 69200 27952
rect 800 26864 69200 27672
rect 880 26584 69200 26864
rect 800 26320 69200 26584
rect 800 26040 69120 26320
rect 800 25640 69200 26040
rect 880 25360 69200 25640
rect 800 24416 69200 25360
rect 880 24136 69200 24416
rect 800 23192 69200 24136
rect 880 22912 69200 23192
rect 800 22104 69200 22912
rect 880 21824 69200 22104
rect 800 20880 69200 21824
rect 880 20600 69200 20880
rect 800 20472 69200 20600
rect 800 20192 69120 20472
rect 800 19656 69200 20192
rect 880 19376 69200 19656
rect 800 18432 69200 19376
rect 880 18152 69200 18432
rect 800 17344 69200 18152
rect 880 17064 69200 17344
rect 800 16120 69200 17064
rect 880 15840 69200 16120
rect 800 14896 69200 15840
rect 880 14624 69200 14896
rect 880 14616 69120 14624
rect 800 14344 69120 14616
rect 800 13808 69200 14344
rect 880 13528 69200 13808
rect 800 12584 69200 13528
rect 880 12304 69200 12584
rect 800 11360 69200 12304
rect 880 11080 69200 11360
rect 800 10136 69200 11080
rect 880 9856 69200 10136
rect 800 9048 69200 9856
rect 880 8776 69200 9048
rect 880 8768 69120 8776
rect 800 8496 69120 8768
rect 800 7824 69200 8496
rect 880 7544 69200 7824
rect 800 6600 69200 7544
rect 880 6320 69200 6600
rect 800 5376 69200 6320
rect 880 5096 69200 5376
rect 800 4288 69200 5096
rect 880 4008 69200 4288
rect 800 3064 69200 4008
rect 880 2784 69120 3064
rect 800 1840 69200 2784
rect 880 1560 69200 1840
rect 800 752 69200 1560
rect 880 579 69200 752
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< labels >>
rlabel metal2 s 17498 0 17554 800 6 clk
port 1 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 peripheralBus_address[0]
port 2 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 peripheralBus_address[10]
port 3 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 peripheralBus_address[11]
port 4 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 peripheralBus_address[12]
port 5 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 peripheralBus_address[13]
port 6 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 peripheralBus_address[14]
port 7 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 peripheralBus_address[15]
port 8 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 peripheralBus_address[16]
port 9 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 peripheralBus_address[17]
port 10 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 peripheralBus_address[18]
port 11 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 peripheralBus_address[19]
port 12 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 peripheralBus_address[1]
port 13 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 peripheralBus_address[20]
port 14 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 peripheralBus_address[21]
port 15 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 peripheralBus_address[22]
port 16 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 peripheralBus_address[23]
port 17 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 peripheralBus_address[2]
port 18 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 peripheralBus_address[3]
port 19 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 peripheralBus_address[4]
port 20 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 peripheralBus_address[5]
port 21 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 peripheralBus_address[6]
port 22 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 peripheralBus_address[7]
port 23 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 peripheralBus_address[8]
port 24 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 peripheralBus_address[9]
port 25 nsew signal input
rlabel metal3 s 0 552 800 672 6 peripheralBus_busy
port 26 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 peripheralBus_data[0]
port 27 nsew signal bidirectional
rlabel metal3 s 0 28976 800 29096 6 peripheralBus_data[10]
port 28 nsew signal bidirectional
rlabel metal3 s 0 31288 800 31408 6 peripheralBus_data[11]
port 29 nsew signal bidirectional
rlabel metal3 s 0 33736 800 33856 6 peripheralBus_data[12]
port 30 nsew signal bidirectional
rlabel metal3 s 0 36048 800 36168 6 peripheralBus_data[13]
port 31 nsew signal bidirectional
rlabel metal3 s 0 38496 800 38616 6 peripheralBus_data[14]
port 32 nsew signal bidirectional
rlabel metal3 s 0 40808 800 40928 6 peripheralBus_data[15]
port 33 nsew signal bidirectional
rlabel metal3 s 0 43256 800 43376 6 peripheralBus_data[16]
port 34 nsew signal bidirectional
rlabel metal3 s 0 45568 800 45688 6 peripheralBus_data[17]
port 35 nsew signal bidirectional
rlabel metal3 s 0 48016 800 48136 6 peripheralBus_data[18]
port 36 nsew signal bidirectional
rlabel metal3 s 0 50328 800 50448 6 peripheralBus_data[19]
port 37 nsew signal bidirectional
rlabel metal3 s 0 7624 800 7744 6 peripheralBus_data[1]
port 38 nsew signal bidirectional
rlabel metal3 s 0 52776 800 52896 6 peripheralBus_data[20]
port 39 nsew signal bidirectional
rlabel metal3 s 0 55088 800 55208 6 peripheralBus_data[21]
port 40 nsew signal bidirectional
rlabel metal3 s 0 57400 800 57520 6 peripheralBus_data[22]
port 41 nsew signal bidirectional
rlabel metal3 s 0 59848 800 59968 6 peripheralBus_data[23]
port 42 nsew signal bidirectional
rlabel metal3 s 0 61072 800 61192 6 peripheralBus_data[24]
port 43 nsew signal bidirectional
rlabel metal3 s 0 62160 800 62280 6 peripheralBus_data[25]
port 44 nsew signal bidirectional
rlabel metal3 s 0 63384 800 63504 6 peripheralBus_data[26]
port 45 nsew signal bidirectional
rlabel metal3 s 0 64608 800 64728 6 peripheralBus_data[27]
port 46 nsew signal bidirectional
rlabel metal3 s 0 65832 800 65952 6 peripheralBus_data[28]
port 47 nsew signal bidirectional
rlabel metal3 s 0 66920 800 67040 6 peripheralBus_data[29]
port 48 nsew signal bidirectional
rlabel metal3 s 0 9936 800 10056 6 peripheralBus_data[2]
port 49 nsew signal bidirectional
rlabel metal3 s 0 68144 800 68264 6 peripheralBus_data[30]
port 50 nsew signal bidirectional
rlabel metal3 s 0 69368 800 69488 6 peripheralBus_data[31]
port 51 nsew signal bidirectional
rlabel metal3 s 0 12384 800 12504 6 peripheralBus_data[3]
port 52 nsew signal bidirectional
rlabel metal3 s 0 14696 800 14816 6 peripheralBus_data[4]
port 53 nsew signal bidirectional
rlabel metal3 s 0 17144 800 17264 6 peripheralBus_data[5]
port 54 nsew signal bidirectional
rlabel metal3 s 0 19456 800 19576 6 peripheralBus_data[6]
port 55 nsew signal bidirectional
rlabel metal3 s 0 21904 800 22024 6 peripheralBus_data[7]
port 56 nsew signal bidirectional
rlabel metal3 s 0 24216 800 24336 6 peripheralBus_data[8]
port 57 nsew signal bidirectional
rlabel metal3 s 0 26664 800 26784 6 peripheralBus_data[9]
port 58 nsew signal bidirectional
rlabel metal3 s 0 1640 800 1760 6 peripheralBus_oe
port 59 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 peripheralBus_we
port 60 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 rst
port 61 nsew signal input
rlabel metal3 s 69200 2864 70000 2984 6 uart_en[0]
port 62 nsew signal output
rlabel metal3 s 69200 20272 70000 20392 6 uart_en[1]
port 63 nsew signal output
rlabel metal3 s 69200 37816 70000 37936 6 uart_en[2]
port 64 nsew signal output
rlabel metal3 s 69200 55360 70000 55480 6 uart_en[3]
port 65 nsew signal output
rlabel metal3 s 69200 8576 70000 8696 6 uart_rx[0]
port 66 nsew signal output
rlabel metal3 s 69200 26120 70000 26240 6 uart_rx[1]
port 67 nsew signal output
rlabel metal3 s 69200 43664 70000 43784 6 uart_rx[2]
port 68 nsew signal output
rlabel metal3 s 69200 61208 70000 61328 6 uart_rx[3]
port 69 nsew signal output
rlabel metal3 s 69200 14424 70000 14544 6 uart_tx[0]
port 70 nsew signal output
rlabel metal3 s 69200 31968 70000 32088 6 uart_tx[1]
port 71 nsew signal output
rlabel metal3 s 69200 49512 70000 49632 6 uart_tx[2]
port 72 nsew signal output
rlabel metal3 s 69200 67056 70000 67176 6 uart_tx[3]
port 73 nsew signal output
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 74 nsew power input
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 74 nsew power input
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 74 nsew power input
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 75 nsew ground input
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 75 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1234398
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_UART/runs/Peripheral_UART/results/finishing/UART.magic.gds
string GDS_START 24092
<< end >>

