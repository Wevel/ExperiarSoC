magic
tech sky130A
magscale 1 2
timestamp 1650758507
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 38824 37584
<< obsm2 >>
rect 1398 2128 38070 37584
<< metal3 >>
rect 0 29928 800 30048
rect 39200 29928 40000 30048
rect 0 9936 800 10056
rect 39200 9936 40000 10056
<< obsm3 >>
rect 800 30128 39200 37569
rect 880 29848 39120 30128
rect 800 10136 39200 29848
rect 880 9856 39120 10136
rect 800 2143 39200 9856
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 19195 9963 19488 23085
rect 19968 9963 23125 23085
<< labels >>
rlabel metal3 s 39200 29928 40000 30048 6 blink[0]
port 1 nsew signal output
rlabel metal3 s 39200 9936 40000 10056 6 blink[1]
port 2 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 clk
port 3 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 rst
port 4 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 5 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 5 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 6 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 807820
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Blink/runs/Blink/results/finishing/Blink.magic.gds
string GDS_START 123934
<< end >>

