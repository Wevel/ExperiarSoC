VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Video
  CLASS BLOCK ;
  FOREIGN Video ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 500.000 ;
  PIN sram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 17.040 350.000 17.640 ;
    END
  END sram_addr0[0]
  PIN sram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 29.280 350.000 29.880 ;
    END
  END sram_addr0[1]
  PIN sram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 41.520 350.000 42.120 ;
    END
  END sram_addr0[2]
  PIN sram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 53.760 350.000 54.360 ;
    END
  END sram_addr0[3]
  PIN sram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 66.000 350.000 66.600 ;
    END
  END sram_addr0[4]
  PIN sram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 73.480 350.000 74.080 ;
    END
  END sram_addr0[5]
  PIN sram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 80.960 350.000 81.560 ;
    END
  END sram_addr0[6]
  PIN sram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 88.440 350.000 89.040 ;
    END
  END sram_addr0[7]
  PIN sram_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 95.920 350.000 96.520 ;
    END
  END sram_addr0[8]
  PIN sram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 18.400 350.000 19.000 ;
    END
  END sram_addr1[0]
  PIN sram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 30.640 350.000 31.240 ;
    END
  END sram_addr1[1]
  PIN sram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 42.880 350.000 43.480 ;
    END
  END sram_addr1[2]
  PIN sram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 55.120 350.000 55.720 ;
    END
  END sram_addr1[3]
  PIN sram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 67.360 350.000 67.960 ;
    END
  END sram_addr1[4]
  PIN sram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 74.840 350.000 75.440 ;
    END
  END sram_addr1[5]
  PIN sram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 82.320 350.000 82.920 ;
    END
  END sram_addr1[6]
  PIN sram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 89.800 350.000 90.400 ;
    END
  END sram_addr1[7]
  PIN sram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 97.280 350.000 97.880 ;
    END
  END sram_addr1[8]
  PIN sram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 12.280 350.000 12.880 ;
    END
  END sram_clk0
  PIN sram_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 14.320 350.000 14.920 ;
    END
  END sram_clk1
  PIN sram_csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 20.440 350.000 21.040 ;
    END
  END sram_csb0[0]
  PIN sram_csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 32.000 350.000 32.600 ;
    END
  END sram_csb0[1]
  PIN sram_csb0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 44.240 350.000 44.840 ;
    END
  END sram_csb0[2]
  PIN sram_csb0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 56.480 350.000 57.080 ;
    END
  END sram_csb0[3]
  PIN sram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 21.800 350.000 22.400 ;
    END
  END sram_csb1[0]
  PIN sram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.040 350.000 34.640 ;
    END
  END sram_csb1[1]
  PIN sram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 46.280 350.000 46.880 ;
    END
  END sram_csb1[2]
  PIN sram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 57.840 350.000 58.440 ;
    END
  END sram_csb1[3]
  PIN sram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 23.160 350.000 23.760 ;
    END
  END sram_din0[0]
  PIN sram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 108.160 350.000 108.760 ;
    END
  END sram_din0[10]
  PIN sram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 112.920 350.000 113.520 ;
    END
  END sram_din0[11]
  PIN sram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 117.680 350.000 118.280 ;
    END
  END sram_din0[12]
  PIN sram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 121.760 350.000 122.360 ;
    END
  END sram_din0[13]
  PIN sram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 126.520 350.000 127.120 ;
    END
  END sram_din0[14]
  PIN sram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 131.280 350.000 131.880 ;
    END
  END sram_din0[15]
  PIN sram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 135.360 350.000 135.960 ;
    END
  END sram_din0[16]
  PIN sram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 140.120 350.000 140.720 ;
    END
  END sram_din0[17]
  PIN sram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 144.880 350.000 145.480 ;
    END
  END sram_din0[18]
  PIN sram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 148.960 350.000 149.560 ;
    END
  END sram_din0[19]
  PIN sram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 35.400 350.000 36.000 ;
    END
  END sram_din0[1]
  PIN sram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 153.720 350.000 154.320 ;
    END
  END sram_din0[20]
  PIN sram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 158.480 350.000 159.080 ;
    END
  END sram_din0[21]
  PIN sram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 163.240 350.000 163.840 ;
    END
  END sram_din0[22]
  PIN sram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 167.320 350.000 167.920 ;
    END
  END sram_din0[23]
  PIN sram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 172.080 350.000 172.680 ;
    END
  END sram_din0[24]
  PIN sram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 176.840 350.000 177.440 ;
    END
  END sram_din0[25]
  PIN sram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 180.920 350.000 181.520 ;
    END
  END sram_din0[26]
  PIN sram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 185.680 350.000 186.280 ;
    END
  END sram_din0[27]
  PIN sram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 190.440 350.000 191.040 ;
    END
  END sram_din0[28]
  PIN sram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 194.520 350.000 195.120 ;
    END
  END sram_din0[29]
  PIN sram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 47.640 350.000 48.240 ;
    END
  END sram_din0[2]
  PIN sram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 199.280 350.000 199.880 ;
    END
  END sram_din0[30]
  PIN sram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.040 350.000 204.640 ;
    END
  END sram_din0[31]
  PIN sram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 59.880 350.000 60.480 ;
    END
  END sram_din0[3]
  PIN sram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 68.720 350.000 69.320 ;
    END
  END sram_din0[4]
  PIN sram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 76.200 350.000 76.800 ;
    END
  END sram_din0[5]
  PIN sram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 83.680 350.000 84.280 ;
    END
  END sram_din0[6]
  PIN sram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 91.840 350.000 92.440 ;
    END
  END sram_din0[7]
  PIN sram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 99.320 350.000 99.920 ;
    END
  END sram_din0[8]
  PIN sram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 103.400 350.000 104.000 ;
    END
  END sram_din0[9]
  PIN sram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 24.520 350.000 25.120 ;
    END
  END sram_dout0[0]
  PIN sram_dout0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 414.840 350.000 415.440 ;
    END
  END sram_dout0[100]
  PIN sram_dout0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 418.240 350.000 418.840 ;
    END
  END sram_dout0[101]
  PIN sram_dout0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 420.960 350.000 421.560 ;
    END
  END sram_dout0[102]
  PIN sram_dout0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 424.360 350.000 424.960 ;
    END
  END sram_dout0[103]
  PIN sram_dout0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 427.080 350.000 427.680 ;
    END
  END sram_dout0[104]
  PIN sram_dout0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 430.480 350.000 431.080 ;
    END
  END sram_dout0[105]
  PIN sram_dout0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 433.200 350.000 433.800 ;
    END
  END sram_dout0[106]
  PIN sram_dout0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 436.600 350.000 437.200 ;
    END
  END sram_dout0[107]
  PIN sram_dout0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 439.320 350.000 439.920 ;
    END
  END sram_dout0[108]
  PIN sram_dout0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 442.720 350.000 443.320 ;
    END
  END sram_dout0[109]
  PIN sram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 109.520 350.000 110.120 ;
    END
  END sram_dout0[10]
  PIN sram_dout0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 445.440 350.000 446.040 ;
    END
  END sram_dout0[110]
  PIN sram_dout0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 448.840 350.000 449.440 ;
    END
  END sram_dout0[111]
  PIN sram_dout0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 451.560 350.000 452.160 ;
    END
  END sram_dout0[112]
  PIN sram_dout0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 454.280 350.000 454.880 ;
    END
  END sram_dout0[113]
  PIN sram_dout0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 457.680 350.000 458.280 ;
    END
  END sram_dout0[114]
  PIN sram_dout0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 460.400 350.000 461.000 ;
    END
  END sram_dout0[115]
  PIN sram_dout0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 463.800 350.000 464.400 ;
    END
  END sram_dout0[116]
  PIN sram_dout0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 466.520 350.000 467.120 ;
    END
  END sram_dout0[117]
  PIN sram_dout0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 469.920 350.000 470.520 ;
    END
  END sram_dout0[118]
  PIN sram_dout0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 472.640 350.000 473.240 ;
    END
  END sram_dout0[119]
  PIN sram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 114.280 350.000 114.880 ;
    END
  END sram_dout0[11]
  PIN sram_dout0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 476.040 350.000 476.640 ;
    END
  END sram_dout0[120]
  PIN sram_dout0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 478.760 350.000 479.360 ;
    END
  END sram_dout0[121]
  PIN sram_dout0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 482.160 350.000 482.760 ;
    END
  END sram_dout0[122]
  PIN sram_dout0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 484.880 350.000 485.480 ;
    END
  END sram_dout0[123]
  PIN sram_dout0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 488.280 350.000 488.880 ;
    END
  END sram_dout0[124]
  PIN sram_dout0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 491.000 350.000 491.600 ;
    END
  END sram_dout0[125]
  PIN sram_dout0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 494.400 350.000 495.000 ;
    END
  END sram_dout0[126]
  PIN sram_dout0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 497.120 350.000 497.720 ;
    END
  END sram_dout0[127]
  PIN sram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 119.040 350.000 119.640 ;
    END
  END sram_dout0[12]
  PIN sram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 123.120 350.000 123.720 ;
    END
  END sram_dout0[13]
  PIN sram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 127.880 350.000 128.480 ;
    END
  END sram_dout0[14]
  PIN sram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 132.640 350.000 133.240 ;
    END
  END sram_dout0[15]
  PIN sram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 137.400 350.000 138.000 ;
    END
  END sram_dout0[16]
  PIN sram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 141.480 350.000 142.080 ;
    END
  END sram_dout0[17]
  PIN sram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 146.240 350.000 146.840 ;
    END
  END sram_dout0[18]
  PIN sram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 151.000 350.000 151.600 ;
    END
  END sram_dout0[19]
  PIN sram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 36.760 350.000 37.360 ;
    END
  END sram_dout0[1]
  PIN sram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 155.080 350.000 155.680 ;
    END
  END sram_dout0[20]
  PIN sram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 159.840 350.000 160.440 ;
    END
  END sram_dout0[21]
  PIN sram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 164.600 350.000 165.200 ;
    END
  END sram_dout0[22]
  PIN sram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 168.680 350.000 169.280 ;
    END
  END sram_dout0[23]
  PIN sram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 173.440 350.000 174.040 ;
    END
  END sram_dout0[24]
  PIN sram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 178.200 350.000 178.800 ;
    END
  END sram_dout0[25]
  PIN sram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 182.960 350.000 183.560 ;
    END
  END sram_dout0[26]
  PIN sram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 187.040 350.000 187.640 ;
    END
  END sram_dout0[27]
  PIN sram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 191.800 350.000 192.400 ;
    END
  END sram_dout0[28]
  PIN sram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 196.560 350.000 197.160 ;
    END
  END sram_dout0[29]
  PIN sram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 49.000 350.000 49.600 ;
    END
  END sram_dout0[2]
  PIN sram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 200.640 350.000 201.240 ;
    END
  END sram_dout0[30]
  PIN sram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 205.400 350.000 206.000 ;
    END
  END sram_dout0[31]
  PIN sram_dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 208.800 350.000 209.400 ;
    END
  END sram_dout0[32]
  PIN sram_dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 211.520 350.000 212.120 ;
    END
  END sram_dout0[33]
  PIN sram_dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 214.920 350.000 215.520 ;
    END
  END sram_dout0[34]
  PIN sram_dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 217.640 350.000 218.240 ;
    END
  END sram_dout0[35]
  PIN sram_dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 220.360 350.000 220.960 ;
    END
  END sram_dout0[36]
  PIN sram_dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 223.760 350.000 224.360 ;
    END
  END sram_dout0[37]
  PIN sram_dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 226.480 350.000 227.080 ;
    END
  END sram_dout0[38]
  PIN sram_dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 229.880 350.000 230.480 ;
    END
  END sram_dout0[39]
  PIN sram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 61.240 350.000 61.840 ;
    END
  END sram_dout0[3]
  PIN sram_dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 232.600 350.000 233.200 ;
    END
  END sram_dout0[40]
  PIN sram_dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 236.000 350.000 236.600 ;
    END
  END sram_dout0[41]
  PIN sram_dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 238.720 350.000 239.320 ;
    END
  END sram_dout0[42]
  PIN sram_dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 242.120 350.000 242.720 ;
    END
  END sram_dout0[43]
  PIN sram_dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 244.840 350.000 245.440 ;
    END
  END sram_dout0[44]
  PIN sram_dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 248.240 350.000 248.840 ;
    END
  END sram_dout0[45]
  PIN sram_dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 250.960 350.000 251.560 ;
    END
  END sram_dout0[46]
  PIN sram_dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 254.360 350.000 254.960 ;
    END
  END sram_dout0[47]
  PIN sram_dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 257.080 350.000 257.680 ;
    END
  END sram_dout0[48]
  PIN sram_dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 260.480 350.000 261.080 ;
    END
  END sram_dout0[49]
  PIN sram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 70.080 350.000 70.680 ;
    END
  END sram_dout0[4]
  PIN sram_dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 263.200 350.000 263.800 ;
    END
  END sram_dout0[50]
  PIN sram_dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 265.920 350.000 266.520 ;
    END
  END sram_dout0[51]
  PIN sram_dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 269.320 350.000 269.920 ;
    END
  END sram_dout0[52]
  PIN sram_dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 272.040 350.000 272.640 ;
    END
  END sram_dout0[53]
  PIN sram_dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 275.440 350.000 276.040 ;
    END
  END sram_dout0[54]
  PIN sram_dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 278.160 350.000 278.760 ;
    END
  END sram_dout0[55]
  PIN sram_dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 281.560 350.000 282.160 ;
    END
  END sram_dout0[56]
  PIN sram_dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 284.280 350.000 284.880 ;
    END
  END sram_dout0[57]
  PIN sram_dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 287.680 350.000 288.280 ;
    END
  END sram_dout0[58]
  PIN sram_dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 290.400 350.000 291.000 ;
    END
  END sram_dout0[59]
  PIN sram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 77.560 350.000 78.160 ;
    END
  END sram_dout0[5]
  PIN sram_dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 293.800 350.000 294.400 ;
    END
  END sram_dout0[60]
  PIN sram_dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 296.520 350.000 297.120 ;
    END
  END sram_dout0[61]
  PIN sram_dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 299.920 350.000 300.520 ;
    END
  END sram_dout0[62]
  PIN sram_dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 302.640 350.000 303.240 ;
    END
  END sram_dout0[63]
  PIN sram_dout0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 306.040 350.000 306.640 ;
    END
  END sram_dout0[64]
  PIN sram_dout0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 308.760 350.000 309.360 ;
    END
  END sram_dout0[65]
  PIN sram_dout0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 311.480 350.000 312.080 ;
    END
  END sram_dout0[66]
  PIN sram_dout0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 314.880 350.000 315.480 ;
    END
  END sram_dout0[67]
  PIN sram_dout0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 317.600 350.000 318.200 ;
    END
  END sram_dout0[68]
  PIN sram_dout0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 321.000 350.000 321.600 ;
    END
  END sram_dout0[69]
  PIN sram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 85.720 350.000 86.320 ;
    END
  END sram_dout0[6]
  PIN sram_dout0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 323.720 350.000 324.320 ;
    END
  END sram_dout0[70]
  PIN sram_dout0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 327.120 350.000 327.720 ;
    END
  END sram_dout0[71]
  PIN sram_dout0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 329.840 350.000 330.440 ;
    END
  END sram_dout0[72]
  PIN sram_dout0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 333.240 350.000 333.840 ;
    END
  END sram_dout0[73]
  PIN sram_dout0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.960 350.000 336.560 ;
    END
  END sram_dout0[74]
  PIN sram_dout0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 339.360 350.000 339.960 ;
    END
  END sram_dout0[75]
  PIN sram_dout0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 342.080 350.000 342.680 ;
    END
  END sram_dout0[76]
  PIN sram_dout0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 345.480 350.000 346.080 ;
    END
  END sram_dout0[77]
  PIN sram_dout0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 348.200 350.000 348.800 ;
    END
  END sram_dout0[78]
  PIN sram_dout0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 351.600 350.000 352.200 ;
    END
  END sram_dout0[79]
  PIN sram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 93.200 350.000 93.800 ;
    END
  END sram_dout0[7]
  PIN sram_dout0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 354.320 350.000 354.920 ;
    END
  END sram_dout0[80]
  PIN sram_dout0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 357.720 350.000 358.320 ;
    END
  END sram_dout0[81]
  PIN sram_dout0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 360.440 350.000 361.040 ;
    END
  END sram_dout0[82]
  PIN sram_dout0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 363.160 350.000 363.760 ;
    END
  END sram_dout0[83]
  PIN sram_dout0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 366.560 350.000 367.160 ;
    END
  END sram_dout0[84]
  PIN sram_dout0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 369.280 350.000 369.880 ;
    END
  END sram_dout0[85]
  PIN sram_dout0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 372.680 350.000 373.280 ;
    END
  END sram_dout0[86]
  PIN sram_dout0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 375.400 350.000 376.000 ;
    END
  END sram_dout0[87]
  PIN sram_dout0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 378.800 350.000 379.400 ;
    END
  END sram_dout0[88]
  PIN sram_dout0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 381.520 350.000 382.120 ;
    END
  END sram_dout0[89]
  PIN sram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 100.680 350.000 101.280 ;
    END
  END sram_dout0[8]
  PIN sram_dout0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 384.920 350.000 385.520 ;
    END
  END sram_dout0[90]
  PIN sram_dout0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 387.640 350.000 388.240 ;
    END
  END sram_dout0[91]
  PIN sram_dout0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 391.040 350.000 391.640 ;
    END
  END sram_dout0[92]
  PIN sram_dout0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 393.760 350.000 394.360 ;
    END
  END sram_dout0[93]
  PIN sram_dout0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 397.160 350.000 397.760 ;
    END
  END sram_dout0[94]
  PIN sram_dout0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 399.880 350.000 400.480 ;
    END
  END sram_dout0[95]
  PIN sram_dout0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 403.280 350.000 403.880 ;
    END
  END sram_dout0[96]
  PIN sram_dout0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 406.000 350.000 406.600 ;
    END
  END sram_dout0[97]
  PIN sram_dout0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 408.720 350.000 409.320 ;
    END
  END sram_dout0[98]
  PIN sram_dout0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 412.120 350.000 412.720 ;
    END
  END sram_dout0[99]
  PIN sram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 105.440 350.000 106.040 ;
    END
  END sram_dout0[9]
  PIN sram_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 25.880 350.000 26.480 ;
    END
  END sram_dout1[0]
  PIN sram_dout1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 416.880 350.000 417.480 ;
    END
  END sram_dout1[100]
  PIN sram_dout1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 419.600 350.000 420.200 ;
    END
  END sram_dout1[101]
  PIN sram_dout1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 423.000 350.000 423.600 ;
    END
  END sram_dout1[102]
  PIN sram_dout1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 425.720 350.000 426.320 ;
    END
  END sram_dout1[103]
  PIN sram_dout1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 429.120 350.000 429.720 ;
    END
  END sram_dout1[104]
  PIN sram_dout1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 431.840 350.000 432.440 ;
    END
  END sram_dout1[105]
  PIN sram_dout1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 434.560 350.000 435.160 ;
    END
  END sram_dout1[106]
  PIN sram_dout1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 437.960 350.000 438.560 ;
    END
  END sram_dout1[107]
  PIN sram_dout1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 440.680 350.000 441.280 ;
    END
  END sram_dout1[108]
  PIN sram_dout1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 444.080 350.000 444.680 ;
    END
  END sram_dout1[109]
  PIN sram_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 111.560 350.000 112.160 ;
    END
  END sram_dout1[10]
  PIN sram_dout1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 446.800 350.000 447.400 ;
    END
  END sram_dout1[110]
  PIN sram_dout1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 450.200 350.000 450.800 ;
    END
  END sram_dout1[111]
  PIN sram_dout1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 452.920 350.000 453.520 ;
    END
  END sram_dout1[112]
  PIN sram_dout1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 456.320 350.000 456.920 ;
    END
  END sram_dout1[113]
  PIN sram_dout1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 459.040 350.000 459.640 ;
    END
  END sram_dout1[114]
  PIN sram_dout1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 462.440 350.000 463.040 ;
    END
  END sram_dout1[115]
  PIN sram_dout1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 465.160 350.000 465.760 ;
    END
  END sram_dout1[116]
  PIN sram_dout1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 468.560 350.000 469.160 ;
    END
  END sram_dout1[117]
  PIN sram_dout1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 471.280 350.000 471.880 ;
    END
  END sram_dout1[118]
  PIN sram_dout1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 474.680 350.000 475.280 ;
    END
  END sram_dout1[119]
  PIN sram_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 115.640 350.000 116.240 ;
    END
  END sram_dout1[11]
  PIN sram_dout1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 477.400 350.000 478.000 ;
    END
  END sram_dout1[120]
  PIN sram_dout1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 480.120 350.000 480.720 ;
    END
  END sram_dout1[121]
  PIN sram_dout1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 483.520 350.000 484.120 ;
    END
  END sram_dout1[122]
  PIN sram_dout1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 486.240 350.000 486.840 ;
    END
  END sram_dout1[123]
  PIN sram_dout1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 489.640 350.000 490.240 ;
    END
  END sram_dout1[124]
  PIN sram_dout1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 492.360 350.000 492.960 ;
    END
  END sram_dout1[125]
  PIN sram_dout1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 495.760 350.000 496.360 ;
    END
  END sram_dout1[126]
  PIN sram_dout1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 498.480 350.000 499.080 ;
    END
  END sram_dout1[127]
  PIN sram_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 120.400 350.000 121.000 ;
    END
  END sram_dout1[12]
  PIN sram_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 125.160 350.000 125.760 ;
    END
  END sram_dout1[13]
  PIN sram_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 129.240 350.000 129.840 ;
    END
  END sram_dout1[14]
  PIN sram_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 134.000 350.000 134.600 ;
    END
  END sram_dout1[15]
  PIN sram_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 138.760 350.000 139.360 ;
    END
  END sram_dout1[16]
  PIN sram_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 143.520 350.000 144.120 ;
    END
  END sram_dout1[17]
  PIN sram_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 147.600 350.000 148.200 ;
    END
  END sram_dout1[18]
  PIN sram_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 152.360 350.000 152.960 ;
    END
  END sram_dout1[19]
  PIN sram_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 38.120 350.000 38.720 ;
    END
  END sram_dout1[1]
  PIN sram_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 157.120 350.000 157.720 ;
    END
  END sram_dout1[20]
  PIN sram_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 161.200 350.000 161.800 ;
    END
  END sram_dout1[21]
  PIN sram_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 165.960 350.000 166.560 ;
    END
  END sram_dout1[22]
  PIN sram_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 170.720 350.000 171.320 ;
    END
  END sram_dout1[23]
  PIN sram_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 174.800 350.000 175.400 ;
    END
  END sram_dout1[24]
  PIN sram_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 179.560 350.000 180.160 ;
    END
  END sram_dout1[25]
  PIN sram_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 184.320 350.000 184.920 ;
    END
  END sram_dout1[26]
  PIN sram_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 189.080 350.000 189.680 ;
    END
  END sram_dout1[27]
  PIN sram_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 193.160 350.000 193.760 ;
    END
  END sram_dout1[28]
  PIN sram_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 197.920 350.000 198.520 ;
    END
  END sram_dout1[29]
  PIN sram_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 50.360 350.000 50.960 ;
    END
  END sram_dout1[2]
  PIN sram_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 202.680 350.000 203.280 ;
    END
  END sram_dout1[30]
  PIN sram_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 206.760 350.000 207.360 ;
    END
  END sram_dout1[31]
  PIN sram_dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 210.160 350.000 210.760 ;
    END
  END sram_dout1[32]
  PIN sram_dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 212.880 350.000 213.480 ;
    END
  END sram_dout1[33]
  PIN sram_dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.280 350.000 216.880 ;
    END
  END sram_dout1[34]
  PIN sram_dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 219.000 350.000 219.600 ;
    END
  END sram_dout1[35]
  PIN sram_dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 222.400 350.000 223.000 ;
    END
  END sram_dout1[36]
  PIN sram_dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 225.120 350.000 225.720 ;
    END
  END sram_dout1[37]
  PIN sram_dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 228.520 350.000 229.120 ;
    END
  END sram_dout1[38]
  PIN sram_dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 231.240 350.000 231.840 ;
    END
  END sram_dout1[39]
  PIN sram_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 62.600 350.000 63.200 ;
    END
  END sram_dout1[3]
  PIN sram_dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 234.640 350.000 235.240 ;
    END
  END sram_dout1[40]
  PIN sram_dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 237.360 350.000 237.960 ;
    END
  END sram_dout1[41]
  PIN sram_dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 240.080 350.000 240.680 ;
    END
  END sram_dout1[42]
  PIN sram_dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.480 350.000 244.080 ;
    END
  END sram_dout1[43]
  PIN sram_dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 246.200 350.000 246.800 ;
    END
  END sram_dout1[44]
  PIN sram_dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 249.600 350.000 250.200 ;
    END
  END sram_dout1[45]
  PIN sram_dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 252.320 350.000 252.920 ;
    END
  END sram_dout1[46]
  PIN sram_dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 255.720 350.000 256.320 ;
    END
  END sram_dout1[47]
  PIN sram_dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 258.440 350.000 259.040 ;
    END
  END sram_dout1[48]
  PIN sram_dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 261.840 350.000 262.440 ;
    END
  END sram_dout1[49]
  PIN sram_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 72.120 350.000 72.720 ;
    END
  END sram_dout1[4]
  PIN sram_dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 264.560 350.000 265.160 ;
    END
  END sram_dout1[50]
  PIN sram_dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 267.960 350.000 268.560 ;
    END
  END sram_dout1[51]
  PIN sram_dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 270.680 350.000 271.280 ;
    END
  END sram_dout1[52]
  PIN sram_dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 274.080 350.000 274.680 ;
    END
  END sram_dout1[53]
  PIN sram_dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 276.800 350.000 277.400 ;
    END
  END sram_dout1[54]
  PIN sram_dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.200 350.000 280.800 ;
    END
  END sram_dout1[55]
  PIN sram_dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 282.920 350.000 283.520 ;
    END
  END sram_dout1[56]
  PIN sram_dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 286.320 350.000 286.920 ;
    END
  END sram_dout1[57]
  PIN sram_dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 289.040 350.000 289.640 ;
    END
  END sram_dout1[58]
  PIN sram_dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 291.760 350.000 292.360 ;
    END
  END sram_dout1[59]
  PIN sram_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 79.600 350.000 80.200 ;
    END
  END sram_dout1[5]
  PIN sram_dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 295.160 350.000 295.760 ;
    END
  END sram_dout1[60]
  PIN sram_dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 297.880 350.000 298.480 ;
    END
  END sram_dout1[61]
  PIN sram_dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 301.280 350.000 301.880 ;
    END
  END sram_dout1[62]
  PIN sram_dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 304.000 350.000 304.600 ;
    END
  END sram_dout1[63]
  PIN sram_dout1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 307.400 350.000 308.000 ;
    END
  END sram_dout1[64]
  PIN sram_dout1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 310.120 350.000 310.720 ;
    END
  END sram_dout1[65]
  PIN sram_dout1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 313.520 350.000 314.120 ;
    END
  END sram_dout1[66]
  PIN sram_dout1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 316.240 350.000 316.840 ;
    END
  END sram_dout1[67]
  PIN sram_dout1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 319.640 350.000 320.240 ;
    END
  END sram_dout1[68]
  PIN sram_dout1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 322.360 350.000 322.960 ;
    END
  END sram_dout1[69]
  PIN sram_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 87.080 350.000 87.680 ;
    END
  END sram_dout1[6]
  PIN sram_dout1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 325.760 350.000 326.360 ;
    END
  END sram_dout1[70]
  PIN sram_dout1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 328.480 350.000 329.080 ;
    END
  END sram_dout1[71]
  PIN sram_dout1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 331.880 350.000 332.480 ;
    END
  END sram_dout1[72]
  PIN sram_dout1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 334.600 350.000 335.200 ;
    END
  END sram_dout1[73]
  PIN sram_dout1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 337.320 350.000 337.920 ;
    END
  END sram_dout1[74]
  PIN sram_dout1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 340.720 350.000 341.320 ;
    END
  END sram_dout1[75]
  PIN sram_dout1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 343.440 350.000 344.040 ;
    END
  END sram_dout1[76]
  PIN sram_dout1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 346.840 350.000 347.440 ;
    END
  END sram_dout1[77]
  PIN sram_dout1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 349.560 350.000 350.160 ;
    END
  END sram_dout1[78]
  PIN sram_dout1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 352.960 350.000 353.560 ;
    END
  END sram_dout1[79]
  PIN sram_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 94.560 350.000 95.160 ;
    END
  END sram_dout1[7]
  PIN sram_dout1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 355.680 350.000 356.280 ;
    END
  END sram_dout1[80]
  PIN sram_dout1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 359.080 350.000 359.680 ;
    END
  END sram_dout1[81]
  PIN sram_dout1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 361.800 350.000 362.400 ;
    END
  END sram_dout1[82]
  PIN sram_dout1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 365.200 350.000 365.800 ;
    END
  END sram_dout1[83]
  PIN sram_dout1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 367.920 350.000 368.520 ;
    END
  END sram_dout1[84]
  PIN sram_dout1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 371.320 350.000 371.920 ;
    END
  END sram_dout1[85]
  PIN sram_dout1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 374.040 350.000 374.640 ;
    END
  END sram_dout1[86]
  PIN sram_dout1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 377.440 350.000 378.040 ;
    END
  END sram_dout1[87]
  PIN sram_dout1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 380.160 350.000 380.760 ;
    END
  END sram_dout1[88]
  PIN sram_dout1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 382.880 350.000 383.480 ;
    END
  END sram_dout1[89]
  PIN sram_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 102.040 350.000 102.640 ;
    END
  END sram_dout1[8]
  PIN sram_dout1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 386.280 350.000 386.880 ;
    END
  END sram_dout1[90]
  PIN sram_dout1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 389.000 350.000 389.600 ;
    END
  END sram_dout1[91]
  PIN sram_dout1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 392.400 350.000 393.000 ;
    END
  END sram_dout1[92]
  PIN sram_dout1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 395.120 350.000 395.720 ;
    END
  END sram_dout1[93]
  PIN sram_dout1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 398.520 350.000 399.120 ;
    END
  END sram_dout1[94]
  PIN sram_dout1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 401.240 350.000 401.840 ;
    END
  END sram_dout1[95]
  PIN sram_dout1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 404.640 350.000 405.240 ;
    END
  END sram_dout1[96]
  PIN sram_dout1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 407.360 350.000 407.960 ;
    END
  END sram_dout1[97]
  PIN sram_dout1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 410.760 350.000 411.360 ;
    END
  END sram_dout1[98]
  PIN sram_dout1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 413.480 350.000 414.080 ;
    END
  END sram_dout1[99]
  PIN sram_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 106.800 350.000 107.400 ;
    END
  END sram_dout1[9]
  PIN sram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 15.680 350.000 16.280 ;
    END
  END sram_web0
  PIN sram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 27.920 350.000 28.520 ;
    END
  END sram_wmask0[0]
  PIN sram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.160 350.000 40.760 ;
    END
  END sram_wmask0[1]
  PIN sram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 51.720 350.000 52.320 ;
    END
  END sram_wmask0[2]
  PIN sram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 63.960 350.000 64.560 ;
    END
  END sram_wmask0[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 3.440 350.000 4.040 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 8.200 350.000 8.800 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 4.800 350.000 5.400 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 9.560 350.000 10.160 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 0.720 350.000 1.320 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 6.160 350.000 6.760 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 10.920 350.000 11.520 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 2.080 350.000 2.680 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 486.965 ;
      LAYER met1 ;
        RECT 0.070 2.420 349.990 487.120 ;
      LAYER met2 ;
        RECT 0.100 4.280 349.960 497.605 ;
        RECT 0.100 0.835 1.190 4.280 ;
        RECT 2.030 0.835 4.410 4.280 ;
        RECT 5.250 0.835 8.090 4.280 ;
        RECT 8.930 0.835 11.310 4.280 ;
        RECT 12.150 0.835 14.990 4.280 ;
        RECT 15.830 0.835 18.670 4.280 ;
        RECT 19.510 0.835 21.890 4.280 ;
        RECT 22.730 0.835 25.570 4.280 ;
        RECT 26.410 0.835 28.790 4.280 ;
        RECT 29.630 0.835 32.470 4.280 ;
        RECT 33.310 0.835 36.150 4.280 ;
        RECT 36.990 0.835 39.370 4.280 ;
        RECT 40.210 0.835 43.050 4.280 ;
        RECT 43.890 0.835 46.270 4.280 ;
        RECT 47.110 0.835 49.950 4.280 ;
        RECT 50.790 0.835 53.630 4.280 ;
        RECT 54.470 0.835 56.850 4.280 ;
        RECT 57.690 0.835 60.530 4.280 ;
        RECT 61.370 0.835 63.750 4.280 ;
        RECT 64.590 0.835 67.430 4.280 ;
        RECT 68.270 0.835 71.110 4.280 ;
        RECT 71.950 0.835 74.330 4.280 ;
        RECT 75.170 0.835 78.010 4.280 ;
        RECT 78.850 0.835 81.690 4.280 ;
        RECT 82.530 0.835 84.910 4.280 ;
        RECT 85.750 0.835 88.590 4.280 ;
        RECT 89.430 0.835 91.810 4.280 ;
        RECT 92.650 0.835 95.490 4.280 ;
        RECT 96.330 0.835 99.170 4.280 ;
        RECT 100.010 0.835 102.390 4.280 ;
        RECT 103.230 0.835 106.070 4.280 ;
        RECT 106.910 0.835 109.290 4.280 ;
        RECT 110.130 0.835 112.970 4.280 ;
        RECT 113.810 0.835 116.650 4.280 ;
        RECT 117.490 0.835 119.870 4.280 ;
        RECT 120.710 0.835 123.550 4.280 ;
        RECT 124.390 0.835 126.770 4.280 ;
        RECT 127.610 0.835 130.450 4.280 ;
        RECT 131.290 0.835 134.130 4.280 ;
        RECT 134.970 0.835 137.350 4.280 ;
        RECT 138.190 0.835 141.030 4.280 ;
        RECT 141.870 0.835 144.710 4.280 ;
        RECT 145.550 0.835 147.930 4.280 ;
        RECT 148.770 0.835 151.610 4.280 ;
        RECT 152.450 0.835 154.830 4.280 ;
        RECT 155.670 0.835 158.510 4.280 ;
        RECT 159.350 0.835 162.190 4.280 ;
        RECT 163.030 0.835 165.410 4.280 ;
        RECT 166.250 0.835 169.090 4.280 ;
        RECT 169.930 0.835 172.310 4.280 ;
        RECT 173.150 0.835 175.990 4.280 ;
        RECT 176.830 0.835 179.670 4.280 ;
        RECT 180.510 0.835 182.890 4.280 ;
        RECT 183.730 0.835 186.570 4.280 ;
        RECT 187.410 0.835 189.790 4.280 ;
        RECT 190.630 0.835 193.470 4.280 ;
        RECT 194.310 0.835 197.150 4.280 ;
        RECT 197.990 0.835 200.370 4.280 ;
        RECT 201.210 0.835 204.050 4.280 ;
        RECT 204.890 0.835 207.270 4.280 ;
        RECT 208.110 0.835 210.950 4.280 ;
        RECT 211.790 0.835 214.630 4.280 ;
        RECT 215.470 0.835 217.850 4.280 ;
        RECT 218.690 0.835 221.530 4.280 ;
        RECT 222.370 0.835 225.210 4.280 ;
        RECT 226.050 0.835 228.430 4.280 ;
        RECT 229.270 0.835 232.110 4.280 ;
        RECT 232.950 0.835 235.330 4.280 ;
        RECT 236.170 0.835 239.010 4.280 ;
        RECT 239.850 0.835 242.690 4.280 ;
        RECT 243.530 0.835 245.910 4.280 ;
        RECT 246.750 0.835 249.590 4.280 ;
        RECT 250.430 0.835 252.810 4.280 ;
        RECT 253.650 0.835 256.490 4.280 ;
        RECT 257.330 0.835 260.170 4.280 ;
        RECT 261.010 0.835 263.390 4.280 ;
        RECT 264.230 0.835 267.070 4.280 ;
        RECT 267.910 0.835 270.290 4.280 ;
        RECT 271.130 0.835 273.970 4.280 ;
        RECT 274.810 0.835 277.650 4.280 ;
        RECT 278.490 0.835 280.870 4.280 ;
        RECT 281.710 0.835 284.550 4.280 ;
        RECT 285.390 0.835 288.230 4.280 ;
        RECT 289.070 0.835 291.450 4.280 ;
        RECT 292.290 0.835 295.130 4.280 ;
        RECT 295.970 0.835 298.350 4.280 ;
        RECT 299.190 0.835 302.030 4.280 ;
        RECT 302.870 0.835 305.710 4.280 ;
        RECT 306.550 0.835 308.930 4.280 ;
        RECT 309.770 0.835 312.610 4.280 ;
        RECT 313.450 0.835 315.830 4.280 ;
        RECT 316.670 0.835 319.510 4.280 ;
        RECT 320.350 0.835 323.190 4.280 ;
        RECT 324.030 0.835 326.410 4.280 ;
        RECT 327.250 0.835 330.090 4.280 ;
        RECT 330.930 0.835 333.310 4.280 ;
        RECT 334.150 0.835 336.990 4.280 ;
        RECT 337.830 0.835 340.670 4.280 ;
        RECT 341.510 0.835 343.890 4.280 ;
        RECT 344.730 0.835 347.570 4.280 ;
        RECT 348.410 0.835 349.960 4.280 ;
      LAYER met3 ;
        RECT 21.050 494.000 345.600 497.585 ;
        RECT 21.050 493.360 349.530 494.000 ;
        RECT 21.050 487.880 345.600 493.360 ;
        RECT 21.050 487.240 349.530 487.880 ;
        RECT 21.050 481.760 345.600 487.240 ;
        RECT 21.050 481.120 349.530 481.760 ;
        RECT 21.050 474.280 345.600 481.120 ;
        RECT 21.050 473.640 349.530 474.280 ;
        RECT 21.050 468.160 345.600 473.640 ;
        RECT 21.050 467.520 349.530 468.160 ;
        RECT 21.050 462.040 345.600 467.520 ;
        RECT 21.050 461.400 349.530 462.040 ;
        RECT 21.050 455.920 345.600 461.400 ;
        RECT 21.050 455.280 349.530 455.920 ;
        RECT 21.050 448.440 345.600 455.280 ;
        RECT 21.050 447.800 349.530 448.440 ;
        RECT 21.050 442.320 345.600 447.800 ;
        RECT 21.050 441.680 349.530 442.320 ;
        RECT 21.050 436.200 345.600 441.680 ;
        RECT 21.050 435.560 349.530 436.200 ;
        RECT 21.050 428.720 345.600 435.560 ;
        RECT 21.050 428.080 349.530 428.720 ;
        RECT 21.050 422.600 345.600 428.080 ;
        RECT 21.050 421.960 349.530 422.600 ;
        RECT 21.050 416.480 345.600 421.960 ;
        RECT 21.050 415.840 349.530 416.480 ;
        RECT 21.050 410.360 345.600 415.840 ;
        RECT 21.050 409.720 349.530 410.360 ;
        RECT 21.050 402.880 345.600 409.720 ;
        RECT 21.050 402.240 349.530 402.880 ;
        RECT 21.050 396.760 345.600 402.240 ;
        RECT 21.050 396.120 349.530 396.760 ;
        RECT 21.050 390.640 345.600 396.120 ;
        RECT 21.050 390.000 349.530 390.640 ;
        RECT 21.050 384.520 345.600 390.000 ;
        RECT 21.050 383.880 349.530 384.520 ;
        RECT 21.050 377.040 345.600 383.880 ;
        RECT 21.050 376.400 349.530 377.040 ;
        RECT 21.050 370.920 345.600 376.400 ;
        RECT 21.050 370.280 349.530 370.920 ;
        RECT 21.050 364.800 345.600 370.280 ;
        RECT 21.050 364.160 349.530 364.800 ;
        RECT 21.050 357.320 345.600 364.160 ;
        RECT 21.050 356.680 349.530 357.320 ;
        RECT 21.050 351.200 345.600 356.680 ;
        RECT 21.050 350.560 349.530 351.200 ;
        RECT 21.050 345.080 345.600 350.560 ;
        RECT 21.050 344.440 349.530 345.080 ;
        RECT 21.050 338.960 345.600 344.440 ;
        RECT 21.050 338.320 349.530 338.960 ;
        RECT 21.050 331.480 345.600 338.320 ;
        RECT 21.050 330.840 349.530 331.480 ;
        RECT 21.050 325.360 345.600 330.840 ;
        RECT 21.050 324.720 349.530 325.360 ;
        RECT 21.050 319.240 345.600 324.720 ;
        RECT 21.050 318.600 349.530 319.240 ;
        RECT 21.050 313.120 345.600 318.600 ;
        RECT 21.050 312.480 349.530 313.120 ;
        RECT 21.050 305.640 345.600 312.480 ;
        RECT 21.050 305.000 349.530 305.640 ;
        RECT 21.050 299.520 345.600 305.000 ;
        RECT 21.050 298.880 349.530 299.520 ;
        RECT 21.050 293.400 345.600 298.880 ;
        RECT 21.050 292.760 349.530 293.400 ;
        RECT 21.050 285.920 345.600 292.760 ;
        RECT 21.050 285.280 349.530 285.920 ;
        RECT 21.050 279.800 345.600 285.280 ;
        RECT 21.050 279.160 349.530 279.800 ;
        RECT 21.050 273.680 345.600 279.160 ;
        RECT 21.050 273.040 349.530 273.680 ;
        RECT 21.050 267.560 345.600 273.040 ;
        RECT 21.050 266.920 349.530 267.560 ;
        RECT 21.050 260.080 345.600 266.920 ;
        RECT 21.050 259.440 349.530 260.080 ;
        RECT 21.050 253.960 345.600 259.440 ;
        RECT 21.050 253.320 349.530 253.960 ;
        RECT 21.050 247.840 345.600 253.320 ;
        RECT 21.050 247.200 349.530 247.840 ;
        RECT 21.050 241.720 345.600 247.200 ;
        RECT 21.050 241.080 349.530 241.720 ;
        RECT 21.050 234.240 345.600 241.080 ;
        RECT 21.050 233.600 349.530 234.240 ;
        RECT 21.050 228.120 345.600 233.600 ;
        RECT 21.050 227.480 349.530 228.120 ;
        RECT 21.050 222.000 345.600 227.480 ;
        RECT 21.050 221.360 349.530 222.000 ;
        RECT 21.050 214.520 345.600 221.360 ;
        RECT 21.050 213.880 349.530 214.520 ;
        RECT 21.050 208.400 345.600 213.880 ;
        RECT 21.050 207.760 349.530 208.400 ;
        RECT 21.050 202.280 345.600 207.760 ;
        RECT 21.050 201.640 349.530 202.280 ;
        RECT 21.050 196.160 345.600 201.640 ;
        RECT 21.050 195.520 349.530 196.160 ;
        RECT 21.050 188.680 345.600 195.520 ;
        RECT 21.050 188.040 349.530 188.680 ;
        RECT 21.050 182.560 345.600 188.040 ;
        RECT 21.050 181.920 349.530 182.560 ;
        RECT 21.050 176.440 345.600 181.920 ;
        RECT 21.050 175.800 349.530 176.440 ;
        RECT 21.050 170.320 345.600 175.800 ;
        RECT 21.050 169.680 349.530 170.320 ;
        RECT 21.050 162.840 345.600 169.680 ;
        RECT 21.050 162.200 349.530 162.840 ;
        RECT 21.050 156.720 345.600 162.200 ;
        RECT 21.050 156.080 349.530 156.720 ;
        RECT 21.050 150.600 345.600 156.080 ;
        RECT 21.050 149.960 349.530 150.600 ;
        RECT 21.050 143.120 345.600 149.960 ;
        RECT 21.050 142.480 349.530 143.120 ;
        RECT 21.050 137.000 345.600 142.480 ;
        RECT 21.050 136.360 349.530 137.000 ;
        RECT 21.050 130.880 345.600 136.360 ;
        RECT 21.050 130.240 349.530 130.880 ;
        RECT 21.050 124.760 345.600 130.240 ;
        RECT 21.050 124.120 349.530 124.760 ;
        RECT 21.050 117.280 345.600 124.120 ;
        RECT 21.050 116.640 349.530 117.280 ;
        RECT 21.050 111.160 345.600 116.640 ;
        RECT 21.050 110.520 349.530 111.160 ;
        RECT 21.050 105.040 345.600 110.520 ;
        RECT 21.050 104.400 349.530 105.040 ;
        RECT 21.050 98.920 345.600 104.400 ;
        RECT 21.050 98.280 349.530 98.920 ;
        RECT 21.050 91.440 345.600 98.280 ;
        RECT 21.050 90.800 349.530 91.440 ;
        RECT 21.050 85.320 345.600 90.800 ;
        RECT 21.050 84.680 349.530 85.320 ;
        RECT 21.050 79.200 345.600 84.680 ;
        RECT 21.050 78.560 349.530 79.200 ;
        RECT 21.050 71.720 345.600 78.560 ;
        RECT 21.050 71.080 349.530 71.720 ;
        RECT 21.050 65.600 345.600 71.080 ;
        RECT 21.050 64.960 349.530 65.600 ;
        RECT 21.050 59.480 345.600 64.960 ;
        RECT 21.050 58.840 349.530 59.480 ;
        RECT 21.050 53.360 345.600 58.840 ;
        RECT 21.050 52.720 349.530 53.360 ;
        RECT 21.050 45.880 345.600 52.720 ;
        RECT 21.050 45.240 349.530 45.880 ;
        RECT 21.050 39.760 345.600 45.240 ;
        RECT 21.050 39.120 349.530 39.760 ;
        RECT 21.050 33.640 345.600 39.120 ;
        RECT 21.050 33.000 349.530 33.640 ;
        RECT 21.050 27.520 345.600 33.000 ;
        RECT 21.050 26.880 349.530 27.520 ;
        RECT 21.050 20.040 345.600 26.880 ;
        RECT 21.050 19.400 349.530 20.040 ;
        RECT 21.050 13.920 345.600 19.400 ;
        RECT 21.050 13.280 349.530 13.920 ;
        RECT 21.050 7.800 345.600 13.280 ;
        RECT 21.050 7.160 349.530 7.800 ;
        RECT 21.050 0.855 345.600 7.160 ;
      LAYER met4 ;
        RECT 281.815 13.095 327.840 483.305 ;
        RECT 330.240 13.095 349.305 483.305 ;
  END
END Video
END LIBRARY

