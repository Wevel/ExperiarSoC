magic
tech sky130A
magscale 1 2
timestamp 1651490877
<< viali >>
rect 6377 37417 6411 37451
rect 6929 37349 6963 37383
rect 2053 37281 2087 37315
rect 2789 37281 2823 37315
rect 5273 37281 5307 37315
rect 37289 37281 37323 37315
rect 1869 37213 1903 37247
rect 3893 37213 3927 37247
rect 4537 37213 4571 37247
rect 33885 37213 33919 37247
rect 34989 37213 35023 37247
rect 35725 37213 35759 37247
rect 36461 37213 36495 37247
rect 37565 37213 37599 37247
rect 2605 37145 2639 37179
rect 4077 37145 4111 37179
rect 4721 37077 4755 37111
rect 34069 37077 34103 37111
rect 35173 37077 35207 37111
rect 35909 37077 35943 37111
rect 36645 37077 36679 37111
rect 3341 36873 3375 36907
rect 5273 36873 5307 36907
rect 29745 36873 29779 36907
rect 35265 36873 35299 36907
rect 1869 36805 1903 36839
rect 4721 36805 4755 36839
rect 2789 36737 2823 36771
rect 3525 36737 3559 36771
rect 3985 36737 4019 36771
rect 24593 36737 24627 36771
rect 33977 36737 34011 36771
rect 34437 36737 34471 36771
rect 35081 36737 35115 36771
rect 36001 36737 36035 36771
rect 37289 36737 37323 36771
rect 37565 36737 37599 36771
rect 2053 36669 2087 36703
rect 24409 36669 24443 36703
rect 35817 36669 35851 36703
rect 23857 36601 23891 36635
rect 34621 36601 34655 36635
rect 2605 36533 2639 36567
rect 4169 36533 4203 36567
rect 24777 36533 24811 36567
rect 25329 36533 25363 36567
rect 30665 36533 30699 36567
rect 36185 36533 36219 36567
rect 3801 36329 3835 36363
rect 5181 36329 5215 36363
rect 33793 36329 33827 36363
rect 36185 36329 36219 36363
rect 36829 36329 36863 36363
rect 2053 36261 2087 36295
rect 24501 36261 24535 36295
rect 26157 36261 26191 36295
rect 35357 36261 35391 36295
rect 20821 36193 20855 36227
rect 21649 36193 21683 36227
rect 25053 36193 25087 36227
rect 25421 36193 25455 36227
rect 29929 36193 29963 36227
rect 30297 36193 30331 36227
rect 31125 36193 31159 36227
rect 35817 36193 35851 36227
rect 37289 36193 37323 36227
rect 2789 36125 2823 36159
rect 3985 36125 4019 36159
rect 4629 36125 4663 36159
rect 20637 36125 20671 36159
rect 21465 36125 21499 36159
rect 22293 36125 22327 36159
rect 22477 36125 22511 36159
rect 25237 36125 25271 36159
rect 25973 36125 26007 36159
rect 26617 36125 26651 36159
rect 30113 36125 30147 36159
rect 30757 36125 30791 36159
rect 30941 36125 30975 36159
rect 32965 36125 32999 36159
rect 33609 36125 33643 36159
rect 35173 36125 35207 36159
rect 36001 36125 36035 36159
rect 37565 36125 37599 36159
rect 1869 36057 1903 36091
rect 22937 36057 22971 36091
rect 2605 35989 2639 36023
rect 4445 35989 4479 36023
rect 20453 35989 20487 36023
rect 21281 35989 21315 36023
rect 22109 35989 22143 36023
rect 26801 35989 26835 36023
rect 33149 35989 33183 36023
rect 2973 35785 3007 35819
rect 3617 35785 3651 35819
rect 4445 35785 4479 35819
rect 21005 35785 21039 35819
rect 21833 35785 21867 35819
rect 24869 35785 24903 35819
rect 26341 35785 26375 35819
rect 35541 35785 35575 35819
rect 4997 35717 5031 35751
rect 1869 35649 1903 35683
rect 3157 35649 3191 35683
rect 3801 35649 3835 35683
rect 4261 35649 4295 35683
rect 24685 35649 24719 35683
rect 26157 35649 26191 35683
rect 30113 35649 30147 35683
rect 30297 35649 30331 35683
rect 32873 35649 32907 35683
rect 36369 35649 36403 35683
rect 37841 35649 37875 35683
rect 23949 35581 23983 35615
rect 24501 35581 24535 35615
rect 29929 35581 29963 35615
rect 36553 35581 36587 35615
rect 2053 35513 2087 35547
rect 29377 35513 29411 35547
rect 33057 35513 33091 35547
rect 25513 35445 25547 35479
rect 36185 35445 36219 35479
rect 37289 35445 37323 35479
rect 38025 35445 38059 35479
rect 2973 35241 3007 35275
rect 3985 35241 4019 35275
rect 36553 35241 36587 35275
rect 35541 35173 35575 35207
rect 1685 35037 1719 35071
rect 2421 35037 2455 35071
rect 3157 35037 3191 35071
rect 3801 35037 3835 35071
rect 36093 35037 36127 35071
rect 36737 35037 36771 35071
rect 37381 35037 37415 35071
rect 37841 35037 37875 35071
rect 1501 34901 1535 34935
rect 2237 34901 2271 34935
rect 4537 34901 4571 34935
rect 25053 34901 25087 34935
rect 37197 34901 37231 34935
rect 38025 34901 38059 34935
rect 2697 34697 2731 34731
rect 3985 34697 4019 34731
rect 37657 34697 37691 34731
rect 2053 34629 2087 34663
rect 29285 34629 29319 34663
rect 36737 34629 36771 34663
rect 1869 34561 1903 34595
rect 2881 34561 2915 34595
rect 3433 34561 3467 34595
rect 29837 34561 29871 34595
rect 30021 34561 30055 34595
rect 30205 34561 30239 34595
rect 32137 34561 32171 34595
rect 37289 34561 37323 34595
rect 37473 34561 37507 34595
rect 32321 34425 32355 34459
rect 3065 34153 3099 34187
rect 37197 34085 37231 34119
rect 35449 34017 35483 34051
rect 2053 33949 2087 33983
rect 35265 33949 35299 33983
rect 36737 33949 36771 33983
rect 37381 33949 37415 33983
rect 37841 33949 37875 33983
rect 1869 33881 1903 33915
rect 2513 33881 2547 33915
rect 34069 33881 34103 33915
rect 35081 33881 35115 33915
rect 33977 33813 34011 33847
rect 38025 33813 38059 33847
rect 2145 33609 2179 33643
rect 29285 33609 29319 33643
rect 32321 33609 32355 33643
rect 1685 33473 1719 33507
rect 29837 33473 29871 33507
rect 30021 33473 30055 33507
rect 30205 33473 30239 33507
rect 32137 33473 32171 33507
rect 37841 33473 37875 33507
rect 37381 33337 37415 33371
rect 1501 33269 1535 33303
rect 38025 33269 38059 33303
rect 35449 33065 35483 33099
rect 37933 32997 37967 33031
rect 2513 32861 2547 32895
rect 3157 32861 3191 32895
rect 26985 32861 27019 32895
rect 35265 32861 35299 32895
rect 36829 32861 36863 32895
rect 37473 32861 37507 32895
rect 38117 32861 38151 32895
rect 1869 32793 1903 32827
rect 1961 32725 1995 32759
rect 2697 32725 2731 32759
rect 27169 32725 27203 32759
rect 35909 32725 35943 32759
rect 37289 32725 37323 32759
rect 25145 32521 25179 32555
rect 26065 32521 26099 32555
rect 29285 32521 29319 32555
rect 2145 32453 2179 32487
rect 1685 32385 1719 32419
rect 2881 32385 2915 32419
rect 25697 32385 25731 32419
rect 25881 32385 25915 32419
rect 29101 32385 29135 32419
rect 29745 32385 29779 32419
rect 37289 32385 37323 32419
rect 37473 32385 37507 32419
rect 2697 32249 2731 32283
rect 3433 32249 3467 32283
rect 37657 32249 37691 32283
rect 1501 32181 1535 32215
rect 1961 31977 1995 32011
rect 33793 31977 33827 32011
rect 38025 31977 38059 32011
rect 3157 31909 3191 31943
rect 25421 31909 25455 31943
rect 37289 31909 37323 31943
rect 23213 31841 23247 31875
rect 1869 31773 1903 31807
rect 2513 31773 2547 31807
rect 7665 31773 7699 31807
rect 11989 31773 12023 31807
rect 16589 31773 16623 31807
rect 18429 31773 18463 31807
rect 21465 31773 21499 31807
rect 21649 31773 21683 31807
rect 21833 31773 21867 31807
rect 22937 31773 22971 31807
rect 25973 31773 26007 31807
rect 26157 31773 26191 31807
rect 26341 31773 26375 31807
rect 27537 31773 27571 31807
rect 33885 31773 33919 31807
rect 37105 31773 37139 31807
rect 37841 31773 37875 31807
rect 16856 31705 16890 31739
rect 7481 31637 7515 31671
rect 11805 31637 11839 31671
rect 17969 31637 18003 31671
rect 21005 31637 21039 31671
rect 27721 31637 27755 31671
rect 2329 31433 2363 31467
rect 7389 31433 7423 31467
rect 16865 31433 16899 31467
rect 26985 31433 27019 31467
rect 35909 31433 35943 31467
rect 1685 31297 1719 31331
rect 2145 31297 2179 31331
rect 2789 31297 2823 31331
rect 7757 31297 7791 31331
rect 11888 31297 11922 31331
rect 16681 31297 16715 31331
rect 22017 31297 22051 31331
rect 27169 31297 27203 31331
rect 36093 31297 36127 31331
rect 37841 31297 37875 31331
rect 7849 31229 7883 31263
rect 8033 31229 8067 31263
rect 8585 31229 8619 31263
rect 10977 31229 11011 31263
rect 11621 31229 11655 31263
rect 21833 31229 21867 31263
rect 22201 31229 22235 31263
rect 23121 31229 23155 31263
rect 23397 31229 23431 31263
rect 36277 31229 36311 31263
rect 13001 31161 13035 31195
rect 1501 31093 1535 31127
rect 3433 31093 3467 31127
rect 21189 31093 21223 31127
rect 27721 31093 27755 31127
rect 38025 31093 38059 31127
rect 9045 30889 9079 30923
rect 11897 30889 11931 30923
rect 33793 30889 33827 30923
rect 35817 30889 35851 30923
rect 16497 30821 16531 30855
rect 7021 30753 7055 30787
rect 12357 30753 12391 30787
rect 12541 30753 12575 30787
rect 15853 30753 15887 30787
rect 21465 30753 21499 30787
rect 7288 30685 7322 30719
rect 12265 30685 12299 30719
rect 21649 30685 21683 30719
rect 35633 30685 35667 30719
rect 36277 30685 36311 30719
rect 37381 30685 37415 30719
rect 37841 30685 37875 30719
rect 1869 30617 1903 30651
rect 2513 30617 2547 30651
rect 16129 30617 16163 30651
rect 33885 30617 33919 30651
rect 1961 30549 1995 30583
rect 8401 30549 8435 30583
rect 16037 30549 16071 30583
rect 21005 30549 21039 30583
rect 21833 30549 21867 30583
rect 37197 30549 37231 30583
rect 38025 30549 38059 30583
rect 36185 30277 36219 30311
rect 1961 30209 1995 30243
rect 23121 30209 23155 30243
rect 23397 30209 23431 30243
rect 27169 30209 27203 30243
rect 27353 30209 27387 30243
rect 28089 30209 28123 30243
rect 36369 30209 36403 30243
rect 36553 30209 36587 30243
rect 37841 30209 37875 30243
rect 2237 30141 2271 30175
rect 2697 30141 2731 30175
rect 26433 30141 26467 30175
rect 26985 30141 27019 30175
rect 28273 30073 28307 30107
rect 3341 30005 3375 30039
rect 37381 30005 37415 30039
rect 38025 30005 38059 30039
rect 2053 29665 2087 29699
rect 2789 29597 2823 29631
rect 36737 29597 36771 29631
rect 37197 29597 37231 29631
rect 37841 29597 37875 29631
rect 1869 29529 1903 29563
rect 2605 29461 2639 29495
rect 37381 29461 37415 29495
rect 38025 29461 38059 29495
rect 26341 29257 26375 29291
rect 35449 29257 35483 29291
rect 3249 29189 3283 29223
rect 1961 29121 1995 29155
rect 26985 29121 27019 29155
rect 27169 29121 27203 29155
rect 27353 29121 27387 29155
rect 27997 29121 28031 29155
rect 35633 29121 35667 29155
rect 37289 29121 37323 29155
rect 37473 29121 37507 29155
rect 37565 29121 37599 29155
rect 2237 29053 2271 29087
rect 2697 29053 2731 29087
rect 28181 28985 28215 29019
rect 23259 28713 23293 28747
rect 16773 28645 16807 28679
rect 25881 28645 25915 28679
rect 16129 28577 16163 28611
rect 16313 28577 16347 28611
rect 21005 28577 21039 28611
rect 1685 28509 1719 28543
rect 17233 28509 17267 28543
rect 21465 28509 21499 28543
rect 21649 28509 21683 28543
rect 21833 28509 21867 28543
rect 23029 28509 23063 28543
rect 26433 28509 26467 28543
rect 26617 28509 26651 28543
rect 36737 28509 36771 28543
rect 37197 28509 37231 28543
rect 37841 28509 37875 28543
rect 2789 28441 2823 28475
rect 1501 28373 1535 28407
rect 2145 28373 2179 28407
rect 16405 28373 16439 28407
rect 17417 28373 17451 28407
rect 26801 28373 26835 28407
rect 37381 28373 37415 28407
rect 38025 28373 38059 28407
rect 17417 28169 17451 28203
rect 35817 28169 35851 28203
rect 2053 28101 2087 28135
rect 18236 28101 18270 28135
rect 1869 28033 1903 28067
rect 2513 28033 2547 28067
rect 3157 28033 3191 28067
rect 17969 28033 18003 28067
rect 27905 28033 27939 28067
rect 36001 28033 36035 28067
rect 37289 28033 37323 28067
rect 37473 28033 37507 28067
rect 37565 28033 37599 28067
rect 28089 27897 28123 27931
rect 2697 27829 2731 27863
rect 19349 27829 19383 27863
rect 9045 27557 9079 27591
rect 37289 27557 37323 27591
rect 1685 27421 1719 27455
rect 7021 27421 7055 27455
rect 11897 27421 11931 27455
rect 37105 27421 37139 27455
rect 37841 27421 37875 27455
rect 7266 27353 7300 27387
rect 1501 27285 1535 27319
rect 2145 27285 2179 27319
rect 2789 27285 2823 27319
rect 8401 27285 8435 27319
rect 12081 27285 12115 27319
rect 38025 27285 38059 27319
rect 12072 27013 12106 27047
rect 1961 26945 1995 26979
rect 25605 26945 25639 26979
rect 37841 26945 37875 26979
rect 2237 26877 2271 26911
rect 2697 26877 2731 26911
rect 10977 26877 11011 26911
rect 11805 26877 11839 26911
rect 3249 26741 3283 26775
rect 13185 26741 13219 26775
rect 25789 26741 25823 26775
rect 38025 26741 38059 26775
rect 7113 26537 7147 26571
rect 11989 26537 12023 26571
rect 29009 26537 29043 26571
rect 31309 26537 31343 26571
rect 35081 26537 35115 26571
rect 2605 26469 2639 26503
rect 23857 26469 23891 26503
rect 2053 26401 2087 26435
rect 12449 26401 12483 26435
rect 12633 26401 12667 26435
rect 23489 26401 23523 26435
rect 29561 26401 29595 26435
rect 1869 26333 1903 26367
rect 2789 26333 2823 26367
rect 3801 26333 3835 26367
rect 6929 26333 6963 26367
rect 12357 26333 12391 26367
rect 23673 26333 23707 26367
rect 29745 26333 29779 26367
rect 29929 26333 29963 26367
rect 31125 26333 31159 26367
rect 35265 26333 35299 26367
rect 37473 26333 37507 26367
rect 38117 26333 38151 26367
rect 37933 26197 37967 26231
rect 16957 25993 16991 26027
rect 27169 25993 27203 26027
rect 36185 25993 36219 26027
rect 1869 25925 1903 25959
rect 2053 25925 2087 25959
rect 2964 25857 2998 25891
rect 17049 25857 17083 25891
rect 23121 25857 23155 25891
rect 23305 25857 23339 25891
rect 26985 25857 27019 25891
rect 29653 25857 29687 25891
rect 35449 25857 35483 25891
rect 36369 25857 36403 25891
rect 36553 25857 36587 25891
rect 37841 25857 37875 25891
rect 2697 25789 2731 25823
rect 16773 25789 16807 25823
rect 22937 25789 22971 25823
rect 29469 25789 29503 25823
rect 38025 25721 38059 25755
rect 4077 25653 4111 25687
rect 4629 25653 4663 25687
rect 17417 25653 17451 25687
rect 29009 25653 29043 25687
rect 29837 25653 29871 25687
rect 35265 25653 35299 25687
rect 2881 25449 2915 25483
rect 6745 25449 6779 25483
rect 36369 25449 36403 25483
rect 2329 25381 2363 25415
rect 37197 25381 37231 25415
rect 38025 25381 38059 25415
rect 4261 25313 4295 25347
rect 4445 25313 4479 25347
rect 7297 25313 7331 25347
rect 36737 25313 36771 25347
rect 1685 25245 1719 25279
rect 2145 25245 2179 25279
rect 3065 25245 3099 25279
rect 7113 25245 7147 25279
rect 17049 25245 17083 25279
rect 23213 25245 23247 25279
rect 23397 25245 23431 25279
rect 26341 25245 26375 25279
rect 28733 25245 28767 25279
rect 31493 25245 31527 25279
rect 36553 25245 36587 25279
rect 37381 25245 37415 25279
rect 37841 25245 37875 25279
rect 7205 25177 7239 25211
rect 8033 25177 8067 25211
rect 22661 25177 22695 25211
rect 1501 25109 1535 25143
rect 3801 25109 3835 25143
rect 4169 25109 4203 25143
rect 5089 25109 5123 25143
rect 17233 25109 17267 25143
rect 23581 25109 23615 25143
rect 26525 25109 26559 25143
rect 28181 25109 28215 25143
rect 28917 25109 28951 25143
rect 31677 25109 31711 25143
rect 2513 24905 2547 24939
rect 19349 24905 19383 24939
rect 37381 24905 37415 24939
rect 1869 24769 1903 24803
rect 3065 24769 3099 24803
rect 7941 24769 7975 24803
rect 8401 24769 8435 24803
rect 14933 24769 14967 24803
rect 18225 24769 18259 24803
rect 23397 24769 23431 24803
rect 23581 24769 23615 24803
rect 37841 24769 37875 24803
rect 17969 24701 18003 24735
rect 23213 24701 23247 24735
rect 14749 24633 14783 24667
rect 1961 24565 1995 24599
rect 7757 24565 7791 24599
rect 17417 24565 17451 24599
rect 22661 24565 22695 24599
rect 38025 24565 38059 24599
rect 29009 24361 29043 24395
rect 31769 24361 31803 24395
rect 1593 24293 1627 24327
rect 37197 24293 37231 24327
rect 29561 24225 29595 24259
rect 36737 24225 36771 24259
rect 1409 24157 1443 24191
rect 2053 24157 2087 24191
rect 2697 24157 2731 24191
rect 14381 24157 14415 24191
rect 26249 24157 26283 24191
rect 29745 24157 29779 24191
rect 29929 24157 29963 24191
rect 31585 24157 31619 24191
rect 34989 24157 35023 24191
rect 35541 24157 35575 24191
rect 36553 24157 36587 24191
rect 37381 24157 37415 24191
rect 37841 24157 37875 24191
rect 36369 24089 36403 24123
rect 14197 24021 14231 24055
rect 26433 24021 26467 24055
rect 34805 24021 34839 24055
rect 35725 24021 35759 24055
rect 38025 24021 38059 24055
rect 8309 23817 8343 23851
rect 37381 23749 37415 23783
rect 1869 23681 1903 23715
rect 2513 23681 2547 23715
rect 9597 23681 9631 23715
rect 10057 23681 10091 23715
rect 37841 23681 37875 23715
rect 2053 23545 2087 23579
rect 29653 23545 29687 23579
rect 3157 23477 3191 23511
rect 35357 23477 35391 23511
rect 38025 23477 38059 23511
rect 1501 23273 1535 23307
rect 34805 23273 34839 23307
rect 8217 23205 8251 23239
rect 37197 23205 37231 23239
rect 7573 23137 7607 23171
rect 9689 23137 9723 23171
rect 29837 23137 29871 23171
rect 36553 23137 36587 23171
rect 1685 23069 1719 23103
rect 2145 23069 2179 23103
rect 2789 23069 2823 23103
rect 8953 23069 8987 23103
rect 23213 23069 23247 23103
rect 23397 23069 23431 23103
rect 30021 23069 30055 23103
rect 30205 23069 30239 23103
rect 31769 23069 31803 23103
rect 34989 23069 35023 23103
rect 36185 23069 36219 23103
rect 36369 23069 36403 23103
rect 37381 23069 37415 23103
rect 37841 23069 37875 23103
rect 7757 23001 7791 23035
rect 7849 23001 7883 23035
rect 9934 23001 9968 23035
rect 21281 23001 21315 23035
rect 21465 23001 21499 23035
rect 2329 22933 2363 22967
rect 9137 22933 9171 22967
rect 11069 22933 11103 22967
rect 22017 22933 22051 22967
rect 23581 22933 23615 22967
rect 31953 22933 31987 22967
rect 38025 22933 38059 22967
rect 9505 22729 9539 22763
rect 23305 22729 23339 22763
rect 1685 22593 1719 22627
rect 23121 22593 23155 22627
rect 24961 22593 24995 22627
rect 30297 22593 30331 22627
rect 34529 22593 34563 22627
rect 37841 22593 37875 22627
rect 23857 22525 23891 22559
rect 30113 22525 30147 22559
rect 37381 22525 37415 22559
rect 3341 22457 3375 22491
rect 34345 22457 34379 22491
rect 1501 22389 1535 22423
rect 2145 22389 2179 22423
rect 2789 22389 2823 22423
rect 25145 22389 25179 22423
rect 29561 22389 29595 22423
rect 30481 22389 30515 22423
rect 38025 22389 38059 22423
rect 21097 22185 21131 22219
rect 35725 22185 35759 22219
rect 1869 21981 1903 22015
rect 2513 21981 2547 22015
rect 3157 21981 3191 22015
rect 16405 21981 16439 22015
rect 20361 21981 20395 22015
rect 32229 21981 32263 22015
rect 35909 21981 35943 22015
rect 36093 21981 36127 22015
rect 37381 21981 37415 22015
rect 37841 21981 37875 22015
rect 2053 21913 2087 21947
rect 16138 21913 16172 21947
rect 36737 21913 36771 21947
rect 2697 21845 2731 21879
rect 15025 21845 15059 21879
rect 16957 21845 16991 21879
rect 20545 21845 20579 21879
rect 32413 21845 32447 21879
rect 37197 21845 37231 21879
rect 38025 21845 38059 21879
rect 4629 21641 4663 21675
rect 15025 21641 15059 21675
rect 25237 21641 25271 21675
rect 26249 21641 26283 21675
rect 1685 21505 1719 21539
rect 2697 21505 2731 21539
rect 2964 21505 2998 21539
rect 14841 21505 14875 21539
rect 20545 21505 20579 21539
rect 25421 21505 25455 21539
rect 26433 21505 26467 21539
rect 26985 21505 27019 21539
rect 28457 21505 28491 21539
rect 37841 21505 37875 21539
rect 20361 21437 20395 21471
rect 20729 21437 20763 21471
rect 21833 21437 21867 21471
rect 22109 21437 22143 21471
rect 1501 21301 1535 21335
rect 2145 21301 2179 21335
rect 4077 21301 4111 21335
rect 27169 21301 27203 21335
rect 28733 21301 28767 21335
rect 38025 21301 38059 21335
rect 2973 21097 3007 21131
rect 26525 21097 26559 21131
rect 3801 21029 3835 21063
rect 15209 21029 15243 21063
rect 26341 21029 26375 21063
rect 35541 21029 35575 21063
rect 4261 20961 4295 20995
rect 4445 20961 4479 20995
rect 14565 20961 14599 20995
rect 3157 20893 3191 20927
rect 4169 20893 4203 20927
rect 7021 20893 7055 20927
rect 14841 20893 14875 20927
rect 15669 20893 15703 20927
rect 20545 20893 20579 20927
rect 20729 20893 20763 20927
rect 35725 20893 35759 20927
rect 37381 20893 37415 20927
rect 37841 20893 37875 20927
rect 1869 20825 1903 20859
rect 2053 20825 2087 20859
rect 26065 20825 26099 20859
rect 36737 20825 36771 20859
rect 7205 20757 7239 20791
rect 14749 20757 14783 20791
rect 17141 20757 17175 20791
rect 20913 20757 20947 20791
rect 25605 20757 25639 20791
rect 37197 20757 37231 20791
rect 38025 20757 38059 20791
rect 6837 20553 6871 20587
rect 15577 20553 15611 20587
rect 26433 20553 26467 20587
rect 32597 20553 32631 20587
rect 1685 20417 1719 20451
rect 2145 20417 2179 20451
rect 2789 20417 2823 20451
rect 7205 20417 7239 20451
rect 20729 20417 20763 20451
rect 30389 20417 30423 20451
rect 30573 20417 30607 20451
rect 32413 20417 32447 20451
rect 37841 20417 37875 20451
rect 7297 20349 7331 20383
rect 7389 20349 7423 20383
rect 20545 20349 20579 20383
rect 25973 20349 26007 20383
rect 29653 20349 29687 20383
rect 30205 20349 30239 20383
rect 2329 20281 2363 20315
rect 26249 20281 26283 20315
rect 1501 20213 1535 20247
rect 3433 20213 3467 20247
rect 20913 20213 20947 20247
rect 25513 20213 25547 20247
rect 38025 20213 38059 20247
rect 8953 20009 8987 20043
rect 10517 20009 10551 20043
rect 35173 20009 35207 20043
rect 36921 20009 36955 20043
rect 6929 19873 6963 19907
rect 11069 19873 11103 19907
rect 22293 19873 22327 19907
rect 37289 19873 37323 19907
rect 7196 19805 7230 19839
rect 22569 19805 22603 19839
rect 37105 19805 37139 19839
rect 37841 19805 37875 19839
rect 1869 19737 1903 19771
rect 2513 19737 2547 19771
rect 11336 19737 11370 19771
rect 35265 19737 35299 19771
rect 1961 19669 1995 19703
rect 8309 19669 8343 19703
rect 12449 19669 12483 19703
rect 38025 19669 38059 19703
rect 11529 19465 11563 19499
rect 32597 19465 32631 19499
rect 35725 19465 35759 19499
rect 37289 19465 37323 19499
rect 1961 19329 1995 19363
rect 11713 19329 11747 19363
rect 22477 19329 22511 19363
rect 30297 19329 30331 19363
rect 30481 19329 30515 19363
rect 32413 19329 32447 19363
rect 35541 19329 35575 19363
rect 37473 19329 37507 19363
rect 2237 19261 2271 19295
rect 2697 19261 2731 19295
rect 22201 19261 22235 19295
rect 30113 19261 30147 19295
rect 37657 19261 37691 19295
rect 29561 19193 29595 19227
rect 36185 19125 36219 19159
rect 11437 18921 11471 18955
rect 26433 18921 26467 18955
rect 37381 18921 37415 18955
rect 12081 18785 12115 18819
rect 16589 18717 16623 18751
rect 26341 18717 26375 18751
rect 36737 18717 36771 18751
rect 37197 18717 37231 18751
rect 37841 18717 37875 18751
rect 1869 18649 1903 18683
rect 2513 18649 2547 18683
rect 11805 18649 11839 18683
rect 16856 18649 16890 18683
rect 26157 18649 26191 18683
rect 1961 18581 1995 18615
rect 11897 18581 11931 18615
rect 17969 18581 18003 18615
rect 18521 18581 18555 18615
rect 25605 18581 25639 18615
rect 38025 18581 38059 18615
rect 1501 18377 1535 18411
rect 32321 18377 32355 18411
rect 3433 18309 3467 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2789 18241 2823 18275
rect 16681 18241 16715 18275
rect 22017 18241 22051 18275
rect 28457 18241 28491 18275
rect 28917 18241 28951 18275
rect 29837 18241 29871 18275
rect 30021 18241 30055 18275
rect 30205 18241 30239 18275
rect 32137 18241 32171 18275
rect 34253 18241 34287 18275
rect 35725 18241 35759 18275
rect 35909 18241 35943 18275
rect 37841 18241 37875 18275
rect 21833 18173 21867 18207
rect 34069 18173 34103 18207
rect 36093 18173 36127 18207
rect 2329 18105 2363 18139
rect 16865 18105 16899 18139
rect 29101 18105 29135 18139
rect 22201 18037 22235 18071
rect 38025 18037 38059 18071
rect 15761 17833 15795 17867
rect 16681 17833 16715 17867
rect 25789 17833 25823 17867
rect 29745 17833 29779 17867
rect 37933 17833 37967 17867
rect 17233 17697 17267 17731
rect 20913 17697 20947 17731
rect 22661 17697 22695 17731
rect 22937 17697 22971 17731
rect 1685 17629 1719 17663
rect 17049 17629 17083 17663
rect 21097 17629 21131 17663
rect 24409 17629 24443 17663
rect 37473 17629 37507 17663
rect 38117 17629 38151 17663
rect 14473 17561 14507 17595
rect 24654 17561 24688 17595
rect 1501 17493 1535 17527
rect 2237 17493 2271 17527
rect 2789 17493 2823 17527
rect 3893 17493 3927 17527
rect 17141 17493 17175 17527
rect 21281 17493 21315 17527
rect 8033 17289 8067 17323
rect 24317 17289 24351 17323
rect 4813 17221 4847 17255
rect 34345 17221 34379 17255
rect 1961 17153 1995 17187
rect 2789 17153 2823 17187
rect 3056 17153 3090 17187
rect 12817 17153 12851 17187
rect 13553 17153 13587 17187
rect 29469 17153 29503 17187
rect 34529 17153 34563 17187
rect 37841 17153 37875 17187
rect 2237 17085 2271 17119
rect 29285 17085 29319 17119
rect 4169 16949 4203 16983
rect 13001 16949 13035 16983
rect 14381 16949 14415 16983
rect 28733 16949 28767 16983
rect 29653 16949 29687 16983
rect 37381 16949 37415 16983
rect 38025 16949 38059 16983
rect 1961 16745 1995 16779
rect 36093 16745 36127 16779
rect 37197 16677 37231 16711
rect 4261 16609 4295 16643
rect 4445 16609 4479 16643
rect 22569 16609 22603 16643
rect 22845 16609 22879 16643
rect 36461 16609 36495 16643
rect 2789 16541 2823 16575
rect 7941 16541 7975 16575
rect 30757 16541 30791 16575
rect 36277 16541 36311 16575
rect 37381 16541 37415 16575
rect 37841 16541 37875 16575
rect 1869 16473 1903 16507
rect 2605 16405 2639 16439
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 5089 16405 5123 16439
rect 7757 16405 7791 16439
rect 30941 16405 30975 16439
rect 38025 16405 38059 16439
rect 2973 16201 3007 16235
rect 8217 16133 8251 16167
rect 8769 16133 8803 16167
rect 1869 16065 1903 16099
rect 3157 16065 3191 16099
rect 29193 16065 29227 16099
rect 29377 16065 29411 16099
rect 30389 16065 30423 16099
rect 36369 16065 36403 16099
rect 37289 16065 37323 16099
rect 37473 16065 37507 16099
rect 3617 15997 3651 16031
rect 29009 15997 29043 16031
rect 37657 15997 37691 16031
rect 2053 15929 2087 15963
rect 28457 15929 28491 15963
rect 4261 15861 4295 15895
rect 7941 15861 7975 15895
rect 30573 15861 30607 15895
rect 36185 15861 36219 15895
rect 38025 15657 38059 15691
rect 6929 15521 6963 15555
rect 16221 15521 16255 15555
rect 1961 15453 1995 15487
rect 2237 15453 2271 15487
rect 2973 15453 3007 15487
rect 8953 15453 8987 15487
rect 11713 15453 11747 15487
rect 37105 15453 37139 15487
rect 37841 15453 37875 15487
rect 7196 15385 7230 15419
rect 16405 15385 16439 15419
rect 16497 15385 16531 15419
rect 2789 15317 2823 15351
rect 3893 15317 3927 15351
rect 8309 15317 8343 15351
rect 11897 15317 11931 15351
rect 16865 15317 16899 15351
rect 36277 15317 36311 15351
rect 37289 15317 37323 15351
rect 2513 15113 2547 15147
rect 7297 15113 7331 15147
rect 10885 15113 10919 15147
rect 17509 15113 17543 15147
rect 24961 15113 24995 15147
rect 36093 15113 36127 15147
rect 18674 15045 18708 15079
rect 1869 14977 1903 15011
rect 3065 14977 3099 15011
rect 7113 14977 7147 15011
rect 11713 14977 11747 15011
rect 11980 14977 12014 15011
rect 17325 14977 17359 15011
rect 23489 14977 23523 15011
rect 23673 14977 23707 15011
rect 24317 14977 24351 15011
rect 33333 14977 33367 15011
rect 35909 14977 35943 15011
rect 36553 14977 36587 15011
rect 37841 14977 37875 15011
rect 18429 14909 18463 14943
rect 33149 14909 33183 14943
rect 33517 14909 33551 14943
rect 19809 14841 19843 14875
rect 36737 14841 36771 14875
rect 1961 14773 1995 14807
rect 13093 14773 13127 14807
rect 24501 14773 24535 14807
rect 38025 14773 38059 14807
rect 24409 14569 24443 14603
rect 26525 14569 26559 14603
rect 37197 14569 37231 14603
rect 32597 14501 32631 14535
rect 12357 14433 12391 14467
rect 13001 14433 13035 14467
rect 33149 14433 33183 14467
rect 1409 14365 1443 14399
rect 2053 14365 2087 14399
rect 12081 14365 12115 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 27077 14365 27111 14399
rect 28181 14365 28215 14399
rect 28365 14365 28399 14399
rect 28549 14365 28583 14399
rect 29653 14365 29687 14399
rect 33333 14365 33367 14399
rect 36737 14365 36771 14399
rect 37381 14365 37415 14399
rect 37841 14365 37875 14399
rect 12173 14297 12207 14331
rect 1593 14229 1627 14263
rect 2697 14229 2731 14263
rect 11713 14229 11747 14263
rect 18337 14229 18371 14263
rect 27261 14229 27295 14263
rect 29837 14229 29871 14263
rect 33517 14229 33551 14263
rect 38025 14229 38059 14263
rect 6929 14025 6963 14059
rect 24317 14025 24351 14059
rect 27997 14025 28031 14059
rect 32505 14025 32539 14059
rect 37933 14025 37967 14059
rect 23029 13957 23063 13991
rect 1869 13889 1903 13923
rect 3065 13889 3099 13923
rect 7297 13889 7331 13923
rect 22017 13889 22051 13923
rect 22293 13889 22327 13923
rect 22477 13889 22511 13923
rect 24409 13889 24443 13923
rect 33057 13889 33091 13923
rect 33241 13889 33275 13923
rect 33425 13889 33459 13923
rect 37289 13889 37323 13923
rect 38117 13889 38151 13923
rect 7389 13821 7423 13855
rect 7573 13821 7607 13855
rect 8217 13821 8251 13855
rect 21281 13821 21315 13855
rect 21833 13821 21867 13855
rect 23489 13821 23523 13855
rect 36737 13821 36771 13855
rect 2053 13753 2087 13787
rect 2513 13685 2547 13719
rect 37473 13685 37507 13719
rect 1501 13481 1535 13515
rect 2329 13481 2363 13515
rect 24869 13481 24903 13515
rect 25237 13345 25271 13379
rect 1685 13277 1719 13311
rect 2145 13277 2179 13311
rect 2789 13277 2823 13311
rect 25053 13277 25087 13311
rect 28273 13277 28307 13311
rect 28457 13277 28491 13311
rect 36093 13277 36127 13311
rect 36737 13277 36771 13311
rect 37841 13277 37875 13311
rect 27721 13209 27755 13243
rect 28641 13141 28675 13175
rect 36277 13141 36311 13175
rect 36921 13141 36955 13175
rect 38025 13141 38059 13175
rect 4813 12937 4847 12971
rect 15117 12937 15151 12971
rect 1869 12801 1903 12835
rect 2881 12801 2915 12835
rect 3148 12801 3182 12835
rect 14933 12801 14967 12835
rect 15117 12801 15151 12835
rect 15301 12801 15335 12835
rect 15945 12801 15979 12835
rect 33149 12801 33183 12835
rect 37841 12801 37875 12835
rect 14289 12733 14323 12767
rect 32965 12733 32999 12767
rect 2053 12665 2087 12699
rect 32413 12665 32447 12699
rect 38025 12665 38059 12699
rect 4261 12597 4295 12631
rect 33333 12597 33367 12631
rect 1501 12393 1535 12427
rect 3065 12393 3099 12427
rect 29837 12393 29871 12427
rect 2329 12325 2363 12359
rect 32321 12325 32355 12359
rect 4261 12257 4295 12291
rect 4353 12257 4387 12291
rect 5089 12257 5123 12291
rect 32781 12257 32815 12291
rect 1685 12189 1719 12223
rect 2145 12189 2179 12223
rect 3249 12189 3283 12223
rect 4169 12189 4203 12223
rect 28365 12189 28399 12223
rect 28549 12189 28583 12223
rect 30389 12189 30423 12223
rect 30665 12189 30699 12223
rect 32137 12189 32171 12223
rect 32965 12189 32999 12223
rect 36645 12189 36679 12223
rect 37841 12189 37875 12223
rect 23213 12121 23247 12155
rect 27813 12121 27847 12155
rect 3801 12053 3835 12087
rect 14565 12053 14599 12087
rect 23121 12053 23155 12087
rect 28733 12053 28767 12087
rect 33149 12053 33183 12087
rect 36829 12053 36863 12087
rect 38025 12053 38059 12087
rect 2145 11849 2179 11883
rect 24225 11849 24259 11883
rect 32597 11849 32631 11883
rect 2789 11781 2823 11815
rect 1685 11713 1719 11747
rect 15853 11713 15887 11747
rect 24409 11713 24443 11747
rect 36553 11713 36587 11747
rect 37841 11713 37875 11747
rect 24593 11645 24627 11679
rect 3341 11577 3375 11611
rect 36737 11577 36771 11611
rect 1501 11509 1535 11543
rect 8769 11509 8803 11543
rect 16037 11509 16071 11543
rect 38025 11509 38059 11543
rect 2697 11305 2731 11339
rect 37197 11305 37231 11339
rect 8217 11237 8251 11271
rect 23397 11237 23431 11271
rect 34897 11237 34931 11271
rect 38025 11237 38059 11271
rect 22109 11169 22143 11203
rect 28641 11169 28675 11203
rect 2513 11101 2547 11135
rect 3157 11101 3191 11135
rect 8033 11101 8067 11135
rect 8953 11101 8987 11135
rect 9209 11101 9243 11135
rect 18061 11101 18095 11135
rect 21281 11101 21315 11135
rect 21465 11101 21499 11135
rect 21649 11101 21683 11135
rect 28273 11101 28307 11135
rect 28457 11101 28491 11135
rect 34713 11101 34747 11135
rect 36737 11101 36771 11135
rect 37381 11101 37415 11135
rect 37841 11101 37875 11135
rect 1869 11033 1903 11067
rect 2053 11033 2087 11067
rect 23581 11033 23615 11067
rect 27721 11033 27755 11067
rect 10333 10965 10367 10999
rect 18245 10965 18279 10999
rect 2145 10761 2179 10795
rect 10149 10761 10183 10795
rect 15301 10761 15335 10795
rect 19441 10761 19475 10795
rect 24409 10761 24443 10795
rect 9597 10693 9631 10727
rect 13001 10693 13035 10727
rect 1685 10625 1719 10659
rect 12357 10625 12391 10659
rect 14749 10625 14783 10659
rect 17601 10625 17635 10659
rect 18061 10625 18095 10659
rect 18328 10625 18362 10659
rect 24593 10625 24627 10659
rect 36553 10625 36587 10659
rect 37841 10625 37875 10659
rect 2789 10557 2823 10591
rect 24777 10557 24811 10591
rect 1501 10421 1535 10455
rect 8309 10421 8343 10455
rect 12541 10421 12575 10455
rect 36737 10421 36771 10455
rect 38025 10421 38059 10455
rect 8125 10217 8159 10251
rect 12265 10217 12299 10251
rect 17877 10217 17911 10251
rect 36369 10217 36403 10251
rect 37197 10217 37231 10251
rect 23029 10149 23063 10183
rect 7481 10081 7515 10115
rect 9045 10081 9079 10115
rect 12725 10081 12759 10115
rect 12817 10081 12851 10115
rect 14381 10081 14415 10115
rect 14841 10081 14875 10115
rect 18429 10081 18463 10115
rect 28641 10081 28675 10115
rect 2053 10013 2087 10047
rect 27721 10013 27755 10047
rect 28273 10013 28307 10047
rect 28457 10013 28491 10047
rect 30113 10013 30147 10047
rect 35909 10013 35943 10047
rect 36553 10013 36587 10047
rect 37013 10013 37047 10047
rect 37841 10013 37875 10047
rect 1869 9945 1903 9979
rect 2513 9945 2547 9979
rect 7757 9945 7791 9979
rect 15086 9945 15120 9979
rect 17325 9945 17359 9979
rect 18245 9945 18279 9979
rect 23213 9945 23247 9979
rect 29929 9945 29963 9979
rect 3065 9877 3099 9911
rect 7665 9877 7699 9911
rect 11713 9877 11747 9911
rect 12633 9877 12667 9911
rect 13553 9877 13587 9911
rect 16221 9877 16255 9911
rect 18337 9877 18371 9911
rect 38025 9877 38059 9911
rect 1593 9673 1627 9707
rect 29837 9673 29871 9707
rect 36737 9673 36771 9707
rect 24133 9605 24167 9639
rect 31493 9605 31527 9639
rect 1409 9537 1443 9571
rect 2053 9537 2087 9571
rect 3249 9537 3283 9571
rect 24317 9537 24351 9571
rect 24501 9537 24535 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 34345 9537 34379 9571
rect 36553 9537 36587 9571
rect 37841 9537 37875 9571
rect 2697 9469 2731 9503
rect 27077 9469 27111 9503
rect 27537 9469 27571 9503
rect 27813 9469 27847 9503
rect 34161 9469 34195 9503
rect 2237 9401 2271 9435
rect 32505 9401 32539 9435
rect 38025 9401 38059 9435
rect 3433 9333 3467 9367
rect 33609 9333 33643 9367
rect 34529 9333 34563 9367
rect 3249 9129 3283 9163
rect 5181 9061 5215 9095
rect 2605 8993 2639 9027
rect 32781 8993 32815 9027
rect 37565 8993 37599 9027
rect 1685 8925 1719 8959
rect 3801 8925 3835 8959
rect 33057 8925 33091 8959
rect 36645 8925 36679 8959
rect 37289 8925 37323 8959
rect 2881 8857 2915 8891
rect 4046 8857 4080 8891
rect 1501 8789 1535 8823
rect 2789 8789 2823 8823
rect 5825 8789 5859 8823
rect 36829 8789 36863 8823
rect 2697 8585 2731 8619
rect 3985 8585 4019 8619
rect 33793 8585 33827 8619
rect 37381 8517 37415 8551
rect 1869 8449 1903 8483
rect 2881 8449 2915 8483
rect 27169 8449 27203 8483
rect 34345 8449 34379 8483
rect 34529 8449 34563 8483
rect 36553 8449 36587 8483
rect 37841 8449 37875 8483
rect 3433 8381 3467 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 2053 8313 2087 8347
rect 27353 8313 27387 8347
rect 36737 8313 36771 8347
rect 38025 8313 38059 8347
rect 34713 8245 34747 8279
rect 1593 8041 1627 8075
rect 20085 7905 20119 7939
rect 1409 7837 1443 7871
rect 2053 7837 2087 7871
rect 19257 7837 19291 7871
rect 29653 7837 29687 7871
rect 29837 7837 29871 7871
rect 30021 7837 30055 7871
rect 37013 7837 37047 7871
rect 37841 7837 37875 7871
rect 2697 7769 2731 7803
rect 20330 7769 20364 7803
rect 2237 7701 2271 7735
rect 8125 7701 8159 7735
rect 19441 7701 19475 7735
rect 21465 7701 21499 7735
rect 37197 7701 37231 7735
rect 38025 7701 38059 7735
rect 2145 7497 2179 7531
rect 7297 7497 7331 7531
rect 7389 7497 7423 7531
rect 18613 7497 18647 7531
rect 19993 7497 20027 7531
rect 2789 7429 2823 7463
rect 18245 7429 18279 7463
rect 1685 7361 1719 7395
rect 8217 7361 8251 7395
rect 8484 7361 8518 7395
rect 18153 7361 18187 7395
rect 31401 7361 31435 7395
rect 32137 7361 32171 7395
rect 32321 7361 32355 7395
rect 36553 7361 36587 7395
rect 37841 7361 37875 7395
rect 7205 7293 7239 7327
rect 10057 7293 10091 7327
rect 17969 7293 18003 7327
rect 31217 7293 31251 7327
rect 31585 7225 31619 7259
rect 1501 7157 1535 7191
rect 7757 7157 7791 7191
rect 9597 7157 9631 7191
rect 30665 7157 30699 7191
rect 32505 7157 32539 7191
rect 36737 7157 36771 7191
rect 38025 7157 38059 7191
rect 7665 6953 7699 6987
rect 8309 6953 8343 6987
rect 37197 6953 37231 6987
rect 16037 6817 16071 6851
rect 8125 6749 8159 6783
rect 13001 6749 13035 6783
rect 14105 6749 14139 6783
rect 27721 6749 27755 6783
rect 27905 6749 27939 6783
rect 28089 6749 28123 6783
rect 36737 6749 36771 6783
rect 37381 6749 37415 6783
rect 37841 6749 37875 6783
rect 1869 6681 1903 6715
rect 2053 6681 2087 6715
rect 14350 6681 14384 6715
rect 2513 6613 2547 6647
rect 13185 6613 13219 6647
rect 15485 6613 15519 6647
rect 27169 6613 27203 6647
rect 38025 6613 38059 6647
rect 2697 6409 2731 6443
rect 11989 6409 12023 6443
rect 13277 6409 13311 6443
rect 13829 6409 13863 6443
rect 36737 6409 36771 6443
rect 1961 6273 1995 6307
rect 2881 6273 2915 6307
rect 12909 6273 12943 6307
rect 24584 6273 24618 6307
rect 33333 6273 33367 6307
rect 36553 6273 36587 6307
rect 37841 6273 37875 6307
rect 2237 6205 2271 6239
rect 3893 6205 3927 6239
rect 12633 6205 12667 6239
rect 12817 6205 12851 6239
rect 23857 6205 23891 6239
rect 24317 6205 24351 6239
rect 3433 6069 3467 6103
rect 25697 6069 25731 6103
rect 33517 6069 33551 6103
rect 38025 6069 38059 6103
rect 29653 5865 29687 5899
rect 34069 5865 34103 5899
rect 37197 5797 37231 5831
rect 30021 5729 30055 5763
rect 1685 5661 1719 5695
rect 2145 5661 2179 5695
rect 2789 5661 2823 5695
rect 29837 5661 29871 5695
rect 34713 5661 34747 5695
rect 34897 5661 34931 5695
rect 36737 5661 36771 5695
rect 37381 5661 37415 5695
rect 37841 5661 37875 5695
rect 1501 5525 1535 5559
rect 2329 5525 2363 5559
rect 35081 5525 35115 5559
rect 38025 5525 38059 5559
rect 36737 5321 36771 5355
rect 1869 5185 1903 5219
rect 2513 5185 2547 5219
rect 3157 5185 3191 5219
rect 36553 5185 36587 5219
rect 37841 5185 37875 5219
rect 3709 5117 3743 5151
rect 2053 5049 2087 5083
rect 2697 4981 2731 5015
rect 38025 4981 38059 5015
rect 2697 4777 2731 4811
rect 24409 4777 24443 4811
rect 27261 4777 27295 4811
rect 2053 4641 2087 4675
rect 6009 4641 6043 4675
rect 27813 4641 27847 4675
rect 2881 4573 2915 4607
rect 24593 4573 24627 4607
rect 24961 4573 24995 4607
rect 27997 4573 28031 4607
rect 32873 4573 32907 4607
rect 37197 4573 37231 4607
rect 37841 4573 37875 4607
rect 1869 4505 1903 4539
rect 4353 4505 4387 4539
rect 5825 4505 5859 4539
rect 24685 4505 24719 4539
rect 24777 4505 24811 4539
rect 3893 4437 3927 4471
rect 5365 4437 5399 4471
rect 5733 4437 5767 4471
rect 6653 4437 6687 4471
rect 23765 4437 23799 4471
rect 28181 4437 28215 4471
rect 33057 4437 33091 4471
rect 36185 4437 36219 4471
rect 37013 4437 37047 4471
rect 38025 4437 38059 4471
rect 5733 4233 5767 4267
rect 6469 4233 6503 4267
rect 24225 4165 24259 4199
rect 1685 4097 1719 4131
rect 2881 4097 2915 4131
rect 3433 4097 3467 4131
rect 4620 4097 4654 4131
rect 16865 4097 16899 4131
rect 17049 4097 17083 4131
rect 17141 4097 17175 4131
rect 18981 4097 19015 4131
rect 20554 4097 20588 4131
rect 20821 4097 20855 4131
rect 23029 4097 23063 4131
rect 23213 4097 23247 4131
rect 24041 4097 24075 4131
rect 24317 4097 24351 4131
rect 24409 4097 24443 4131
rect 28181 4097 28215 4131
rect 28825 4097 28859 4131
rect 30113 4097 30147 4131
rect 33609 4097 33643 4131
rect 36093 4097 36127 4131
rect 36553 4097 36587 4131
rect 37841 4097 37875 4131
rect 4353 4029 4387 4063
rect 23121 4029 23155 4063
rect 28273 4029 28307 4063
rect 30297 4029 30331 4063
rect 33425 4029 33459 4063
rect 2697 3961 2731 3995
rect 19441 3961 19475 3995
rect 24593 3961 24627 3995
rect 29929 3961 29963 3995
rect 35909 3961 35943 3995
rect 36737 3961 36771 3995
rect 1501 3893 1535 3927
rect 2145 3893 2179 3927
rect 16681 3893 16715 3927
rect 22477 3893 22511 3927
rect 32873 3893 32907 3927
rect 33793 3893 33827 3927
rect 38025 3893 38059 3927
rect 4905 3689 4939 3723
rect 15117 3689 15151 3723
rect 19625 3689 19659 3723
rect 20637 3689 20671 3723
rect 24501 3689 24535 3723
rect 35081 3689 35115 3723
rect 6009 3621 6043 3655
rect 15577 3621 15611 3655
rect 20269 3621 20303 3655
rect 35725 3621 35759 3655
rect 2605 3553 2639 3587
rect 9137 3553 9171 3587
rect 16957 3553 16991 3587
rect 29929 3553 29963 3587
rect 2697 3485 2731 3519
rect 2973 3485 3007 3519
rect 5089 3485 5123 3519
rect 10241 3485 10275 3519
rect 11069 3485 11103 3519
rect 16690 3485 16724 3519
rect 20177 3485 20211 3519
rect 20453 3485 20487 3519
rect 24593 3485 24627 3519
rect 25053 3485 25087 3519
rect 27721 3485 27755 3519
rect 27905 3485 27939 3519
rect 30113 3485 30147 3519
rect 30297 3485 30331 3519
rect 33333 3485 33367 3519
rect 33517 3485 33551 3519
rect 33701 3485 33735 3519
rect 34897 3485 34931 3519
rect 35541 3485 35575 3519
rect 36461 3485 36495 3519
rect 37105 3485 37139 3519
rect 37841 3485 37875 3519
rect 1869 3417 1903 3451
rect 9321 3417 9355 3451
rect 11314 3417 11348 3451
rect 32781 3417 32815 3451
rect 1961 3349 1995 3383
rect 3801 3349 3835 3383
rect 9413 3349 9447 3383
rect 9781 3349 9815 3383
rect 10425 3349 10459 3383
rect 12449 3349 12483 3383
rect 27169 3349 27203 3383
rect 28089 3349 28123 3383
rect 36645 3349 36679 3383
rect 37289 3349 37323 3383
rect 38025 3349 38059 3383
rect 9965 3145 9999 3179
rect 10977 3145 11011 3179
rect 1869 3077 1903 3111
rect 36645 3077 36679 3111
rect 2789 3009 2823 3043
rect 3249 3009 3283 3043
rect 3893 3009 3927 3043
rect 8861 3009 8895 3043
rect 35449 3009 35483 3043
rect 35909 3009 35943 3043
rect 36553 3009 36587 3043
rect 37841 3009 37875 3043
rect 2053 2873 2087 2907
rect 36093 2873 36127 2907
rect 2605 2805 2639 2839
rect 3433 2805 3467 2839
rect 4445 2805 4479 2839
rect 4997 2805 5031 2839
rect 34805 2805 34839 2839
rect 38025 2805 38059 2839
rect 3801 2601 3835 2635
rect 4445 2601 4479 2635
rect 35081 2601 35115 2635
rect 2145 2533 2179 2567
rect 36645 2533 36679 2567
rect 5089 2465 5123 2499
rect 1869 2397 1903 2431
rect 2973 2397 3007 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 35265 2397 35299 2431
rect 36001 2397 36035 2431
rect 36461 2397 36495 2431
rect 37841 2397 37875 2431
rect 5641 2329 5675 2363
rect 2789 2261 2823 2295
rect 35817 2261 35851 2295
rect 38025 2261 38059 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 2590 37408 2596 37460
rect 2648 37448 2654 37460
rect 6365 37451 6423 37457
rect 6365 37448 6377 37451
rect 2648 37420 6377 37448
rect 2648 37408 2654 37420
rect 6365 37417 6377 37420
rect 6411 37417 6423 37451
rect 6365 37411 6423 37417
rect 3878 37340 3884 37392
rect 3936 37380 3942 37392
rect 6917 37383 6975 37389
rect 6917 37380 6929 37383
rect 3936 37352 6929 37380
rect 3936 37340 3942 37352
rect 6917 37349 6929 37352
rect 6963 37349 6975 37383
rect 6917 37343 6975 37349
rect 2038 37312 2044 37324
rect 1999 37284 2044 37312
rect 2038 37272 2044 37284
rect 2096 37272 2102 37324
rect 2777 37315 2835 37321
rect 2777 37281 2789 37315
rect 2823 37312 2835 37315
rect 3694 37312 3700 37324
rect 2823 37284 3700 37312
rect 2823 37281 2835 37284
rect 2777 37275 2835 37281
rect 3694 37272 3700 37284
rect 3752 37272 3758 37324
rect 5261 37315 5319 37321
rect 5261 37312 5273 37315
rect 3804 37284 5273 37312
rect 1854 37244 1860 37256
rect 1767 37216 1860 37244
rect 1854 37204 1860 37216
rect 1912 37244 1918 37256
rect 3804 37244 3832 37284
rect 5261 37281 5273 37284
rect 5307 37281 5319 37315
rect 5261 37275 5319 37281
rect 35544 37284 35848 37312
rect 1912 37216 3832 37244
rect 1912 37204 1918 37216
rect 3878 37204 3884 37256
rect 3936 37244 3942 37256
rect 4525 37247 4583 37253
rect 3936 37216 3981 37244
rect 3936 37204 3942 37216
rect 4525 37213 4537 37247
rect 4571 37244 4583 37247
rect 4614 37244 4620 37256
rect 4571 37216 4620 37244
rect 4571 37213 4583 37216
rect 4525 37207 4583 37213
rect 4614 37204 4620 37216
rect 4672 37204 4678 37256
rect 33870 37244 33876 37256
rect 33831 37216 33876 37244
rect 33870 37204 33876 37216
rect 33928 37204 33934 37256
rect 34977 37247 35035 37253
rect 34977 37213 34989 37247
rect 35023 37213 35035 37247
rect 34977 37207 35035 37213
rect 2590 37176 2596 37188
rect 2551 37148 2596 37176
rect 2590 37136 2596 37148
rect 2648 37136 2654 37188
rect 4062 37176 4068 37188
rect 4023 37148 4068 37176
rect 4062 37136 4068 37148
rect 4120 37136 4126 37188
rect 26786 37136 26792 37188
rect 26844 37176 26850 37188
rect 34992 37176 35020 37207
rect 35066 37204 35072 37256
rect 35124 37244 35130 37256
rect 35544 37244 35572 37284
rect 35710 37244 35716 37256
rect 35124 37216 35572 37244
rect 35671 37216 35716 37244
rect 35124 37204 35130 37216
rect 35710 37204 35716 37216
rect 35768 37204 35774 37256
rect 35820 37244 35848 37284
rect 36372 37284 36584 37312
rect 36372 37244 36400 37284
rect 35820 37216 36400 37244
rect 36449 37247 36507 37253
rect 36449 37213 36461 37247
rect 36495 37213 36507 37247
rect 36556 37244 36584 37284
rect 37182 37272 37188 37324
rect 37240 37312 37246 37324
rect 37277 37315 37335 37321
rect 37277 37312 37289 37315
rect 37240 37284 37289 37312
rect 37240 37272 37246 37284
rect 37277 37281 37289 37284
rect 37323 37281 37335 37315
rect 37277 37275 37335 37281
rect 37553 37247 37611 37253
rect 37553 37244 37565 37247
rect 36556 37216 37565 37244
rect 36449 37207 36507 37213
rect 37553 37213 37565 37216
rect 37599 37213 37611 37247
rect 37553 37207 37611 37213
rect 26844 37148 35020 37176
rect 26844 37136 26850 37148
rect 35434 37136 35440 37188
rect 35492 37176 35498 37188
rect 35492 37148 36216 37176
rect 35492 37136 35498 37148
rect 1762 37068 1768 37120
rect 1820 37108 1826 37120
rect 3878 37108 3884 37120
rect 1820 37080 3884 37108
rect 1820 37068 1826 37080
rect 3878 37068 3884 37080
rect 3936 37068 3942 37120
rect 3970 37068 3976 37120
rect 4028 37108 4034 37120
rect 4709 37111 4767 37117
rect 4709 37108 4721 37111
rect 4028 37080 4721 37108
rect 4028 37068 4034 37080
rect 4709 37077 4721 37080
rect 4755 37077 4767 37111
rect 4709 37071 4767 37077
rect 34057 37111 34115 37117
rect 34057 37077 34069 37111
rect 34103 37108 34115 37111
rect 34514 37108 34520 37120
rect 34103 37080 34520 37108
rect 34103 37077 34115 37080
rect 34057 37071 34115 37077
rect 34514 37068 34520 37080
rect 34572 37068 34578 37120
rect 35161 37111 35219 37117
rect 35161 37077 35173 37111
rect 35207 37108 35219 37111
rect 35342 37108 35348 37120
rect 35207 37080 35348 37108
rect 35207 37077 35219 37080
rect 35161 37071 35219 37077
rect 35342 37068 35348 37080
rect 35400 37068 35406 37120
rect 35802 37068 35808 37120
rect 35860 37108 35866 37120
rect 35897 37111 35955 37117
rect 35897 37108 35909 37111
rect 35860 37080 35909 37108
rect 35860 37068 35866 37080
rect 35897 37077 35909 37080
rect 35943 37077 35955 37111
rect 36188 37108 36216 37148
rect 36464 37108 36492 37207
rect 36630 37108 36636 37120
rect 36188 37080 36492 37108
rect 36591 37080 36636 37108
rect 35897 37071 35955 37077
rect 36630 37068 36636 37080
rect 36688 37068 36694 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 3326 36904 3332 36916
rect 3287 36876 3332 36904
rect 3326 36864 3332 36876
rect 3384 36864 3390 36916
rect 3878 36864 3884 36916
rect 3936 36904 3942 36916
rect 5261 36907 5319 36913
rect 5261 36904 5273 36907
rect 3936 36876 5273 36904
rect 3936 36864 3942 36876
rect 5261 36873 5273 36876
rect 5307 36873 5319 36907
rect 29730 36904 29736 36916
rect 29691 36876 29736 36904
rect 5261 36867 5319 36873
rect 29730 36864 29736 36876
rect 29788 36864 29794 36916
rect 35253 36907 35311 36913
rect 35253 36873 35265 36907
rect 35299 36904 35311 36907
rect 35526 36904 35532 36916
rect 35299 36876 35532 36904
rect 35299 36873 35311 36876
rect 35253 36867 35311 36873
rect 35526 36864 35532 36876
rect 35584 36864 35590 36916
rect 1762 36796 1768 36848
rect 1820 36836 1826 36848
rect 1857 36839 1915 36845
rect 1857 36836 1869 36839
rect 1820 36808 1869 36836
rect 1820 36796 1826 36808
rect 1857 36805 1869 36808
rect 1903 36805 1915 36839
rect 1857 36799 1915 36805
rect 2866 36796 2872 36848
rect 2924 36836 2930 36848
rect 4709 36839 4767 36845
rect 4709 36836 4721 36839
rect 2924 36808 4721 36836
rect 2924 36796 2930 36808
rect 4709 36805 4721 36808
rect 4755 36805 4767 36839
rect 4709 36799 4767 36805
rect 22462 36796 22468 36848
rect 22520 36836 22526 36848
rect 22520 36808 37596 36836
rect 22520 36796 22526 36808
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36768 2835 36771
rect 3326 36768 3332 36780
rect 2823 36740 3332 36768
rect 2823 36737 2835 36740
rect 2777 36731 2835 36737
rect 3326 36728 3332 36740
rect 3384 36728 3390 36780
rect 3510 36768 3516 36780
rect 3471 36740 3516 36768
rect 3510 36728 3516 36740
rect 3568 36728 3574 36780
rect 3970 36768 3976 36780
rect 3931 36740 3976 36768
rect 3970 36728 3976 36740
rect 4028 36728 4034 36780
rect 24581 36771 24639 36777
rect 24581 36737 24593 36771
rect 24627 36768 24639 36771
rect 33965 36771 34023 36777
rect 24627 36740 25360 36768
rect 24627 36737 24639 36740
rect 24581 36731 24639 36737
rect 2041 36703 2099 36709
rect 2041 36669 2053 36703
rect 2087 36700 2099 36703
rect 24302 36700 24308 36712
rect 2087 36672 24308 36700
rect 2087 36669 2099 36672
rect 2041 36663 2099 36669
rect 24302 36660 24308 36672
rect 24360 36660 24366 36712
rect 24397 36703 24455 36709
rect 24397 36669 24409 36703
rect 24443 36669 24455 36703
rect 24397 36663 24455 36669
rect 4062 36592 4068 36644
rect 4120 36632 4126 36644
rect 23845 36635 23903 36641
rect 23845 36632 23857 36635
rect 4120 36604 23857 36632
rect 4120 36592 4126 36604
rect 23845 36601 23857 36604
rect 23891 36632 23903 36635
rect 24412 36632 24440 36663
rect 23891 36604 24440 36632
rect 23891 36601 23903 36604
rect 23845 36595 23903 36601
rect 2593 36567 2651 36573
rect 2593 36533 2605 36567
rect 2639 36564 2651 36567
rect 2774 36564 2780 36576
rect 2639 36536 2780 36564
rect 2639 36533 2651 36536
rect 2593 36527 2651 36533
rect 2774 36524 2780 36536
rect 2832 36524 2838 36576
rect 3786 36524 3792 36576
rect 3844 36564 3850 36576
rect 4157 36567 4215 36573
rect 4157 36564 4169 36567
rect 3844 36536 4169 36564
rect 3844 36524 3850 36536
rect 4157 36533 4169 36536
rect 4203 36533 4215 36567
rect 24762 36564 24768 36576
rect 24723 36536 24768 36564
rect 4157 36527 4215 36533
rect 24762 36524 24768 36536
rect 24820 36524 24826 36576
rect 25332 36573 25360 36740
rect 33965 36737 33977 36771
rect 34011 36768 34023 36771
rect 34425 36771 34483 36777
rect 34425 36768 34437 36771
rect 34011 36740 34437 36768
rect 34011 36737 34023 36740
rect 33965 36731 34023 36737
rect 34425 36737 34437 36740
rect 34471 36768 34483 36771
rect 34698 36768 34704 36780
rect 34471 36740 34704 36768
rect 34471 36737 34483 36740
rect 34425 36731 34483 36737
rect 34698 36728 34704 36740
rect 34756 36728 34762 36780
rect 34790 36728 34796 36780
rect 34848 36768 34854 36780
rect 35069 36771 35127 36777
rect 35069 36768 35081 36771
rect 34848 36740 35081 36768
rect 34848 36728 34854 36740
rect 35069 36737 35081 36740
rect 35115 36737 35127 36771
rect 35986 36768 35992 36780
rect 35947 36740 35992 36768
rect 35069 36731 35127 36737
rect 35986 36728 35992 36740
rect 36044 36728 36050 36780
rect 37274 36768 37280 36780
rect 37235 36740 37280 36768
rect 37274 36728 37280 36740
rect 37332 36728 37338 36780
rect 37568 36777 37596 36808
rect 37553 36771 37611 36777
rect 37553 36737 37565 36771
rect 37599 36737 37611 36771
rect 37553 36731 37611 36737
rect 35805 36703 35863 36709
rect 35805 36669 35817 36703
rect 35851 36669 35863 36703
rect 35805 36663 35863 36669
rect 34609 36635 34667 36641
rect 34609 36601 34621 36635
rect 34655 36632 34667 36635
rect 35820 36632 35848 36663
rect 34655 36604 35848 36632
rect 34655 36601 34667 36604
rect 34609 36595 34667 36601
rect 25317 36567 25375 36573
rect 25317 36533 25329 36567
rect 25363 36564 25375 36567
rect 25498 36564 25504 36576
rect 25363 36536 25504 36564
rect 25363 36533 25375 36536
rect 25317 36527 25375 36533
rect 25498 36524 25504 36536
rect 25556 36524 25562 36576
rect 30653 36567 30711 36573
rect 30653 36533 30665 36567
rect 30699 36564 30711 36567
rect 30742 36564 30748 36576
rect 30699 36536 30748 36564
rect 30699 36533 30711 36536
rect 30653 36527 30711 36533
rect 30742 36524 30748 36536
rect 30800 36524 30806 36576
rect 35894 36524 35900 36576
rect 35952 36564 35958 36576
rect 36173 36567 36231 36573
rect 36173 36564 36185 36567
rect 35952 36536 36185 36564
rect 35952 36524 35958 36536
rect 36173 36533 36185 36536
rect 36219 36533 36231 36567
rect 36173 36527 36231 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 3326 36320 3332 36372
rect 3384 36360 3390 36372
rect 3789 36363 3847 36369
rect 3789 36360 3801 36363
rect 3384 36332 3801 36360
rect 3384 36320 3390 36332
rect 3789 36329 3801 36332
rect 3835 36329 3847 36363
rect 5166 36360 5172 36372
rect 5127 36332 5172 36360
rect 3789 36323 3847 36329
rect 5166 36320 5172 36332
rect 5224 36320 5230 36372
rect 30282 36360 30288 36372
rect 20824 36332 30288 36360
rect 2041 36295 2099 36301
rect 2041 36261 2053 36295
rect 2087 36292 2099 36295
rect 2130 36292 2136 36304
rect 2087 36264 2136 36292
rect 2087 36261 2099 36264
rect 2041 36255 2099 36261
rect 2130 36252 2136 36264
rect 2188 36252 2194 36304
rect 5184 36224 5212 36320
rect 20824 36233 20852 36332
rect 30282 36320 30288 36332
rect 30340 36320 30346 36372
rect 33781 36363 33839 36369
rect 33781 36329 33793 36363
rect 33827 36360 33839 36363
rect 35710 36360 35716 36372
rect 33827 36332 35716 36360
rect 33827 36329 33839 36332
rect 33781 36323 33839 36329
rect 35710 36320 35716 36332
rect 35768 36320 35774 36372
rect 36170 36360 36176 36372
rect 36131 36332 36176 36360
rect 36170 36320 36176 36332
rect 36228 36320 36234 36372
rect 36817 36363 36875 36369
rect 36817 36329 36829 36363
rect 36863 36360 36875 36363
rect 37182 36360 37188 36372
rect 36863 36332 37188 36360
rect 36863 36329 36875 36332
rect 36817 36323 36875 36329
rect 37182 36320 37188 36332
rect 37240 36320 37246 36372
rect 24302 36252 24308 36304
rect 24360 36292 24366 36304
rect 24489 36295 24547 36301
rect 24489 36292 24501 36295
rect 24360 36264 24501 36292
rect 24360 36252 24366 36264
rect 24489 36261 24501 36264
rect 24535 36292 24547 36295
rect 26145 36295 26203 36301
rect 24535 36264 25084 36292
rect 24535 36261 24547 36264
rect 24489 36255 24547 36261
rect 25056 36233 25084 36264
rect 26145 36261 26157 36295
rect 26191 36292 26203 36295
rect 34790 36292 34796 36304
rect 26191 36264 34796 36292
rect 26191 36261 26203 36264
rect 26145 36255 26203 36261
rect 34790 36252 34796 36264
rect 34848 36252 34854 36304
rect 35345 36295 35403 36301
rect 35345 36261 35357 36295
rect 35391 36292 35403 36295
rect 35391 36264 35848 36292
rect 35391 36261 35403 36264
rect 35345 36255 35403 36261
rect 3988 36196 5212 36224
rect 20809 36227 20867 36233
rect 2774 36156 2780 36168
rect 2735 36128 2780 36156
rect 2774 36116 2780 36128
rect 2832 36116 2838 36168
rect 3988 36165 4016 36196
rect 20809 36193 20821 36227
rect 20855 36193 20867 36227
rect 20809 36187 20867 36193
rect 21637 36227 21695 36233
rect 21637 36193 21649 36227
rect 21683 36224 21695 36227
rect 25041 36227 25099 36233
rect 21683 36196 23980 36224
rect 21683 36193 21695 36196
rect 21637 36187 21695 36193
rect 3973 36159 4031 36165
rect 3973 36125 3985 36159
rect 4019 36125 4031 36159
rect 3973 36119 4031 36125
rect 4617 36159 4675 36165
rect 4617 36125 4629 36159
rect 4663 36156 4675 36159
rect 20625 36159 20683 36165
rect 4663 36128 6914 36156
rect 4663 36125 4675 36128
rect 4617 36119 4675 36125
rect 1854 36088 1860 36100
rect 1767 36060 1860 36088
rect 1854 36048 1860 36060
rect 1912 36088 1918 36100
rect 2866 36088 2872 36100
rect 1912 36060 2872 36088
rect 1912 36048 1918 36060
rect 2866 36048 2872 36060
rect 2924 36048 2930 36100
rect 6886 36088 6914 36128
rect 20625 36125 20637 36159
rect 20671 36156 20683 36159
rect 21450 36156 21456 36168
rect 20671 36128 21456 36156
rect 20671 36125 20683 36128
rect 20625 36119 20683 36125
rect 21450 36116 21456 36128
rect 21508 36116 21514 36168
rect 22281 36159 22339 36165
rect 22281 36125 22293 36159
rect 22327 36125 22339 36159
rect 22462 36156 22468 36168
rect 22423 36128 22468 36156
rect 22281 36119 22339 36125
rect 6886 36060 21404 36088
rect 2590 36020 2596 36032
rect 2551 35992 2596 36020
rect 2590 35980 2596 35992
rect 2648 35980 2654 36032
rect 4154 35980 4160 36032
rect 4212 36020 4218 36032
rect 4433 36023 4491 36029
rect 4433 36020 4445 36023
rect 4212 35992 4445 36020
rect 4212 35980 4218 35992
rect 4433 35989 4445 35992
rect 4479 35989 4491 36023
rect 20438 36020 20444 36032
rect 20399 35992 20444 36020
rect 4433 35983 4491 35989
rect 20438 35980 20444 35992
rect 20496 35980 20502 36032
rect 20530 35980 20536 36032
rect 20588 36020 20594 36032
rect 21269 36023 21327 36029
rect 21269 36020 21281 36023
rect 20588 35992 21281 36020
rect 20588 35980 20594 35992
rect 21269 35989 21281 35992
rect 21315 35989 21327 36023
rect 21376 36020 21404 36060
rect 21910 36048 21916 36100
rect 21968 36088 21974 36100
rect 22296 36088 22324 36119
rect 22462 36116 22468 36128
rect 22520 36116 22526 36168
rect 22925 36091 22983 36097
rect 22925 36088 22937 36091
rect 21968 36060 22937 36088
rect 21968 36048 21974 36060
rect 22925 36057 22937 36060
rect 22971 36057 22983 36091
rect 23952 36088 23980 36196
rect 25041 36193 25053 36227
rect 25087 36193 25099 36227
rect 25041 36187 25099 36193
rect 25409 36227 25467 36233
rect 25409 36193 25421 36227
rect 25455 36224 25467 36227
rect 25455 36196 26234 36224
rect 25455 36193 25467 36196
rect 25409 36187 25467 36193
rect 25225 36159 25283 36165
rect 25225 36125 25237 36159
rect 25271 36156 25283 36159
rect 25498 36156 25504 36168
rect 25271 36128 25504 36156
rect 25271 36125 25283 36128
rect 25225 36119 25283 36125
rect 25498 36116 25504 36128
rect 25556 36116 25562 36168
rect 25958 36156 25964 36168
rect 25919 36128 25964 36156
rect 25958 36116 25964 36128
rect 26016 36116 26022 36168
rect 26206 36156 26234 36196
rect 29730 36184 29736 36236
rect 29788 36224 29794 36236
rect 35820 36233 35848 36264
rect 29917 36227 29975 36233
rect 29917 36224 29929 36227
rect 29788 36196 29929 36224
rect 29788 36184 29794 36196
rect 29917 36193 29929 36196
rect 29963 36193 29975 36227
rect 29917 36187 29975 36193
rect 30285 36227 30343 36233
rect 30285 36193 30297 36227
rect 30331 36224 30343 36227
rect 31113 36227 31171 36233
rect 30331 36196 31064 36224
rect 30331 36193 30343 36196
rect 30285 36187 30343 36193
rect 26605 36159 26663 36165
rect 26605 36156 26617 36159
rect 26206 36128 26617 36156
rect 26605 36125 26617 36128
rect 26651 36125 26663 36159
rect 26605 36119 26663 36125
rect 30006 36116 30012 36168
rect 30064 36156 30070 36168
rect 30101 36159 30159 36165
rect 30101 36156 30113 36159
rect 30064 36128 30113 36156
rect 30064 36116 30070 36128
rect 30101 36125 30113 36128
rect 30147 36125 30159 36159
rect 30742 36156 30748 36168
rect 30703 36128 30748 36156
rect 30101 36119 30159 36125
rect 29822 36088 29828 36100
rect 23952 36060 29828 36088
rect 22925 36051 22983 36057
rect 29822 36048 29828 36060
rect 29880 36048 29886 36100
rect 30116 36088 30144 36119
rect 30742 36116 30748 36128
rect 30800 36116 30806 36168
rect 30929 36159 30987 36165
rect 30929 36125 30941 36159
rect 30975 36125 30987 36159
rect 31036 36156 31064 36196
rect 31113 36193 31125 36227
rect 31159 36224 31171 36227
rect 35805 36227 35863 36233
rect 31159 36196 33640 36224
rect 31159 36193 31171 36196
rect 31113 36187 31171 36193
rect 33612 36165 33640 36196
rect 35805 36193 35817 36227
rect 35851 36193 35863 36227
rect 35805 36187 35863 36193
rect 37277 36227 37335 36233
rect 37277 36193 37289 36227
rect 37323 36224 37335 36227
rect 37366 36224 37372 36236
rect 37323 36196 37372 36224
rect 37323 36193 37335 36196
rect 37277 36187 37335 36193
rect 37366 36184 37372 36196
rect 37424 36184 37430 36236
rect 32953 36159 33011 36165
rect 32953 36156 32965 36159
rect 31036 36128 32965 36156
rect 30929 36119 30987 36125
rect 32953 36125 32965 36128
rect 32999 36125 33011 36159
rect 32953 36119 33011 36125
rect 33597 36159 33655 36165
rect 33597 36125 33609 36159
rect 33643 36125 33655 36159
rect 33597 36119 33655 36125
rect 35161 36159 35219 36165
rect 35161 36125 35173 36159
rect 35207 36156 35219 36159
rect 35526 36156 35532 36168
rect 35207 36128 35532 36156
rect 35207 36125 35219 36128
rect 35161 36119 35219 36125
rect 30944 36088 30972 36119
rect 35526 36116 35532 36128
rect 35584 36116 35590 36168
rect 35986 36156 35992 36168
rect 35899 36128 35992 36156
rect 35986 36116 35992 36128
rect 36044 36156 36050 36168
rect 36354 36156 36360 36168
rect 36044 36128 36360 36156
rect 36044 36116 36050 36128
rect 36354 36116 36360 36128
rect 36412 36116 36418 36168
rect 37553 36159 37611 36165
rect 37553 36125 37565 36159
rect 37599 36125 37611 36159
rect 37553 36119 37611 36125
rect 30116 36060 30972 36088
rect 34514 36048 34520 36100
rect 34572 36088 34578 36100
rect 37568 36088 37596 36119
rect 34572 36060 37596 36088
rect 34572 36048 34578 36060
rect 22097 36023 22155 36029
rect 22097 36020 22109 36023
rect 21376 35992 22109 36020
rect 21269 35983 21327 35989
rect 22097 35989 22109 35992
rect 22143 35989 22155 36023
rect 26786 36020 26792 36032
rect 26747 35992 26792 36020
rect 22097 35983 22155 35989
rect 26786 35980 26792 35992
rect 26844 35980 26850 36032
rect 33137 36023 33195 36029
rect 33137 35989 33149 36023
rect 33183 36020 33195 36023
rect 35434 36020 35440 36032
rect 33183 35992 35440 36020
rect 33183 35989 33195 35992
rect 33137 35983 33195 35989
rect 35434 35980 35440 35992
rect 35492 35980 35498 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 2958 35816 2964 35828
rect 2919 35788 2964 35816
rect 2958 35776 2964 35788
rect 3016 35776 3022 35828
rect 3510 35776 3516 35828
rect 3568 35816 3574 35828
rect 3605 35819 3663 35825
rect 3605 35816 3617 35819
rect 3568 35788 3617 35816
rect 3568 35776 3574 35788
rect 3605 35785 3617 35788
rect 3651 35785 3663 35819
rect 4154 35816 4160 35828
rect 3605 35779 3663 35785
rect 4080 35788 4160 35816
rect 4080 35748 4108 35788
rect 4154 35776 4160 35788
rect 4212 35776 4218 35828
rect 4433 35819 4491 35825
rect 4433 35785 4445 35819
rect 4479 35816 4491 35819
rect 4614 35816 4620 35828
rect 4479 35788 4620 35816
rect 4479 35785 4491 35788
rect 4433 35779 4491 35785
rect 4614 35776 4620 35788
rect 4672 35776 4678 35828
rect 20993 35819 21051 35825
rect 20993 35785 21005 35819
rect 21039 35816 21051 35819
rect 21450 35816 21456 35828
rect 21039 35788 21456 35816
rect 21039 35785 21051 35788
rect 20993 35779 21051 35785
rect 21450 35776 21456 35788
rect 21508 35816 21514 35828
rect 21821 35819 21879 35825
rect 21821 35816 21833 35819
rect 21508 35788 21833 35816
rect 21508 35776 21514 35788
rect 21821 35785 21833 35788
rect 21867 35816 21879 35819
rect 21910 35816 21916 35828
rect 21867 35788 21916 35816
rect 21867 35785 21879 35788
rect 21821 35779 21879 35785
rect 21910 35776 21916 35788
rect 21968 35776 21974 35828
rect 24857 35819 24915 35825
rect 24857 35785 24869 35819
rect 24903 35816 24915 35819
rect 25958 35816 25964 35828
rect 24903 35788 25964 35816
rect 24903 35785 24915 35788
rect 24857 35779 24915 35785
rect 25958 35776 25964 35788
rect 26016 35776 26022 35828
rect 26329 35819 26387 35825
rect 26329 35785 26341 35819
rect 26375 35816 26387 35819
rect 33870 35816 33876 35828
rect 26375 35788 33876 35816
rect 26375 35785 26387 35788
rect 26329 35779 26387 35785
rect 33870 35776 33876 35788
rect 33928 35776 33934 35828
rect 35526 35816 35532 35828
rect 35487 35788 35532 35816
rect 35526 35776 35532 35788
rect 35584 35776 35590 35828
rect 4985 35751 5043 35757
rect 4985 35748 4997 35751
rect 3160 35720 4108 35748
rect 4172 35720 4997 35748
rect 1857 35683 1915 35689
rect 1857 35649 1869 35683
rect 1903 35680 1915 35683
rect 3050 35680 3056 35692
rect 1903 35652 3056 35680
rect 1903 35649 1915 35652
rect 1857 35643 1915 35649
rect 3050 35640 3056 35652
rect 3108 35640 3114 35692
rect 3160 35689 3188 35720
rect 3145 35683 3203 35689
rect 3145 35649 3157 35683
rect 3191 35649 3203 35683
rect 3145 35643 3203 35649
rect 3789 35683 3847 35689
rect 3789 35649 3801 35683
rect 3835 35680 3847 35683
rect 4172 35680 4200 35720
rect 4985 35717 4997 35720
rect 5031 35748 5043 35751
rect 35894 35748 35900 35760
rect 5031 35720 35900 35748
rect 5031 35717 5043 35720
rect 4985 35711 5043 35717
rect 35894 35708 35900 35720
rect 35952 35708 35958 35760
rect 3835 35652 4200 35680
rect 4249 35683 4307 35689
rect 3835 35649 3847 35652
rect 3789 35643 3847 35649
rect 4249 35649 4261 35683
rect 4295 35680 4307 35683
rect 20530 35680 20536 35692
rect 4295 35652 20536 35680
rect 4295 35649 4307 35652
rect 4249 35643 4307 35649
rect 20530 35640 20536 35652
rect 20588 35640 20594 35692
rect 24673 35683 24731 35689
rect 24673 35649 24685 35683
rect 24719 35649 24731 35683
rect 24673 35643 24731 35649
rect 3694 35572 3700 35624
rect 3752 35612 3758 35624
rect 23937 35615 23995 35621
rect 23937 35612 23949 35615
rect 3752 35584 23949 35612
rect 3752 35572 3758 35584
rect 23937 35581 23949 35584
rect 23983 35612 23995 35615
rect 24489 35615 24547 35621
rect 24489 35612 24501 35615
rect 23983 35584 24501 35612
rect 23983 35581 23995 35584
rect 23937 35575 23995 35581
rect 24489 35581 24501 35584
rect 24535 35581 24547 35615
rect 24688 35612 24716 35643
rect 24762 35640 24768 35692
rect 24820 35680 24826 35692
rect 26145 35683 26203 35689
rect 26145 35680 26157 35683
rect 24820 35652 26157 35680
rect 24820 35640 24826 35652
rect 26145 35649 26157 35652
rect 26191 35649 26203 35683
rect 26145 35643 26203 35649
rect 30006 35640 30012 35692
rect 30064 35680 30070 35692
rect 30101 35683 30159 35689
rect 30101 35680 30113 35683
rect 30064 35652 30113 35680
rect 30064 35640 30070 35652
rect 30101 35649 30113 35652
rect 30147 35649 30159 35683
rect 30101 35643 30159 35649
rect 30285 35683 30343 35689
rect 30285 35649 30297 35683
rect 30331 35680 30343 35683
rect 32861 35683 32919 35689
rect 32861 35680 32873 35683
rect 30331 35652 32873 35680
rect 30331 35649 30343 35652
rect 30285 35643 30343 35649
rect 32861 35649 32873 35652
rect 32907 35649 32919 35683
rect 36354 35680 36360 35692
rect 36315 35652 36360 35680
rect 32861 35643 32919 35649
rect 36354 35640 36360 35652
rect 36412 35640 36418 35692
rect 37829 35683 37887 35689
rect 37829 35649 37841 35683
rect 37875 35649 37887 35683
rect 37829 35643 37887 35649
rect 25498 35612 25504 35624
rect 24688 35584 25504 35612
rect 24489 35575 24547 35581
rect 25498 35572 25504 35584
rect 25556 35572 25562 35624
rect 29917 35615 29975 35621
rect 29917 35581 29929 35615
rect 29963 35581 29975 35615
rect 36538 35612 36544 35624
rect 36499 35584 36544 35612
rect 29917 35575 29975 35581
rect 2041 35547 2099 35553
rect 2041 35513 2053 35547
rect 2087 35544 2099 35547
rect 29365 35547 29423 35553
rect 29365 35544 29377 35547
rect 2087 35516 29377 35544
rect 2087 35513 2099 35516
rect 2041 35507 2099 35513
rect 29365 35513 29377 35516
rect 29411 35544 29423 35547
rect 29932 35544 29960 35575
rect 36538 35572 36544 35584
rect 36596 35572 36602 35624
rect 29411 35516 29960 35544
rect 33045 35547 33103 35553
rect 29411 35513 29423 35516
rect 29365 35507 29423 35513
rect 33045 35513 33057 35547
rect 33091 35544 33103 35547
rect 37844 35544 37872 35643
rect 33091 35516 37872 35544
rect 33091 35513 33103 35516
rect 33045 35507 33103 35513
rect 25498 35476 25504 35488
rect 25459 35448 25504 35476
rect 25498 35436 25504 35448
rect 25556 35436 25562 35488
rect 36170 35476 36176 35488
rect 36131 35448 36176 35476
rect 36170 35436 36176 35448
rect 36228 35436 36234 35488
rect 37182 35436 37188 35488
rect 37240 35476 37246 35488
rect 37277 35479 37335 35485
rect 37277 35476 37289 35479
rect 37240 35448 37289 35476
rect 37240 35436 37246 35448
rect 37277 35445 37289 35448
rect 37323 35445 37335 35479
rect 38010 35476 38016 35488
rect 37971 35448 38016 35476
rect 37277 35439 37335 35445
rect 38010 35436 38016 35448
rect 38068 35436 38074 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 2774 35232 2780 35284
rect 2832 35272 2838 35284
rect 2961 35275 3019 35281
rect 2961 35272 2973 35275
rect 2832 35244 2973 35272
rect 2832 35232 2838 35244
rect 2961 35241 2973 35244
rect 3007 35241 3019 35275
rect 3970 35272 3976 35284
rect 3931 35244 3976 35272
rect 2961 35235 3019 35241
rect 3970 35232 3976 35244
rect 4028 35232 4034 35284
rect 36538 35272 36544 35284
rect 36499 35244 36544 35272
rect 36538 35232 36544 35244
rect 36596 35232 36602 35284
rect 35529 35207 35587 35213
rect 35529 35173 35541 35207
rect 35575 35204 35587 35207
rect 37366 35204 37372 35216
rect 35575 35176 37372 35204
rect 35575 35173 35587 35176
rect 35529 35167 35587 35173
rect 37366 35164 37372 35176
rect 37424 35164 37430 35216
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35068 1731 35071
rect 2409 35071 2467 35077
rect 1719 35040 2360 35068
rect 1719 35037 1731 35040
rect 1673 35031 1731 35037
rect 1486 34932 1492 34944
rect 1447 34904 1492 34932
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 2222 34932 2228 34944
rect 2183 34904 2228 34932
rect 2222 34892 2228 34904
rect 2280 34892 2286 34944
rect 2332 34932 2360 35040
rect 2409 35037 2421 35071
rect 2455 35068 2467 35071
rect 2682 35068 2688 35080
rect 2455 35040 2688 35068
rect 2455 35037 2467 35040
rect 2409 35031 2467 35037
rect 2682 35028 2688 35040
rect 2740 35028 2746 35080
rect 3145 35071 3203 35077
rect 3145 35037 3157 35071
rect 3191 35037 3203 35071
rect 3145 35031 3203 35037
rect 3789 35071 3847 35077
rect 3789 35037 3801 35071
rect 3835 35068 3847 35071
rect 20438 35068 20444 35080
rect 3835 35040 20444 35068
rect 3835 35037 3847 35040
rect 3789 35031 3847 35037
rect 3160 35000 3188 35031
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 36081 35071 36139 35077
rect 36081 35037 36093 35071
rect 36127 35068 36139 35071
rect 36722 35068 36728 35080
rect 36127 35040 36728 35068
rect 36127 35037 36139 35040
rect 36081 35031 36139 35037
rect 36722 35028 36728 35040
rect 36780 35028 36786 35080
rect 37182 35028 37188 35080
rect 37240 35068 37246 35080
rect 37369 35071 37427 35077
rect 37369 35068 37381 35071
rect 37240 35040 37381 35068
rect 37240 35028 37246 35040
rect 37369 35037 37381 35040
rect 37415 35037 37427 35071
rect 37369 35031 37427 35037
rect 37829 35071 37887 35077
rect 37829 35037 37841 35071
rect 37875 35037 37887 35071
rect 37829 35031 37887 35037
rect 3970 35000 3976 35012
rect 3160 34972 3976 35000
rect 3970 34960 3976 34972
rect 4028 35000 4034 35012
rect 36170 35000 36176 35012
rect 4028 34972 36176 35000
rect 4028 34960 4034 34972
rect 36170 34960 36176 34972
rect 36228 34960 36234 35012
rect 36814 34960 36820 35012
rect 36872 35000 36878 35012
rect 37844 35000 37872 35031
rect 36872 34972 37872 35000
rect 36872 34960 36878 34972
rect 4525 34935 4583 34941
rect 4525 34932 4537 34935
rect 2332 34904 4537 34932
rect 4525 34901 4537 34904
rect 4571 34932 4583 34935
rect 4614 34932 4620 34944
rect 4571 34904 4620 34932
rect 4571 34901 4583 34904
rect 4525 34895 4583 34901
rect 4614 34892 4620 34904
rect 4672 34892 4678 34944
rect 25041 34935 25099 34941
rect 25041 34901 25053 34935
rect 25087 34932 25099 34935
rect 25498 34932 25504 34944
rect 25087 34904 25504 34932
rect 25087 34901 25099 34904
rect 25041 34895 25099 34901
rect 25498 34892 25504 34904
rect 25556 34892 25562 34944
rect 37185 34935 37243 34941
rect 37185 34901 37197 34935
rect 37231 34932 37243 34935
rect 37274 34932 37280 34944
rect 37231 34904 37280 34932
rect 37231 34901 37243 34904
rect 37185 34895 37243 34901
rect 37274 34892 37280 34904
rect 37332 34892 37338 34944
rect 38010 34932 38016 34944
rect 37971 34904 38016 34932
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2682 34728 2688 34740
rect 2643 34700 2688 34728
rect 2682 34688 2688 34700
rect 2740 34688 2746 34740
rect 3970 34728 3976 34740
rect 3931 34700 3976 34728
rect 3970 34688 3976 34700
rect 4028 34688 4034 34740
rect 37645 34731 37703 34737
rect 37645 34728 37657 34731
rect 29932 34700 37657 34728
rect 2041 34663 2099 34669
rect 2041 34629 2053 34663
rect 2087 34660 2099 34663
rect 29273 34663 29331 34669
rect 29273 34660 29285 34663
rect 2087 34632 29285 34660
rect 2087 34629 2099 34632
rect 2041 34623 2099 34629
rect 29273 34629 29285 34632
rect 29319 34660 29331 34663
rect 29319 34632 29868 34660
rect 29319 34629 29331 34632
rect 29273 34623 29331 34629
rect 1854 34592 1860 34604
rect 1815 34564 1860 34592
rect 1854 34552 1860 34564
rect 1912 34552 1918 34604
rect 29840 34601 29868 34632
rect 2869 34595 2927 34601
rect 2869 34561 2881 34595
rect 2915 34592 2927 34595
rect 3421 34595 3479 34601
rect 3421 34592 3433 34595
rect 2915 34564 3433 34592
rect 2915 34561 2927 34564
rect 2869 34555 2927 34561
rect 3421 34561 3433 34564
rect 3467 34592 3479 34595
rect 29825 34595 29883 34601
rect 3467 34564 26234 34592
rect 3467 34561 3479 34564
rect 3421 34555 3479 34561
rect 26206 34524 26234 34564
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 29932 34524 29960 34700
rect 37645 34697 37657 34700
rect 37691 34697 37703 34731
rect 37645 34691 37703 34697
rect 36725 34663 36783 34669
rect 36725 34629 36737 34663
rect 36771 34660 36783 34663
rect 37366 34660 37372 34672
rect 36771 34632 37372 34660
rect 36771 34629 36783 34632
rect 36725 34623 36783 34629
rect 37366 34620 37372 34632
rect 37424 34620 37430 34672
rect 30006 34552 30012 34604
rect 30064 34592 30070 34604
rect 30193 34595 30251 34601
rect 30064 34564 30109 34592
rect 30064 34552 30070 34564
rect 30193 34561 30205 34595
rect 30239 34592 30251 34595
rect 32125 34595 32183 34601
rect 32125 34592 32137 34595
rect 30239 34564 32137 34592
rect 30239 34561 30251 34564
rect 30193 34555 30251 34561
rect 32125 34561 32137 34564
rect 32171 34561 32183 34595
rect 37274 34592 37280 34604
rect 37235 34564 37280 34592
rect 32125 34555 32183 34561
rect 37274 34552 37280 34564
rect 37332 34552 37338 34604
rect 37461 34595 37519 34601
rect 37461 34592 37473 34595
rect 37384 34564 37473 34592
rect 36814 34524 36820 34536
rect 26206 34496 29960 34524
rect 32324 34496 36820 34524
rect 32324 34465 32352 34496
rect 36814 34484 36820 34496
rect 36872 34484 36878 34536
rect 32309 34459 32367 34465
rect 32309 34425 32321 34459
rect 32355 34425 32367 34459
rect 32309 34419 32367 34425
rect 36354 34416 36360 34468
rect 36412 34456 36418 34468
rect 37384 34456 37412 34564
rect 37461 34561 37473 34564
rect 37507 34561 37519 34595
rect 37461 34555 37519 34561
rect 36412 34428 37412 34456
rect 36412 34416 36418 34428
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 3050 34184 3056 34196
rect 3011 34156 3056 34184
rect 3050 34144 3056 34156
rect 3108 34144 3114 34196
rect 37185 34119 37243 34125
rect 37185 34116 37197 34119
rect 35866 34088 37197 34116
rect 35437 34051 35495 34057
rect 35437 34017 35449 34051
rect 35483 34048 35495 34051
rect 35866 34048 35894 34088
rect 37185 34085 37197 34088
rect 37231 34085 37243 34119
rect 37185 34079 37243 34085
rect 35483 34020 35894 34048
rect 35483 34017 35495 34020
rect 35437 34011 35495 34017
rect 2041 33983 2099 33989
rect 2041 33949 2053 33983
rect 2087 33980 2099 33983
rect 29270 33980 29276 33992
rect 2087 33952 29276 33980
rect 2087 33949 2099 33952
rect 2041 33943 2099 33949
rect 29270 33940 29276 33952
rect 29328 33940 29334 33992
rect 35253 33983 35311 33989
rect 35253 33949 35265 33983
rect 35299 33980 35311 33983
rect 35342 33980 35348 33992
rect 35299 33952 35348 33980
rect 35299 33949 35311 33952
rect 35253 33943 35311 33949
rect 35342 33940 35348 33952
rect 35400 33980 35406 33992
rect 36354 33980 36360 33992
rect 35400 33952 36360 33980
rect 35400 33940 35406 33952
rect 36354 33940 36360 33952
rect 36412 33940 36418 33992
rect 36725 33983 36783 33989
rect 36725 33949 36737 33983
rect 36771 33980 36783 33983
rect 37366 33980 37372 33992
rect 36771 33952 37372 33980
rect 36771 33949 36783 33952
rect 36725 33943 36783 33949
rect 37366 33940 37372 33952
rect 37424 33940 37430 33992
rect 37826 33980 37832 33992
rect 37787 33952 37832 33980
rect 37826 33940 37832 33952
rect 37884 33940 37890 33992
rect 1854 33912 1860 33924
rect 1815 33884 1860 33912
rect 1854 33872 1860 33884
rect 1912 33912 1918 33924
rect 2501 33915 2559 33921
rect 2501 33912 2513 33915
rect 1912 33884 2513 33912
rect 1912 33872 1918 33884
rect 2501 33881 2513 33884
rect 2547 33881 2559 33915
rect 2501 33875 2559 33881
rect 34057 33915 34115 33921
rect 34057 33881 34069 33915
rect 34103 33912 34115 33915
rect 35069 33915 35127 33921
rect 35069 33912 35081 33915
rect 34103 33884 35081 33912
rect 34103 33881 34115 33884
rect 34057 33875 34115 33881
rect 35069 33881 35081 33884
rect 35115 33881 35127 33915
rect 35069 33875 35127 33881
rect 4614 33804 4620 33856
rect 4672 33844 4678 33856
rect 33965 33847 34023 33853
rect 33965 33844 33977 33847
rect 4672 33816 33977 33844
rect 4672 33804 4678 33816
rect 33965 33813 33977 33816
rect 34011 33813 34023 33847
rect 38010 33844 38016 33856
rect 37971 33816 38016 33844
rect 33965 33807 34023 33813
rect 38010 33804 38016 33816
rect 38068 33804 38074 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1946 33600 1952 33652
rect 2004 33640 2010 33652
rect 2133 33643 2191 33649
rect 2133 33640 2145 33643
rect 2004 33612 2145 33640
rect 2004 33600 2010 33612
rect 2133 33609 2145 33612
rect 2179 33609 2191 33643
rect 29270 33640 29276 33652
rect 29231 33612 29276 33640
rect 2133 33603 2191 33609
rect 29270 33600 29276 33612
rect 29328 33600 29334 33652
rect 32309 33643 32367 33649
rect 32309 33609 32321 33643
rect 32355 33640 32367 33643
rect 37826 33640 37832 33652
rect 32355 33612 37832 33640
rect 32355 33609 32367 33612
rect 32309 33603 32367 33609
rect 37826 33600 37832 33612
rect 37884 33600 37890 33652
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 2682 33504 2688 33516
rect 1719 33476 2688 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 2682 33464 2688 33476
rect 2740 33464 2746 33516
rect 29288 33504 29316 33600
rect 29825 33507 29883 33513
rect 29825 33504 29837 33507
rect 29288 33476 29837 33504
rect 29825 33473 29837 33476
rect 29871 33473 29883 33507
rect 30006 33504 30012 33516
rect 29967 33476 30012 33504
rect 29825 33467 29883 33473
rect 30006 33464 30012 33476
rect 30064 33464 30070 33516
rect 30193 33507 30251 33513
rect 30193 33473 30205 33507
rect 30239 33504 30251 33507
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 30239 33476 32137 33504
rect 30239 33473 30251 33476
rect 30193 33467 30251 33473
rect 32125 33473 32137 33476
rect 32171 33473 32183 33507
rect 37826 33504 37832 33516
rect 37787 33476 37832 33504
rect 32125 33467 32183 33473
rect 37826 33464 37832 33476
rect 37884 33464 37890 33516
rect 37369 33371 37427 33377
rect 37369 33337 37381 33371
rect 37415 33368 37427 33371
rect 38102 33368 38108 33380
rect 37415 33340 38108 33368
rect 37415 33337 37427 33340
rect 37369 33331 37427 33337
rect 38102 33328 38108 33340
rect 38160 33328 38166 33380
rect 1486 33300 1492 33312
rect 1447 33272 1492 33300
rect 1486 33260 1492 33272
rect 1544 33260 1550 33312
rect 38010 33300 38016 33312
rect 37971 33272 38016 33300
rect 38010 33260 38016 33272
rect 38068 33260 38074 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 35342 33056 35348 33108
rect 35400 33096 35406 33108
rect 35437 33099 35495 33105
rect 35437 33096 35449 33099
rect 35400 33068 35449 33096
rect 35400 33056 35406 33068
rect 35437 33065 35449 33068
rect 35483 33065 35495 33099
rect 35437 33059 35495 33065
rect 36262 32988 36268 33040
rect 36320 33028 36326 33040
rect 37921 33031 37979 33037
rect 37921 33028 37933 33031
rect 36320 33000 37933 33028
rect 36320 32988 36326 33000
rect 37921 32997 37933 33000
rect 37967 32997 37979 33031
rect 37921 32991 37979 32997
rect 2501 32895 2559 32901
rect 2501 32861 2513 32895
rect 2547 32892 2559 32895
rect 2774 32892 2780 32904
rect 2547 32864 2780 32892
rect 2547 32861 2559 32864
rect 2501 32855 2559 32861
rect 2774 32852 2780 32864
rect 2832 32892 2838 32904
rect 3145 32895 3203 32901
rect 3145 32892 3157 32895
rect 2832 32864 3157 32892
rect 2832 32852 2838 32864
rect 3145 32861 3157 32864
rect 3191 32861 3203 32895
rect 3145 32855 3203 32861
rect 26050 32852 26056 32904
rect 26108 32892 26114 32904
rect 26973 32895 27031 32901
rect 26973 32892 26985 32895
rect 26108 32864 26985 32892
rect 26108 32852 26114 32864
rect 26973 32861 26985 32864
rect 27019 32861 27031 32895
rect 26973 32855 27031 32861
rect 35253 32895 35311 32901
rect 35253 32861 35265 32895
rect 35299 32892 35311 32895
rect 35802 32892 35808 32904
rect 35299 32864 35808 32892
rect 35299 32861 35311 32864
rect 35253 32855 35311 32861
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 36817 32895 36875 32901
rect 36817 32861 36829 32895
rect 36863 32892 36875 32895
rect 37458 32892 37464 32904
rect 36863 32864 37464 32892
rect 36863 32861 36875 32864
rect 36817 32855 36875 32861
rect 37458 32852 37464 32864
rect 37516 32852 37522 32904
rect 38102 32892 38108 32904
rect 38063 32864 38108 32892
rect 38102 32852 38108 32864
rect 38160 32852 38166 32904
rect 1854 32824 1860 32836
rect 1815 32796 1860 32824
rect 1854 32784 1860 32796
rect 1912 32784 1918 32836
rect 37826 32824 37832 32836
rect 27172 32796 37832 32824
rect 1946 32756 1952 32768
rect 1907 32728 1952 32756
rect 1946 32716 1952 32728
rect 2004 32716 2010 32768
rect 2685 32759 2743 32765
rect 2685 32725 2697 32759
rect 2731 32756 2743 32759
rect 6178 32756 6184 32768
rect 2731 32728 6184 32756
rect 2731 32725 2743 32728
rect 2685 32719 2743 32725
rect 6178 32716 6184 32728
rect 6236 32716 6242 32768
rect 27172 32765 27200 32796
rect 37826 32784 37832 32796
rect 37884 32784 37890 32836
rect 27157 32759 27215 32765
rect 27157 32725 27169 32759
rect 27203 32725 27215 32759
rect 27157 32719 27215 32725
rect 35802 32716 35808 32768
rect 35860 32756 35866 32768
rect 35897 32759 35955 32765
rect 35897 32756 35909 32759
rect 35860 32728 35909 32756
rect 35860 32716 35866 32728
rect 35897 32725 35909 32728
rect 35943 32725 35955 32759
rect 37274 32756 37280 32768
rect 37235 32728 37280 32756
rect 35897 32719 35955 32725
rect 37274 32716 37280 32728
rect 37332 32716 37338 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1946 32512 1952 32564
rect 2004 32552 2010 32564
rect 25133 32555 25191 32561
rect 25133 32552 25145 32555
rect 2004 32524 25145 32552
rect 2004 32512 2010 32524
rect 25133 32521 25145 32524
rect 25179 32552 25191 32555
rect 26050 32552 26056 32564
rect 25179 32524 25728 32552
rect 26011 32524 26056 32552
rect 25179 32521 25191 32524
rect 25133 32515 25191 32521
rect 1854 32444 1860 32496
rect 1912 32484 1918 32496
rect 2133 32487 2191 32493
rect 2133 32484 2145 32487
rect 1912 32456 2145 32484
rect 1912 32444 1918 32456
rect 2133 32453 2145 32456
rect 2179 32453 2191 32487
rect 2133 32447 2191 32453
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 25700 32425 25728 32524
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 29273 32555 29331 32561
rect 29273 32521 29285 32555
rect 29319 32552 29331 32555
rect 30006 32552 30012 32564
rect 29319 32524 30012 32552
rect 29319 32521 29331 32524
rect 29273 32515 29331 32521
rect 30006 32512 30012 32524
rect 30064 32512 30070 32564
rect 2869 32419 2927 32425
rect 2869 32385 2881 32419
rect 2915 32416 2927 32419
rect 25685 32419 25743 32425
rect 2915 32388 3464 32416
rect 2915 32385 2927 32388
rect 2869 32379 2927 32385
rect 2682 32280 2688 32292
rect 2643 32252 2688 32280
rect 2682 32240 2688 32252
rect 2740 32240 2746 32292
rect 3436 32289 3464 32388
rect 25685 32385 25697 32419
rect 25731 32385 25743 32419
rect 25685 32379 25743 32385
rect 25869 32419 25927 32425
rect 25869 32385 25881 32419
rect 25915 32416 25927 32419
rect 26234 32416 26240 32428
rect 25915 32388 26240 32416
rect 25915 32385 25927 32388
rect 25869 32379 25927 32385
rect 26234 32376 26240 32388
rect 26292 32376 26298 32428
rect 28718 32376 28724 32428
rect 28776 32416 28782 32428
rect 29089 32419 29147 32425
rect 29089 32416 29101 32419
rect 28776 32388 29101 32416
rect 28776 32376 28782 32388
rect 29089 32385 29101 32388
rect 29135 32416 29147 32419
rect 29733 32419 29791 32425
rect 29733 32416 29745 32419
rect 29135 32388 29745 32416
rect 29135 32385 29147 32388
rect 29089 32379 29147 32385
rect 29733 32385 29745 32388
rect 29779 32385 29791 32419
rect 37274 32416 37280 32428
rect 37235 32388 37280 32416
rect 29733 32379 29791 32385
rect 37274 32376 37280 32388
rect 37332 32376 37338 32428
rect 37461 32419 37519 32425
rect 37461 32385 37473 32419
rect 37507 32416 37519 32419
rect 37642 32416 37648 32428
rect 37507 32388 37648 32416
rect 37507 32385 37519 32388
rect 37461 32379 37519 32385
rect 37642 32376 37648 32388
rect 37700 32376 37706 32428
rect 3510 32308 3516 32360
rect 3568 32348 3574 32360
rect 25406 32348 25412 32360
rect 3568 32320 25412 32348
rect 3568 32308 3574 32320
rect 25406 32308 25412 32320
rect 25464 32308 25470 32360
rect 3421 32283 3479 32289
rect 3421 32249 3433 32283
rect 3467 32280 3479 32283
rect 37645 32283 37703 32289
rect 37645 32280 37657 32283
rect 3467 32252 37657 32280
rect 3467 32249 3479 32252
rect 3421 32243 3479 32249
rect 37645 32249 37657 32252
rect 37691 32249 37703 32283
rect 37645 32243 37703 32249
rect 1486 32212 1492 32224
rect 1447 32184 1492 32212
rect 1486 32172 1492 32184
rect 1544 32172 1550 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1949 32011 2007 32017
rect 1949 31977 1961 32011
rect 1995 32008 2007 32011
rect 3510 32008 3516 32020
rect 1995 31980 3516 32008
rect 1995 31977 2007 31980
rect 1949 31971 2007 31977
rect 3510 31968 3516 31980
rect 3568 31968 3574 32020
rect 33781 32011 33839 32017
rect 33781 32008 33793 32011
rect 6886 31980 33793 32008
rect 1670 31900 1676 31952
rect 1728 31940 1734 31952
rect 3145 31943 3203 31949
rect 3145 31940 3157 31943
rect 1728 31912 3157 31940
rect 1728 31900 1734 31912
rect 3145 31909 3157 31912
rect 3191 31940 3203 31943
rect 6886 31940 6914 31980
rect 33781 31977 33793 31980
rect 33827 31977 33839 32011
rect 38010 32008 38016 32020
rect 33781 31971 33839 31977
rect 35866 31980 37872 32008
rect 37971 31980 38016 32008
rect 25406 31940 25412 31952
rect 3191 31912 6914 31940
rect 25367 31912 25412 31940
rect 3191 31909 3203 31912
rect 3145 31903 3203 31909
rect 25406 31900 25412 31912
rect 25464 31900 25470 31952
rect 35866 31940 35894 31980
rect 37274 31940 37280 31952
rect 26206 31912 35894 31940
rect 37235 31912 37280 31940
rect 23201 31875 23259 31881
rect 23201 31841 23213 31875
rect 23247 31872 23259 31875
rect 26206 31872 26234 31912
rect 37274 31900 37280 31912
rect 37332 31900 37338 31952
rect 23247 31844 26234 31872
rect 27724 31844 37136 31872
rect 23247 31841 23259 31844
rect 23201 31835 23259 31841
rect 1854 31804 1860 31816
rect 1815 31776 1860 31804
rect 1854 31764 1860 31776
rect 1912 31804 1918 31816
rect 2501 31807 2559 31813
rect 2501 31804 2513 31807
rect 1912 31776 2513 31804
rect 1912 31764 1918 31776
rect 2501 31773 2513 31776
rect 2547 31773 2559 31807
rect 7650 31804 7656 31816
rect 7611 31776 7656 31804
rect 2501 31767 2559 31773
rect 7650 31764 7656 31776
rect 7708 31764 7714 31816
rect 11974 31804 11980 31816
rect 11935 31776 11980 31804
rect 11974 31764 11980 31776
rect 12032 31764 12038 31816
rect 16577 31807 16635 31813
rect 16577 31773 16589 31807
rect 16623 31804 16635 31807
rect 17402 31804 17408 31816
rect 16623 31776 17408 31804
rect 16623 31773 16635 31776
rect 16577 31767 16635 31773
rect 17402 31764 17408 31776
rect 17460 31804 17466 31816
rect 18417 31807 18475 31813
rect 18417 31804 18429 31807
rect 17460 31776 18429 31804
rect 17460 31764 17466 31776
rect 18417 31773 18429 31776
rect 18463 31773 18475 31807
rect 18417 31767 18475 31773
rect 19058 31764 19064 31816
rect 19116 31804 19122 31816
rect 21453 31807 21511 31813
rect 21453 31804 21465 31807
rect 19116 31776 21465 31804
rect 19116 31764 19122 31776
rect 21453 31773 21465 31776
rect 21499 31773 21511 31807
rect 21453 31767 21511 31773
rect 21637 31807 21695 31813
rect 21637 31773 21649 31807
rect 21683 31773 21695 31807
rect 21637 31767 21695 31773
rect 21821 31807 21879 31813
rect 21821 31773 21833 31807
rect 21867 31804 21879 31807
rect 22925 31807 22983 31813
rect 22925 31804 22937 31807
rect 21867 31776 22937 31804
rect 21867 31773 21879 31776
rect 21821 31767 21879 31773
rect 22925 31773 22937 31776
rect 22971 31773 22983 31807
rect 22925 31767 22983 31773
rect 16850 31745 16856 31748
rect 16844 31699 16856 31745
rect 16908 31736 16914 31748
rect 21652 31736 21680 31767
rect 25406 31764 25412 31816
rect 25464 31804 25470 31816
rect 25961 31807 26019 31813
rect 25961 31804 25973 31807
rect 25464 31776 25973 31804
rect 25464 31764 25470 31776
rect 25961 31773 25973 31776
rect 26007 31773 26019 31807
rect 25961 31767 26019 31773
rect 26145 31807 26203 31813
rect 26145 31773 26157 31807
rect 26191 31804 26203 31807
rect 26234 31804 26240 31816
rect 26191 31776 26240 31804
rect 26191 31773 26203 31776
rect 26145 31767 26203 31773
rect 26234 31764 26240 31776
rect 26292 31764 26298 31816
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31804 26387 31807
rect 27525 31807 27583 31813
rect 27525 31804 27537 31807
rect 26375 31776 27537 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 27525 31773 27537 31776
rect 27571 31773 27583 31807
rect 27525 31767 27583 31773
rect 16908 31708 16944 31736
rect 21008 31708 21680 31736
rect 16850 31696 16856 31699
rect 16908 31696 16914 31708
rect 21008 31680 21036 31708
rect 7282 31628 7288 31680
rect 7340 31668 7346 31680
rect 7469 31671 7527 31677
rect 7469 31668 7481 31671
rect 7340 31640 7481 31668
rect 7340 31628 7346 31640
rect 7469 31637 7481 31640
rect 7515 31637 7527 31671
rect 7469 31631 7527 31637
rect 11793 31671 11851 31677
rect 11793 31637 11805 31671
rect 11839 31668 11851 31671
rect 11882 31668 11888 31680
rect 11839 31640 11888 31668
rect 11839 31637 11851 31640
rect 11793 31631 11851 31637
rect 11882 31628 11888 31640
rect 11940 31628 11946 31680
rect 17954 31668 17960 31680
rect 17915 31640 17960 31668
rect 17954 31628 17960 31640
rect 18012 31628 18018 31680
rect 20990 31668 20996 31680
rect 20951 31640 20996 31668
rect 20990 31628 20996 31640
rect 21048 31628 21054 31680
rect 27724 31677 27752 31844
rect 33873 31807 33931 31813
rect 33873 31773 33885 31807
rect 33919 31804 33931 31807
rect 35894 31804 35900 31816
rect 33919 31776 35900 31804
rect 33919 31773 33931 31776
rect 33873 31767 33931 31773
rect 35894 31764 35900 31776
rect 35952 31764 35958 31816
rect 37108 31813 37136 31844
rect 37844 31813 37872 31980
rect 38010 31968 38016 31980
rect 38068 31968 38074 32020
rect 37093 31807 37151 31813
rect 37093 31773 37105 31807
rect 37139 31773 37151 31807
rect 37093 31767 37151 31773
rect 37829 31807 37887 31813
rect 37829 31773 37841 31807
rect 37875 31773 37887 31807
rect 37829 31767 37887 31773
rect 27709 31671 27767 31677
rect 27709 31637 27721 31671
rect 27755 31637 27767 31671
rect 27709 31631 27767 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 2317 31467 2375 31473
rect 2317 31433 2329 31467
rect 2363 31464 2375 31467
rect 7377 31467 7435 31473
rect 2363 31436 6914 31464
rect 2363 31433 2375 31436
rect 2317 31427 2375 31433
rect 6886 31396 6914 31436
rect 7377 31433 7389 31467
rect 7423 31464 7435 31467
rect 7650 31464 7656 31476
rect 7423 31436 7656 31464
rect 7423 31433 7435 31436
rect 7377 31427 7435 31433
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 16850 31464 16856 31476
rect 16811 31436 16856 31464
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 26234 31424 26240 31476
rect 26292 31464 26298 31476
rect 26973 31467 27031 31473
rect 26973 31464 26985 31467
rect 26292 31436 26985 31464
rect 26292 31424 26298 31436
rect 26973 31433 26985 31436
rect 27019 31464 27031 31467
rect 27154 31464 27160 31476
rect 27019 31436 27160 31464
rect 27019 31433 27031 31436
rect 26973 31427 27031 31433
rect 27154 31424 27160 31436
rect 27212 31424 27218 31476
rect 35894 31424 35900 31476
rect 35952 31464 35958 31476
rect 35952 31436 35997 31464
rect 35952 31424 35958 31436
rect 12342 31396 12348 31408
rect 6886 31368 12348 31396
rect 12342 31356 12348 31368
rect 12400 31356 12406 31408
rect 1673 31331 1731 31337
rect 1673 31297 1685 31331
rect 1719 31297 1731 31331
rect 2130 31328 2136 31340
rect 2091 31300 2136 31328
rect 1673 31291 1731 31297
rect 1688 31260 1716 31291
rect 2130 31288 2136 31300
rect 2188 31328 2194 31340
rect 2777 31331 2835 31337
rect 2777 31328 2789 31331
rect 2188 31300 2789 31328
rect 2188 31288 2194 31300
rect 2777 31297 2789 31300
rect 2823 31297 2835 31331
rect 7742 31328 7748 31340
rect 7703 31300 7748 31328
rect 2777 31291 2835 31297
rect 7742 31288 7748 31300
rect 7800 31288 7806 31340
rect 11882 31337 11888 31340
rect 11876 31328 11888 31337
rect 11843 31300 11888 31328
rect 11876 31291 11888 31300
rect 11882 31288 11888 31291
rect 11940 31288 11946 31340
rect 16482 31288 16488 31340
rect 16540 31328 16546 31340
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16540 31300 16681 31328
rect 16540 31288 16546 31300
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21048 31300 22017 31328
rect 21048 31288 21054 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 27157 31331 27215 31337
rect 27157 31297 27169 31331
rect 27203 31328 27215 31331
rect 27706 31328 27712 31340
rect 27203 31300 27712 31328
rect 27203 31297 27215 31300
rect 27157 31291 27215 31297
rect 27706 31288 27712 31300
rect 27764 31288 27770 31340
rect 36078 31328 36084 31340
rect 36039 31300 36084 31328
rect 36078 31288 36084 31300
rect 36136 31288 36142 31340
rect 37829 31331 37887 31337
rect 37829 31328 37841 31331
rect 36188 31300 37841 31328
rect 1688 31232 3464 31260
rect 1486 31124 1492 31136
rect 1447 31096 1492 31124
rect 1486 31084 1492 31096
rect 1544 31084 1550 31136
rect 3436 31133 3464 31232
rect 6178 31220 6184 31272
rect 6236 31260 6242 31272
rect 7837 31263 7895 31269
rect 7837 31260 7849 31263
rect 6236 31232 7849 31260
rect 6236 31220 6242 31232
rect 7837 31229 7849 31232
rect 7883 31229 7895 31263
rect 8018 31260 8024 31272
rect 7979 31232 8024 31260
rect 7837 31223 7895 31229
rect 8018 31220 8024 31232
rect 8076 31260 8082 31272
rect 8573 31263 8631 31269
rect 8573 31260 8585 31263
rect 8076 31232 8585 31260
rect 8076 31220 8082 31232
rect 8573 31229 8585 31232
rect 8619 31229 8631 31263
rect 8573 31223 8631 31229
rect 9030 31220 9036 31272
rect 9088 31260 9094 31272
rect 10965 31263 11023 31269
rect 10965 31260 10977 31263
rect 9088 31232 10977 31260
rect 9088 31220 9094 31232
rect 10965 31229 10977 31232
rect 11011 31260 11023 31263
rect 11609 31263 11667 31269
rect 11609 31260 11621 31263
rect 11011 31232 11621 31260
rect 11011 31229 11023 31232
rect 10965 31223 11023 31229
rect 11609 31229 11621 31232
rect 11655 31229 11667 31263
rect 21821 31263 21879 31269
rect 21821 31260 21833 31263
rect 11609 31223 11667 31229
rect 13004 31232 21833 31260
rect 13004 31204 13032 31232
rect 21821 31229 21833 31232
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31260 22247 31263
rect 23109 31263 23167 31269
rect 23109 31260 23121 31263
rect 22235 31232 23121 31260
rect 22235 31229 22247 31232
rect 22189 31223 22247 31229
rect 23109 31229 23121 31232
rect 23155 31229 23167 31263
rect 23109 31223 23167 31229
rect 23385 31263 23443 31269
rect 23385 31229 23397 31263
rect 23431 31260 23443 31263
rect 36188 31260 36216 31300
rect 37829 31297 37841 31300
rect 37875 31297 37887 31331
rect 37829 31291 37887 31297
rect 23431 31232 36216 31260
rect 23431 31229 23443 31232
rect 23385 31223 23443 31229
rect 36262 31220 36268 31272
rect 36320 31260 36326 31272
rect 36320 31232 36365 31260
rect 36320 31220 36326 31232
rect 12986 31192 12992 31204
rect 12899 31164 12992 31192
rect 12986 31152 12992 31164
rect 13044 31152 13050 31204
rect 3421 31127 3479 31133
rect 3421 31093 3433 31127
rect 3467 31124 3479 31127
rect 8478 31124 8484 31136
rect 3467 31096 8484 31124
rect 3467 31093 3479 31096
rect 3421 31087 3479 31093
rect 8478 31084 8484 31096
rect 8536 31084 8542 31136
rect 20990 31084 20996 31136
rect 21048 31124 21054 31136
rect 21177 31127 21235 31133
rect 21177 31124 21189 31127
rect 21048 31096 21189 31124
rect 21048 31084 21054 31096
rect 21177 31093 21189 31096
rect 21223 31093 21235 31127
rect 27706 31124 27712 31136
rect 27619 31096 27712 31124
rect 21177 31087 21235 31093
rect 27706 31084 27712 31096
rect 27764 31124 27770 31136
rect 28718 31124 28724 31136
rect 27764 31096 28724 31124
rect 27764 31084 27770 31096
rect 28718 31084 28724 31096
rect 28776 31084 28782 31136
rect 38010 31124 38016 31136
rect 37971 31096 38016 31124
rect 38010 31084 38016 31096
rect 38068 31084 38074 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 9030 30920 9036 30932
rect 7024 30892 9036 30920
rect 7024 30793 7052 30892
rect 9030 30880 9036 30892
rect 9088 30880 9094 30932
rect 11885 30923 11943 30929
rect 11885 30889 11897 30923
rect 11931 30920 11943 30923
rect 11974 30920 11980 30932
rect 11931 30892 11980 30920
rect 11931 30889 11943 30892
rect 11885 30883 11943 30889
rect 11974 30880 11980 30892
rect 12032 30880 12038 30932
rect 33781 30923 33839 30929
rect 33781 30920 33793 30923
rect 12084 30892 33793 30920
rect 8478 30812 8484 30864
rect 8536 30852 8542 30864
rect 12084 30852 12112 30892
rect 33781 30889 33793 30892
rect 33827 30889 33839 30923
rect 33781 30883 33839 30889
rect 35805 30923 35863 30929
rect 35805 30889 35817 30923
rect 35851 30920 35863 30923
rect 36078 30920 36084 30932
rect 35851 30892 36084 30920
rect 35851 30889 35863 30892
rect 35805 30883 35863 30889
rect 36078 30880 36084 30892
rect 36136 30920 36142 30932
rect 37642 30920 37648 30932
rect 36136 30892 37648 30920
rect 36136 30880 36142 30892
rect 37642 30880 37648 30892
rect 37700 30880 37706 30932
rect 16482 30852 16488 30864
rect 8536 30824 12112 30852
rect 16443 30824 16488 30852
rect 8536 30812 8542 30824
rect 16482 30812 16488 30824
rect 16540 30812 16546 30864
rect 19058 30852 19064 30864
rect 17880 30824 19064 30852
rect 7009 30787 7067 30793
rect 7009 30753 7021 30787
rect 7055 30753 7067 30787
rect 12342 30784 12348 30796
rect 12303 30756 12348 30784
rect 7009 30747 7067 30753
rect 12342 30744 12348 30756
rect 12400 30744 12406 30796
rect 12529 30787 12587 30793
rect 12529 30753 12541 30787
rect 12575 30784 12587 30787
rect 15841 30787 15899 30793
rect 15841 30784 15853 30787
rect 12575 30756 15853 30784
rect 12575 30753 12587 30756
rect 12529 30747 12587 30753
rect 15841 30753 15853 30756
rect 15887 30784 15899 30787
rect 16114 30784 16120 30796
rect 15887 30756 16120 30784
rect 15887 30753 15899 30756
rect 15841 30747 15899 30753
rect 16114 30744 16120 30756
rect 16172 30744 16178 30796
rect 7282 30725 7288 30728
rect 7276 30716 7288 30725
rect 7243 30688 7288 30716
rect 7276 30679 7288 30688
rect 7282 30676 7288 30679
rect 7340 30676 7346 30728
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30716 12311 30719
rect 12986 30716 12992 30728
rect 12299 30688 12992 30716
rect 12299 30685 12311 30688
rect 12253 30679 12311 30685
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 17880 30716 17908 30824
rect 19058 30812 19064 30824
rect 19116 30812 19122 30864
rect 17954 30744 17960 30796
rect 18012 30784 18018 30796
rect 21453 30787 21511 30793
rect 21453 30784 21465 30787
rect 18012 30756 21465 30784
rect 18012 30744 18018 30756
rect 21453 30753 21465 30756
rect 21499 30753 21511 30787
rect 21453 30747 21511 30753
rect 13096 30688 17908 30716
rect 1854 30648 1860 30660
rect 1815 30620 1860 30648
rect 1854 30608 1860 30620
rect 1912 30648 1918 30660
rect 2501 30651 2559 30657
rect 2501 30648 2513 30651
rect 1912 30620 2513 30648
rect 1912 30608 1918 30620
rect 2501 30617 2513 30620
rect 2547 30617 2559 30651
rect 2501 30611 2559 30617
rect 1946 30580 1952 30592
rect 1907 30552 1952 30580
rect 1946 30540 1952 30552
rect 2004 30540 2010 30592
rect 7742 30540 7748 30592
rect 7800 30580 7806 30592
rect 8389 30583 8447 30589
rect 8389 30580 8401 30583
rect 7800 30552 8401 30580
rect 7800 30540 7806 30552
rect 8389 30549 8401 30552
rect 8435 30580 8447 30583
rect 13096 30580 13124 30688
rect 16117 30651 16175 30657
rect 16117 30617 16129 30651
rect 16163 30648 16175 30651
rect 17972 30648 18000 30744
rect 21637 30719 21695 30725
rect 21637 30716 21649 30719
rect 16163 30620 18000 30648
rect 21008 30688 21649 30716
rect 16163 30617 16175 30620
rect 16117 30611 16175 30617
rect 21008 30592 21036 30688
rect 21637 30685 21649 30688
rect 21683 30685 21695 30719
rect 21637 30679 21695 30685
rect 35342 30676 35348 30728
rect 35400 30716 35406 30728
rect 35621 30719 35679 30725
rect 35621 30716 35633 30719
rect 35400 30688 35633 30716
rect 35400 30676 35406 30688
rect 35621 30685 35633 30688
rect 35667 30716 35679 30719
rect 35802 30716 35808 30728
rect 35667 30688 35808 30716
rect 35667 30685 35679 30688
rect 35621 30679 35679 30685
rect 35802 30676 35808 30688
rect 35860 30716 35866 30728
rect 36265 30719 36323 30725
rect 36265 30716 36277 30719
rect 35860 30688 36277 30716
rect 35860 30676 35866 30688
rect 36265 30685 36277 30688
rect 36311 30685 36323 30719
rect 37366 30716 37372 30728
rect 37327 30688 37372 30716
rect 36265 30679 36323 30685
rect 37366 30676 37372 30688
rect 37424 30676 37430 30728
rect 37826 30716 37832 30728
rect 37787 30688 37832 30716
rect 37826 30676 37832 30688
rect 37884 30676 37890 30728
rect 33873 30651 33931 30657
rect 33873 30617 33885 30651
rect 33919 30648 33931 30651
rect 36170 30648 36176 30660
rect 33919 30620 36176 30648
rect 33919 30617 33931 30620
rect 33873 30611 33931 30617
rect 36170 30608 36176 30620
rect 36228 30608 36234 30660
rect 16022 30580 16028 30592
rect 8435 30552 13124 30580
rect 15983 30552 16028 30580
rect 8435 30549 8447 30552
rect 8389 30543 8447 30549
rect 16022 30540 16028 30552
rect 16080 30540 16086 30592
rect 20990 30580 20996 30592
rect 20951 30552 20996 30580
rect 20990 30540 20996 30552
rect 21048 30540 21054 30592
rect 21818 30580 21824 30592
rect 21779 30552 21824 30580
rect 21818 30540 21824 30552
rect 21876 30540 21882 30592
rect 37182 30580 37188 30592
rect 37143 30552 37188 30580
rect 37182 30540 37188 30552
rect 37240 30540 37246 30592
rect 38010 30580 38016 30592
rect 37971 30552 38016 30580
rect 38010 30540 38016 30552
rect 38068 30540 38074 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 36170 30308 36176 30320
rect 36131 30280 36176 30308
rect 36170 30268 36176 30280
rect 36228 30268 36234 30320
rect 37642 30308 37648 30320
rect 36372 30280 37648 30308
rect 1949 30243 2007 30249
rect 1949 30209 1961 30243
rect 1995 30240 2007 30243
rect 16022 30240 16028 30252
rect 1995 30212 16028 30240
rect 1995 30209 2007 30212
rect 1949 30203 2007 30209
rect 16022 30200 16028 30212
rect 16080 30200 16086 30252
rect 21818 30200 21824 30252
rect 21876 30240 21882 30252
rect 23109 30243 23167 30249
rect 23109 30240 23121 30243
rect 21876 30212 23121 30240
rect 21876 30200 21882 30212
rect 23109 30209 23121 30212
rect 23155 30209 23167 30243
rect 23109 30203 23167 30209
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30240 23443 30243
rect 23431 30212 27108 30240
rect 23431 30209 23443 30212
rect 23385 30203 23443 30209
rect 2222 30172 2228 30184
rect 2183 30144 2228 30172
rect 2222 30132 2228 30144
rect 2280 30172 2286 30184
rect 2685 30175 2743 30181
rect 2685 30172 2697 30175
rect 2280 30144 2697 30172
rect 2280 30132 2286 30144
rect 2685 30141 2697 30144
rect 2731 30141 2743 30175
rect 26421 30175 26479 30181
rect 26421 30172 26433 30175
rect 2685 30135 2743 30141
rect 26206 30144 26433 30172
rect 1946 30064 1952 30116
rect 2004 30104 2010 30116
rect 26206 30104 26234 30144
rect 26421 30141 26433 30144
rect 26467 30172 26479 30175
rect 26973 30175 27031 30181
rect 26973 30172 26985 30175
rect 26467 30144 26985 30172
rect 26467 30141 26479 30144
rect 26421 30135 26479 30141
rect 26973 30141 26985 30144
rect 27019 30141 27031 30175
rect 27080 30172 27108 30212
rect 27154 30200 27160 30252
rect 27212 30240 27218 30252
rect 36372 30249 36400 30280
rect 37642 30268 37648 30280
rect 37700 30268 37706 30320
rect 27341 30243 27399 30249
rect 27212 30212 27257 30240
rect 27212 30200 27218 30212
rect 27341 30209 27353 30243
rect 27387 30240 27399 30243
rect 28077 30243 28135 30249
rect 28077 30240 28089 30243
rect 27387 30212 28089 30240
rect 27387 30209 27399 30212
rect 27341 30203 27399 30209
rect 28077 30209 28089 30212
rect 28123 30209 28135 30243
rect 28077 30203 28135 30209
rect 36357 30243 36415 30249
rect 36357 30209 36369 30243
rect 36403 30209 36415 30243
rect 36357 30203 36415 30209
rect 36541 30243 36599 30249
rect 36541 30209 36553 30243
rect 36587 30240 36599 30243
rect 37182 30240 37188 30252
rect 36587 30212 37188 30240
rect 36587 30209 36599 30212
rect 36541 30203 36599 30209
rect 37182 30200 37188 30212
rect 37240 30200 37246 30252
rect 37458 30200 37464 30252
rect 37516 30240 37522 30252
rect 37829 30243 37887 30249
rect 37829 30240 37841 30243
rect 37516 30212 37841 30240
rect 37516 30200 37522 30212
rect 37829 30209 37841 30212
rect 37875 30209 37887 30243
rect 37829 30203 37887 30209
rect 37274 30172 37280 30184
rect 27080 30144 37280 30172
rect 26973 30135 27031 30141
rect 37274 30132 37280 30144
rect 37332 30132 37338 30184
rect 2004 30076 26234 30104
rect 28261 30107 28319 30113
rect 2004 30064 2010 30076
rect 28261 30073 28273 30107
rect 28307 30104 28319 30107
rect 37826 30104 37832 30116
rect 28307 30076 37832 30104
rect 28307 30073 28319 30076
rect 28261 30067 28319 30073
rect 37826 30064 37832 30076
rect 37884 30064 37890 30116
rect 3326 30036 3332 30048
rect 3287 30008 3332 30036
rect 3326 29996 3332 30008
rect 3384 29996 3390 30048
rect 37366 30036 37372 30048
rect 37327 30008 37372 30036
rect 37366 29996 37372 30008
rect 37424 29996 37430 30048
rect 38013 30039 38071 30045
rect 38013 30005 38025 30039
rect 38059 30036 38071 30039
rect 38102 30036 38108 30048
rect 38059 30008 38108 30036
rect 38059 30005 38071 30008
rect 38013 29999 38071 30005
rect 38102 29996 38108 30008
rect 38160 29996 38166 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 3326 29792 3332 29844
rect 3384 29832 3390 29844
rect 35434 29832 35440 29844
rect 3384 29804 35440 29832
rect 3384 29792 3390 29804
rect 35434 29792 35440 29804
rect 35492 29792 35498 29844
rect 2041 29699 2099 29705
rect 2041 29665 2053 29699
rect 2087 29696 2099 29699
rect 2087 29668 6914 29696
rect 2087 29665 2099 29668
rect 2041 29659 2099 29665
rect 2777 29631 2835 29637
rect 2777 29597 2789 29631
rect 2823 29628 2835 29631
rect 3326 29628 3332 29640
rect 2823 29600 3332 29628
rect 2823 29597 2835 29600
rect 2777 29591 2835 29597
rect 3326 29588 3332 29600
rect 3384 29588 3390 29640
rect 6886 29628 6914 29668
rect 26326 29628 26332 29640
rect 6886 29600 26332 29628
rect 26326 29588 26332 29600
rect 26384 29588 26390 29640
rect 36725 29631 36783 29637
rect 36725 29597 36737 29631
rect 36771 29628 36783 29631
rect 37182 29628 37188 29640
rect 36771 29600 37188 29628
rect 36771 29597 36783 29600
rect 36725 29591 36783 29597
rect 37182 29588 37188 29600
rect 37240 29588 37246 29640
rect 37274 29588 37280 29640
rect 37332 29628 37338 29640
rect 37829 29631 37887 29637
rect 37829 29628 37841 29631
rect 37332 29600 37841 29628
rect 37332 29588 37338 29600
rect 37829 29597 37841 29600
rect 37875 29597 37887 29631
rect 37829 29591 37887 29597
rect 1854 29560 1860 29572
rect 1815 29532 1860 29560
rect 1854 29520 1860 29532
rect 1912 29520 1918 29572
rect 2593 29495 2651 29501
rect 2593 29461 2605 29495
rect 2639 29492 2651 29495
rect 2774 29492 2780 29504
rect 2639 29464 2780 29492
rect 2639 29461 2651 29464
rect 2593 29455 2651 29461
rect 2774 29452 2780 29464
rect 2832 29452 2838 29504
rect 37369 29495 37427 29501
rect 37369 29461 37381 29495
rect 37415 29492 37427 29495
rect 37550 29492 37556 29504
rect 37415 29464 37556 29492
rect 37415 29461 37427 29464
rect 37369 29455 37427 29461
rect 37550 29452 37556 29464
rect 37608 29452 37614 29504
rect 38010 29492 38016 29504
rect 37971 29464 38016 29492
rect 38010 29452 38016 29464
rect 38068 29452 38074 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 26326 29288 26332 29300
rect 26287 29260 26332 29288
rect 26326 29248 26332 29260
rect 26384 29248 26390 29300
rect 35434 29288 35440 29300
rect 35395 29260 35440 29288
rect 35434 29248 35440 29260
rect 35492 29248 35498 29300
rect 1854 29180 1860 29232
rect 1912 29220 1918 29232
rect 3237 29223 3295 29229
rect 3237 29220 3249 29223
rect 1912 29192 3249 29220
rect 1912 29180 1918 29192
rect 3237 29189 3249 29192
rect 3283 29189 3295 29223
rect 3237 29183 3295 29189
rect 1949 29155 2007 29161
rect 1949 29121 1961 29155
rect 1995 29152 2007 29155
rect 16298 29152 16304 29164
rect 1995 29124 16304 29152
rect 1995 29121 2007 29124
rect 1949 29115 2007 29121
rect 16298 29112 16304 29124
rect 16356 29112 16362 29164
rect 26344 29152 26372 29248
rect 37642 29220 37648 29232
rect 37476 29192 37648 29220
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26344 29124 26985 29152
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 27154 29152 27160 29164
rect 27115 29124 27160 29152
rect 26973 29115 27031 29121
rect 27154 29112 27160 29124
rect 27212 29112 27218 29164
rect 27341 29155 27399 29161
rect 27341 29121 27353 29155
rect 27387 29152 27399 29155
rect 27985 29155 28043 29161
rect 27985 29152 27997 29155
rect 27387 29124 27997 29152
rect 27387 29121 27399 29124
rect 27341 29115 27399 29121
rect 27985 29121 27997 29124
rect 28031 29121 28043 29155
rect 27985 29115 28043 29121
rect 35621 29155 35679 29161
rect 35621 29121 35633 29155
rect 35667 29152 35679 29155
rect 37277 29155 37335 29161
rect 37277 29152 37289 29155
rect 35667 29124 37289 29152
rect 35667 29121 35679 29124
rect 35621 29115 35679 29121
rect 37277 29121 37289 29124
rect 37323 29121 37335 29155
rect 37277 29115 37335 29121
rect 37366 29112 37372 29164
rect 37424 29152 37430 29164
rect 37476 29161 37504 29192
rect 37642 29180 37648 29192
rect 37700 29180 37706 29232
rect 37461 29155 37519 29161
rect 37461 29152 37473 29155
rect 37424 29124 37473 29152
rect 37424 29112 37430 29124
rect 37461 29121 37473 29124
rect 37507 29121 37519 29155
rect 37461 29115 37519 29121
rect 37550 29112 37556 29164
rect 37608 29152 37614 29164
rect 37608 29124 37653 29152
rect 37608 29112 37614 29124
rect 2222 29084 2228 29096
rect 2183 29056 2228 29084
rect 2222 29044 2228 29056
rect 2280 29084 2286 29096
rect 2685 29087 2743 29093
rect 2685 29084 2697 29087
rect 2280 29056 2697 29084
rect 2280 29044 2286 29056
rect 2685 29053 2697 29056
rect 2731 29053 2743 29087
rect 2685 29047 2743 29053
rect 28169 29019 28227 29025
rect 28169 28985 28181 29019
rect 28215 29016 28227 29019
rect 37458 29016 37464 29028
rect 28215 28988 37464 29016
rect 28215 28985 28227 28988
rect 28169 28979 28227 28985
rect 37458 28976 37464 28988
rect 37516 28976 37522 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 23247 28747 23305 28753
rect 23247 28713 23259 28747
rect 23293 28744 23305 28747
rect 23293 28716 26004 28744
rect 23293 28713 23305 28716
rect 23247 28707 23305 28713
rect 16761 28679 16819 28685
rect 16761 28645 16773 28679
rect 16807 28645 16819 28679
rect 16761 28639 16819 28645
rect 16114 28608 16120 28620
rect 16075 28580 16120 28608
rect 16114 28568 16120 28580
rect 16172 28568 16178 28620
rect 16298 28608 16304 28620
rect 16259 28580 16304 28608
rect 16298 28568 16304 28580
rect 16356 28568 16362 28620
rect 1673 28543 1731 28549
rect 1673 28509 1685 28543
rect 1719 28509 1731 28543
rect 16776 28540 16804 28639
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 25869 28679 25927 28685
rect 25869 28676 25881 28679
rect 17276 28648 25881 28676
rect 17276 28636 17282 28648
rect 20990 28608 20996 28620
rect 20903 28580 20996 28608
rect 20990 28568 20996 28580
rect 21048 28608 21054 28620
rect 21048 28580 21588 28608
rect 21048 28568 21054 28580
rect 21560 28552 21588 28580
rect 17221 28543 17279 28549
rect 17221 28540 17233 28543
rect 16776 28512 17233 28540
rect 1673 28503 1731 28509
rect 17221 28509 17233 28512
rect 17267 28509 17279 28543
rect 21450 28540 21456 28552
rect 21411 28512 21456 28540
rect 17221 28503 17279 28509
rect 1688 28472 1716 28503
rect 21450 28500 21456 28512
rect 21508 28500 21514 28552
rect 21542 28500 21548 28552
rect 21600 28540 21606 28552
rect 21637 28543 21695 28549
rect 21637 28540 21649 28543
rect 21600 28512 21649 28540
rect 21600 28500 21606 28512
rect 21637 28509 21649 28512
rect 21683 28509 21695 28543
rect 21637 28503 21695 28509
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 23017 28543 23075 28549
rect 23017 28540 23029 28543
rect 21867 28512 23029 28540
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 23017 28509 23029 28512
rect 23063 28509 23075 28543
rect 25792 28540 25820 28648
rect 25869 28645 25881 28648
rect 25915 28645 25927 28679
rect 25869 28639 25927 28645
rect 25976 28608 26004 28716
rect 25976 28580 37872 28608
rect 26421 28543 26479 28549
rect 26421 28540 26433 28543
rect 25792 28512 26433 28540
rect 23017 28503 23075 28509
rect 26421 28509 26433 28512
rect 26467 28509 26479 28543
rect 26421 28503 26479 28509
rect 26605 28543 26663 28549
rect 26605 28509 26617 28543
rect 26651 28540 26663 28543
rect 27154 28540 27160 28552
rect 26651 28512 27160 28540
rect 26651 28509 26663 28512
rect 26605 28503 26663 28509
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 36725 28543 36783 28549
rect 36725 28509 36737 28543
rect 36771 28540 36783 28543
rect 37182 28540 37188 28552
rect 36771 28512 37188 28540
rect 36771 28509 36783 28512
rect 36725 28503 36783 28509
rect 37182 28500 37188 28512
rect 37240 28500 37246 28552
rect 37844 28549 37872 28580
rect 37829 28543 37887 28549
rect 37829 28509 37841 28543
rect 37875 28509 37887 28543
rect 37829 28503 37887 28509
rect 2777 28475 2835 28481
rect 2777 28472 2789 28475
rect 1688 28444 2789 28472
rect 2777 28441 2789 28444
rect 2823 28472 2835 28475
rect 35802 28472 35808 28484
rect 2823 28444 35808 28472
rect 2823 28441 2835 28444
rect 2777 28435 2835 28441
rect 35802 28432 35808 28444
rect 35860 28432 35866 28484
rect 1486 28404 1492 28416
rect 1447 28376 1492 28404
rect 1486 28364 1492 28376
rect 1544 28364 1550 28416
rect 1854 28364 1860 28416
rect 1912 28404 1918 28416
rect 2133 28407 2191 28413
rect 2133 28404 2145 28407
rect 1912 28376 2145 28404
rect 1912 28364 1918 28376
rect 2133 28373 2145 28376
rect 2179 28373 2191 28407
rect 2133 28367 2191 28373
rect 16393 28407 16451 28413
rect 16393 28373 16405 28407
rect 16439 28404 16451 28407
rect 17310 28404 17316 28416
rect 16439 28376 17316 28404
rect 16439 28373 16451 28376
rect 16393 28367 16451 28373
rect 17310 28364 17316 28376
rect 17368 28364 17374 28416
rect 17405 28407 17463 28413
rect 17405 28373 17417 28407
rect 17451 28404 17463 28407
rect 18230 28404 18236 28416
rect 17451 28376 18236 28404
rect 17451 28373 17463 28376
rect 17405 28367 17463 28373
rect 18230 28364 18236 28376
rect 18288 28364 18294 28416
rect 26789 28407 26847 28413
rect 26789 28373 26801 28407
rect 26835 28404 26847 28407
rect 27890 28404 27896 28416
rect 26835 28376 27896 28404
rect 26835 28373 26847 28376
rect 26789 28367 26847 28373
rect 27890 28364 27896 28376
rect 27948 28364 27954 28416
rect 37369 28407 37427 28413
rect 37369 28373 37381 28407
rect 37415 28404 37427 28407
rect 37550 28404 37556 28416
rect 37415 28376 37556 28404
rect 37415 28373 37427 28376
rect 37369 28367 37427 28373
rect 37550 28364 37556 28376
rect 37608 28364 37614 28416
rect 38010 28404 38016 28416
rect 37971 28376 38016 28404
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 17402 28200 17408 28212
rect 17363 28172 17408 28200
rect 17402 28160 17408 28172
rect 17460 28160 17466 28212
rect 35802 28200 35808 28212
rect 35763 28172 35808 28200
rect 35802 28160 35808 28172
rect 35860 28160 35866 28212
rect 2041 28135 2099 28141
rect 2041 28101 2053 28135
rect 2087 28132 2099 28135
rect 17218 28132 17224 28144
rect 2087 28104 17224 28132
rect 2087 28101 2099 28104
rect 2041 28095 2099 28101
rect 17218 28092 17224 28104
rect 17276 28092 17282 28144
rect 1854 28064 1860 28076
rect 1815 28036 1860 28064
rect 1854 28024 1860 28036
rect 1912 28024 1918 28076
rect 2501 28067 2559 28073
rect 2501 28033 2513 28067
rect 2547 28064 2559 28067
rect 2774 28064 2780 28076
rect 2547 28036 2780 28064
rect 2547 28033 2559 28036
rect 2501 28027 2559 28033
rect 2774 28024 2780 28036
rect 2832 28064 2838 28076
rect 3145 28067 3203 28073
rect 3145 28064 3157 28067
rect 2832 28036 3157 28064
rect 2832 28024 2838 28036
rect 3145 28033 3157 28036
rect 3191 28033 3203 28067
rect 17420 28064 17448 28160
rect 18230 28141 18236 28144
rect 18224 28132 18236 28141
rect 18191 28104 18236 28132
rect 18224 28095 18236 28104
rect 18230 28092 18236 28095
rect 18288 28092 18294 28144
rect 17957 28067 18015 28073
rect 17957 28064 17969 28067
rect 17420 28036 17969 28064
rect 3145 28027 3203 28033
rect 17957 28033 17969 28036
rect 18003 28033 18015 28067
rect 27890 28064 27896 28076
rect 27851 28036 27896 28064
rect 17957 28027 18015 28033
rect 27890 28024 27896 28036
rect 27948 28024 27954 28076
rect 35989 28067 36047 28073
rect 35989 28033 36001 28067
rect 36035 28064 36047 28067
rect 37277 28067 37335 28073
rect 37277 28064 37289 28067
rect 36035 28036 37289 28064
rect 36035 28033 36047 28036
rect 35989 28027 36047 28033
rect 37277 28033 37289 28036
rect 37323 28033 37335 28067
rect 37277 28027 37335 28033
rect 37366 28024 37372 28076
rect 37424 28064 37430 28076
rect 37461 28067 37519 28073
rect 37461 28064 37473 28067
rect 37424 28036 37473 28064
rect 37424 28024 37430 28036
rect 37461 28033 37473 28036
rect 37507 28033 37519 28067
rect 37461 28027 37519 28033
rect 37550 28024 37556 28076
rect 37608 28064 37614 28076
rect 37608 28036 37653 28064
rect 37608 28024 37614 28036
rect 28077 27931 28135 27937
rect 28077 27897 28089 27931
rect 28123 27928 28135 27931
rect 37090 27928 37096 27940
rect 28123 27900 37096 27928
rect 28123 27897 28135 27900
rect 28077 27891 28135 27897
rect 37090 27888 37096 27900
rect 37148 27888 37154 27940
rect 2682 27860 2688 27872
rect 2643 27832 2688 27860
rect 2682 27820 2688 27832
rect 2740 27820 2746 27872
rect 17310 27820 17316 27872
rect 17368 27860 17374 27872
rect 19337 27863 19395 27869
rect 19337 27860 19349 27863
rect 17368 27832 19349 27860
rect 17368 27820 17374 27832
rect 19337 27829 19349 27832
rect 19383 27860 19395 27863
rect 21450 27860 21456 27872
rect 19383 27832 21456 27860
rect 19383 27829 19395 27832
rect 19337 27823 19395 27829
rect 21450 27820 21456 27832
rect 21508 27820 21514 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2682 27616 2688 27668
rect 2740 27656 2746 27668
rect 12250 27656 12256 27668
rect 2740 27628 12256 27656
rect 2740 27616 2746 27628
rect 12250 27616 12256 27628
rect 12308 27616 12314 27668
rect 9030 27588 9036 27600
rect 8991 27560 9036 27588
rect 9030 27548 9036 27560
rect 9088 27548 9094 27600
rect 37274 27588 37280 27600
rect 37235 27560 37280 27588
rect 37274 27548 37280 27560
rect 37332 27548 37338 27600
rect 1673 27455 1731 27461
rect 1673 27421 1685 27455
rect 1719 27452 1731 27455
rect 7009 27455 7067 27461
rect 1719 27424 2820 27452
rect 1719 27421 1731 27424
rect 1673 27415 1731 27421
rect 1486 27316 1492 27328
rect 1447 27288 1492 27316
rect 1486 27276 1492 27288
rect 1544 27276 1550 27328
rect 1946 27276 1952 27328
rect 2004 27316 2010 27328
rect 2792 27325 2820 27424
rect 7009 27421 7021 27455
rect 7055 27452 7067 27455
rect 8294 27452 8300 27464
rect 7055 27424 8300 27452
rect 7055 27421 7067 27424
rect 7009 27415 7067 27421
rect 8294 27412 8300 27424
rect 8352 27452 8358 27464
rect 9048 27452 9076 27548
rect 8352 27424 9076 27452
rect 11885 27455 11943 27461
rect 8352 27412 8358 27424
rect 11885 27421 11897 27455
rect 11931 27452 11943 27455
rect 11974 27452 11980 27464
rect 11931 27424 11980 27452
rect 11931 27421 11943 27424
rect 11885 27415 11943 27421
rect 11974 27412 11980 27424
rect 12032 27412 12038 27464
rect 37090 27452 37096 27464
rect 37051 27424 37096 27452
rect 37090 27412 37096 27424
rect 37148 27412 37154 27464
rect 37826 27452 37832 27464
rect 37787 27424 37832 27452
rect 37826 27412 37832 27424
rect 37884 27412 37890 27464
rect 7098 27344 7104 27396
rect 7156 27384 7162 27396
rect 7254 27387 7312 27393
rect 7254 27384 7266 27387
rect 7156 27356 7266 27384
rect 7156 27344 7162 27356
rect 7254 27353 7266 27356
rect 7300 27353 7312 27387
rect 34790 27384 34796 27396
rect 7254 27347 7312 27353
rect 8220 27356 34796 27384
rect 2133 27319 2191 27325
rect 2133 27316 2145 27319
rect 2004 27288 2145 27316
rect 2004 27276 2010 27288
rect 2133 27285 2145 27288
rect 2179 27285 2191 27319
rect 2133 27279 2191 27285
rect 2777 27319 2835 27325
rect 2777 27285 2789 27319
rect 2823 27316 2835 27319
rect 8220 27316 8248 27356
rect 34790 27344 34796 27356
rect 34848 27344 34854 27396
rect 8386 27316 8392 27328
rect 2823 27288 8248 27316
rect 8347 27288 8392 27316
rect 2823 27285 2835 27288
rect 2777 27279 2835 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 12066 27316 12072 27328
rect 12027 27288 12072 27316
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 38010 27316 38016 27328
rect 37971 27288 38016 27316
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 12066 27053 12072 27056
rect 12060 27044 12072 27053
rect 12027 27016 12072 27044
rect 12060 27007 12072 27016
rect 12066 27004 12072 27007
rect 12124 27004 12130 27056
rect 1949 26979 2007 26985
rect 1949 26945 1961 26979
rect 1995 26976 2007 26979
rect 16482 26976 16488 26988
rect 1995 26948 16488 26976
rect 1995 26945 2007 26948
rect 1949 26939 2007 26945
rect 16482 26936 16488 26948
rect 16540 26936 16546 26988
rect 23842 26936 23848 26988
rect 23900 26976 23906 26988
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 23900 26948 25605 26976
rect 23900 26936 23906 26948
rect 25593 26945 25605 26948
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 31294 26936 31300 26988
rect 31352 26976 31358 26988
rect 37829 26979 37887 26985
rect 37829 26976 37841 26979
rect 31352 26948 37841 26976
rect 31352 26936 31358 26948
rect 37829 26945 37841 26948
rect 37875 26945 37887 26979
rect 37829 26939 37887 26945
rect 2222 26908 2228 26920
rect 2183 26880 2228 26908
rect 2222 26868 2228 26880
rect 2280 26908 2286 26920
rect 2685 26911 2743 26917
rect 2685 26908 2697 26911
rect 2280 26880 2697 26908
rect 2280 26868 2286 26880
rect 2685 26877 2697 26880
rect 2731 26877 2743 26911
rect 10962 26908 10968 26920
rect 10875 26880 10968 26908
rect 2685 26871 2743 26877
rect 10962 26868 10968 26880
rect 11020 26908 11026 26920
rect 11793 26911 11851 26917
rect 11793 26908 11805 26911
rect 11020 26880 11805 26908
rect 11020 26868 11026 26880
rect 11793 26877 11805 26880
rect 11839 26877 11851 26911
rect 11793 26871 11851 26877
rect 1854 26732 1860 26784
rect 1912 26772 1918 26784
rect 3237 26775 3295 26781
rect 3237 26772 3249 26775
rect 1912 26744 3249 26772
rect 1912 26732 1918 26744
rect 3237 26741 3249 26744
rect 3283 26741 3295 26775
rect 13170 26772 13176 26784
rect 13083 26744 13176 26772
rect 3237 26735 3295 26741
rect 13170 26732 13176 26744
rect 13228 26772 13234 26784
rect 23474 26772 23480 26784
rect 13228 26744 23480 26772
rect 13228 26732 13234 26744
rect 23474 26732 23480 26744
rect 23532 26732 23538 26784
rect 25777 26775 25835 26781
rect 25777 26741 25789 26775
rect 25823 26772 25835 26775
rect 37826 26772 37832 26784
rect 25823 26744 37832 26772
rect 25823 26741 25835 26744
rect 25777 26735 25835 26741
rect 37826 26732 37832 26744
rect 37884 26732 37890 26784
rect 38010 26772 38016 26784
rect 37971 26744 38016 26772
rect 38010 26732 38016 26744
rect 38068 26732 38074 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 7098 26568 7104 26580
rect 7059 26540 7104 26568
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 11974 26568 11980 26580
rect 11935 26540 11980 26568
rect 11974 26528 11980 26540
rect 12032 26528 12038 26580
rect 28997 26571 29055 26577
rect 28997 26568 29009 26571
rect 16546 26540 29009 26568
rect 2593 26503 2651 26509
rect 2593 26469 2605 26503
rect 2639 26500 2651 26503
rect 2774 26500 2780 26512
rect 2639 26472 2780 26500
rect 2639 26469 2651 26472
rect 2593 26463 2651 26469
rect 2774 26460 2780 26472
rect 2832 26460 2838 26512
rect 16546 26500 16574 26540
rect 28997 26537 29009 26540
rect 29043 26568 29055 26571
rect 31294 26568 31300 26580
rect 29043 26540 29592 26568
rect 31255 26540 31300 26568
rect 29043 26537 29055 26540
rect 28997 26531 29055 26537
rect 23842 26500 23848 26512
rect 6886 26472 16574 26500
rect 23803 26472 23848 26500
rect 2041 26435 2099 26441
rect 2041 26401 2053 26435
rect 2087 26432 2099 26435
rect 6886 26432 6914 26472
rect 23842 26460 23848 26472
rect 23900 26460 23906 26512
rect 2087 26404 6914 26432
rect 2087 26401 2099 26404
rect 2041 26395 2099 26401
rect 12250 26392 12256 26444
rect 12308 26432 12314 26444
rect 12437 26435 12495 26441
rect 12437 26432 12449 26435
rect 12308 26404 12449 26432
rect 12308 26392 12314 26404
rect 12437 26401 12449 26404
rect 12483 26401 12495 26435
rect 12437 26395 12495 26401
rect 12621 26435 12679 26441
rect 12621 26401 12633 26435
rect 12667 26432 12679 26435
rect 16114 26432 16120 26444
rect 12667 26404 16120 26432
rect 12667 26401 12679 26404
rect 12621 26395 12679 26401
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 23474 26432 23480 26444
rect 23435 26404 23480 26432
rect 23474 26392 23480 26404
rect 23532 26392 23538 26444
rect 29564 26441 29592 26540
rect 31294 26528 31300 26540
rect 31352 26528 31358 26580
rect 34790 26528 34796 26580
rect 34848 26568 34854 26580
rect 35069 26571 35127 26577
rect 35069 26568 35081 26571
rect 34848 26540 35081 26568
rect 34848 26528 34854 26540
rect 35069 26537 35081 26540
rect 35115 26537 35127 26571
rect 35069 26531 35127 26537
rect 29549 26435 29607 26441
rect 29549 26401 29561 26435
rect 29595 26401 29607 26435
rect 29549 26395 29607 26401
rect 1854 26364 1860 26376
rect 1815 26336 1860 26364
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 2777 26367 2835 26373
rect 2777 26333 2789 26367
rect 2823 26364 2835 26367
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 2823 26336 3801 26364
rect 2823 26333 2835 26336
rect 2777 26327 2835 26333
rect 3789 26333 3801 26336
rect 3835 26364 3847 26367
rect 3878 26364 3884 26376
rect 3835 26336 3884 26364
rect 3835 26333 3847 26336
rect 3789 26327 3847 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 6914 26324 6920 26376
rect 6972 26364 6978 26376
rect 12345 26367 12403 26373
rect 6972 26336 7017 26364
rect 6972 26324 6978 26336
rect 12345 26333 12357 26367
rect 12391 26364 12403 26367
rect 13170 26364 13176 26376
rect 12391 26336 13176 26364
rect 12391 26333 12403 26336
rect 12345 26327 12403 26333
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26333 23719 26367
rect 23661 26327 23719 26333
rect 23382 26256 23388 26308
rect 23440 26296 23446 26308
rect 23676 26296 23704 26327
rect 29638 26324 29644 26376
rect 29696 26364 29702 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 29696 26336 29745 26364
rect 29696 26324 29702 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26364 29975 26367
rect 31113 26367 31171 26373
rect 31113 26364 31125 26367
rect 29963 26336 31125 26364
rect 29963 26333 29975 26336
rect 29917 26327 29975 26333
rect 31113 26333 31125 26336
rect 31159 26333 31171 26367
rect 35250 26364 35256 26376
rect 35211 26336 35256 26364
rect 31113 26327 31171 26333
rect 35250 26324 35256 26336
rect 35308 26324 35314 26376
rect 37461 26367 37519 26373
rect 37461 26333 37473 26367
rect 37507 26364 37519 26367
rect 38102 26364 38108 26376
rect 37507 26336 38108 26364
rect 37507 26333 37519 26336
rect 37461 26327 37519 26333
rect 38102 26324 38108 26336
rect 38160 26324 38166 26376
rect 23440 26268 23704 26296
rect 23440 26256 23446 26268
rect 8294 26188 8300 26240
rect 8352 26228 8358 26240
rect 10962 26228 10968 26240
rect 8352 26200 10968 26228
rect 8352 26188 8358 26200
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 37734 26188 37740 26240
rect 37792 26228 37798 26240
rect 37921 26231 37979 26237
rect 37921 26228 37933 26231
rect 37792 26200 37933 26228
rect 37792 26188 37798 26200
rect 37921 26197 37933 26200
rect 37967 26197 37979 26231
rect 37921 26191 37979 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 16945 26027 17003 26033
rect 16945 26024 16957 26027
rect 16540 25996 16957 26024
rect 16540 25984 16546 25996
rect 16945 25993 16957 25996
rect 16991 25993 17003 26027
rect 16945 25987 17003 25993
rect 27157 26027 27215 26033
rect 27157 25993 27169 26027
rect 27203 26024 27215 26027
rect 27203 25996 35204 26024
rect 27203 25993 27215 25996
rect 27157 25987 27215 25993
rect 1857 25959 1915 25965
rect 1857 25925 1869 25959
rect 1903 25956 1915 25959
rect 1946 25956 1952 25968
rect 1903 25928 1952 25956
rect 1903 25925 1915 25928
rect 1857 25919 1915 25925
rect 1946 25916 1952 25928
rect 2004 25916 2010 25968
rect 2041 25959 2099 25965
rect 2041 25925 2053 25959
rect 2087 25956 2099 25959
rect 3786 25956 3792 25968
rect 2087 25928 3792 25956
rect 2087 25925 2099 25928
rect 2041 25919 2099 25925
rect 3786 25916 3792 25928
rect 3844 25916 3850 25968
rect 3878 25916 3884 25968
rect 3936 25956 3942 25968
rect 35176 25956 35204 25996
rect 35250 25984 35256 26036
rect 35308 26024 35314 26036
rect 36173 26027 36231 26033
rect 36173 26024 36185 26027
rect 35308 25996 36185 26024
rect 35308 25984 35314 25996
rect 36173 25993 36185 25996
rect 36219 25993 36231 26027
rect 36173 25987 36231 25993
rect 3936 25928 31708 25956
rect 35176 25928 35894 25956
rect 3936 25916 3942 25928
rect 2958 25897 2964 25900
rect 2952 25851 2964 25897
rect 3016 25888 3022 25900
rect 17037 25891 17095 25897
rect 3016 25860 3052 25888
rect 2958 25848 2964 25851
rect 3016 25848 3022 25860
rect 17037 25857 17049 25891
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 23109 25891 23167 25897
rect 23109 25857 23121 25891
rect 23155 25857 23167 25891
rect 23109 25851 23167 25857
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25888 23351 25891
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 23339 25860 26985 25888
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 29638 25888 29644 25900
rect 29551 25860 29644 25888
rect 26973 25851 27031 25857
rect 2685 25823 2743 25829
rect 2685 25789 2697 25823
rect 2731 25789 2743 25823
rect 2685 25783 2743 25789
rect 2700 25684 2728 25783
rect 15838 25780 15844 25832
rect 15896 25820 15902 25832
rect 16114 25820 16120 25832
rect 15896 25792 16120 25820
rect 15896 25780 15902 25792
rect 16114 25780 16120 25792
rect 16172 25820 16178 25832
rect 16761 25823 16819 25829
rect 16761 25820 16773 25823
rect 16172 25792 16773 25820
rect 16172 25780 16178 25792
rect 16761 25789 16773 25792
rect 16807 25789 16819 25823
rect 17052 25820 17080 25851
rect 19334 25820 19340 25832
rect 17052 25792 19340 25820
rect 16761 25783 16819 25789
rect 19334 25780 19340 25792
rect 19392 25820 19398 25832
rect 22925 25823 22983 25829
rect 22925 25820 22937 25823
rect 19392 25792 22937 25820
rect 19392 25780 19398 25792
rect 22925 25789 22937 25792
rect 22971 25789 22983 25823
rect 23124 25820 23152 25851
rect 29638 25848 29644 25860
rect 29696 25888 29702 25900
rect 30006 25888 30012 25900
rect 29696 25860 30012 25888
rect 29696 25848 29702 25860
rect 30006 25848 30012 25860
rect 30064 25848 30070 25900
rect 23382 25820 23388 25832
rect 23124 25792 23388 25820
rect 22925 25783 22983 25789
rect 23382 25780 23388 25792
rect 23440 25780 23446 25832
rect 28994 25780 29000 25832
rect 29052 25820 29058 25832
rect 29457 25823 29515 25829
rect 29457 25820 29469 25823
rect 29052 25792 29469 25820
rect 29052 25780 29058 25792
rect 29457 25789 29469 25792
rect 29503 25789 29515 25823
rect 29457 25783 29515 25789
rect 3620 25724 4660 25752
rect 3620 25684 3648 25724
rect 4062 25684 4068 25696
rect 2700 25656 3648 25684
rect 4023 25656 4068 25684
rect 4062 25644 4068 25656
rect 4120 25644 4126 25696
rect 4632 25693 4660 25724
rect 4617 25687 4675 25693
rect 4617 25653 4629 25687
rect 4663 25684 4675 25687
rect 8294 25684 8300 25696
rect 4663 25656 8300 25684
rect 4663 25653 4675 25656
rect 4617 25647 4675 25653
rect 8294 25644 8300 25656
rect 8352 25644 8358 25696
rect 17034 25644 17040 25696
rect 17092 25684 17098 25696
rect 17405 25687 17463 25693
rect 17405 25684 17417 25687
rect 17092 25656 17417 25684
rect 17092 25644 17098 25656
rect 17405 25653 17417 25656
rect 17451 25653 17463 25687
rect 28994 25684 29000 25696
rect 28955 25656 29000 25684
rect 17405 25647 17463 25653
rect 28994 25644 29000 25656
rect 29052 25644 29058 25696
rect 29825 25687 29883 25693
rect 29825 25653 29837 25687
rect 29871 25684 29883 25687
rect 31478 25684 31484 25696
rect 29871 25656 31484 25684
rect 29871 25653 29883 25656
rect 29825 25647 29883 25653
rect 31478 25644 31484 25656
rect 31536 25644 31542 25696
rect 31680 25684 31708 25928
rect 35434 25888 35440 25900
rect 35395 25860 35440 25888
rect 35434 25848 35440 25860
rect 35492 25848 35498 25900
rect 35866 25752 35894 25928
rect 36357 25891 36415 25897
rect 36357 25857 36369 25891
rect 36403 25888 36415 25891
rect 36446 25888 36452 25900
rect 36403 25860 36452 25888
rect 36403 25857 36415 25860
rect 36357 25851 36415 25857
rect 36446 25848 36452 25860
rect 36504 25848 36510 25900
rect 36541 25891 36599 25897
rect 36541 25857 36553 25891
rect 36587 25888 36599 25891
rect 37734 25888 37740 25900
rect 36587 25860 37740 25888
rect 36587 25857 36599 25860
rect 36541 25851 36599 25857
rect 37734 25848 37740 25860
rect 37792 25848 37798 25900
rect 37829 25891 37887 25897
rect 37829 25857 37841 25891
rect 37875 25857 37887 25891
rect 37829 25851 37887 25857
rect 37844 25752 37872 25851
rect 38010 25752 38016 25764
rect 35866 25724 37872 25752
rect 37971 25724 38016 25752
rect 38010 25712 38016 25724
rect 38068 25712 38074 25764
rect 35253 25687 35311 25693
rect 35253 25684 35265 25687
rect 31680 25656 35265 25684
rect 35253 25653 35265 25656
rect 35299 25653 35311 25687
rect 35253 25647 35311 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2869 25483 2927 25489
rect 2869 25449 2881 25483
rect 2915 25480 2927 25483
rect 2958 25480 2964 25492
rect 2915 25452 2964 25480
rect 2915 25449 2927 25452
rect 2869 25443 2927 25449
rect 2958 25440 2964 25452
rect 3016 25440 3022 25492
rect 3786 25440 3792 25492
rect 3844 25480 3850 25492
rect 6733 25483 6791 25489
rect 3844 25452 4476 25480
rect 3844 25440 3850 25452
rect 2317 25415 2375 25421
rect 2317 25381 2329 25415
rect 2363 25412 2375 25415
rect 4448 25412 4476 25452
rect 6733 25449 6745 25483
rect 6779 25480 6791 25483
rect 6914 25480 6920 25492
rect 6779 25452 6920 25480
rect 6779 25449 6791 25452
rect 6733 25443 6791 25449
rect 6914 25440 6920 25452
rect 6972 25440 6978 25492
rect 28994 25480 29000 25492
rect 16546 25452 29000 25480
rect 16546 25412 16574 25452
rect 28994 25440 29000 25452
rect 29052 25440 29058 25492
rect 35434 25440 35440 25492
rect 35492 25480 35498 25492
rect 36357 25483 36415 25489
rect 36357 25480 36369 25483
rect 35492 25452 36369 25480
rect 35492 25440 35498 25452
rect 36357 25449 36369 25452
rect 36403 25449 36415 25483
rect 36357 25443 36415 25449
rect 37185 25415 37243 25421
rect 37185 25412 37197 25415
rect 2363 25384 4292 25412
rect 4448 25384 16574 25412
rect 36740 25384 37197 25412
rect 2363 25381 2375 25384
rect 2317 25375 2375 25381
rect 4264 25353 4292 25384
rect 4249 25347 4307 25353
rect 4249 25313 4261 25347
rect 4295 25313 4307 25347
rect 4249 25307 4307 25313
rect 4433 25347 4491 25353
rect 4433 25313 4445 25347
rect 4479 25344 4491 25347
rect 7285 25347 7343 25353
rect 7285 25344 7297 25347
rect 4479 25316 7297 25344
rect 4479 25313 4491 25316
rect 4433 25307 4491 25313
rect 7285 25313 7297 25316
rect 7331 25344 7343 25347
rect 7374 25344 7380 25356
rect 7331 25316 7380 25344
rect 7331 25313 7343 25316
rect 7285 25307 7343 25313
rect 7374 25304 7380 25316
rect 7432 25304 7438 25356
rect 36740 25353 36768 25384
rect 37185 25381 37197 25384
rect 37231 25381 37243 25415
rect 38010 25412 38016 25424
rect 37971 25384 38016 25412
rect 37185 25375 37243 25381
rect 38010 25372 38016 25384
rect 38068 25372 38074 25424
rect 36725 25347 36783 25353
rect 36725 25313 36737 25347
rect 36771 25313 36783 25347
rect 36725 25307 36783 25313
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25245 1731 25279
rect 2130 25276 2136 25288
rect 2091 25248 2136 25276
rect 1673 25239 1731 25245
rect 1688 25208 1716 25239
rect 2130 25236 2136 25248
rect 2188 25236 2194 25288
rect 3053 25279 3111 25285
rect 3053 25245 3065 25279
rect 3099 25276 3111 25279
rect 7101 25279 7159 25285
rect 3099 25248 3832 25276
rect 3099 25245 3111 25248
rect 3053 25239 3111 25245
rect 2682 25208 2688 25220
rect 1688 25180 2688 25208
rect 2682 25168 2688 25180
rect 2740 25168 2746 25220
rect 1486 25140 1492 25152
rect 1447 25112 1492 25140
rect 1486 25100 1492 25112
rect 1544 25100 1550 25152
rect 3804 25149 3832 25248
rect 7101 25245 7113 25279
rect 7147 25276 7159 25279
rect 17034 25276 17040 25288
rect 7147 25248 8064 25276
rect 16995 25248 17040 25276
rect 7147 25245 7159 25248
rect 7101 25239 7159 25245
rect 8036 25217 8064 25248
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25245 23259 25279
rect 23382 25276 23388 25288
rect 23343 25248 23388 25276
rect 23201 25239 23259 25245
rect 7193 25211 7251 25217
rect 7193 25208 7205 25211
rect 6886 25180 7205 25208
rect 3789 25143 3847 25149
rect 3789 25109 3801 25143
rect 3835 25109 3847 25143
rect 3789 25103 3847 25109
rect 4062 25100 4068 25152
rect 4120 25140 4126 25152
rect 4157 25143 4215 25149
rect 4157 25140 4169 25143
rect 4120 25112 4169 25140
rect 4120 25100 4126 25112
rect 4157 25109 4169 25112
rect 4203 25140 4215 25143
rect 5077 25143 5135 25149
rect 5077 25140 5089 25143
rect 4203 25112 5089 25140
rect 4203 25109 4215 25112
rect 4157 25103 4215 25109
rect 5077 25109 5089 25112
rect 5123 25140 5135 25143
rect 5534 25140 5540 25152
rect 5123 25112 5540 25140
rect 5123 25109 5135 25112
rect 5077 25103 5135 25109
rect 5534 25100 5540 25112
rect 5592 25100 5598 25152
rect 5626 25100 5632 25152
rect 5684 25140 5690 25152
rect 6886 25140 6914 25180
rect 7193 25177 7205 25180
rect 7239 25177 7251 25211
rect 7193 25171 7251 25177
rect 8021 25211 8079 25217
rect 8021 25177 8033 25211
rect 8067 25208 8079 25211
rect 8386 25208 8392 25220
rect 8067 25180 8392 25208
rect 8067 25177 8079 25180
rect 8021 25171 8079 25177
rect 8386 25168 8392 25180
rect 8444 25208 8450 25220
rect 22649 25211 22707 25217
rect 22649 25208 22661 25211
rect 8444 25180 22661 25208
rect 8444 25168 8450 25180
rect 22649 25177 22661 25180
rect 22695 25208 22707 25211
rect 23216 25208 23244 25239
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 24854 25236 24860 25288
rect 24912 25276 24918 25288
rect 26329 25279 26387 25285
rect 26329 25276 26341 25279
rect 24912 25248 26341 25276
rect 24912 25236 24918 25248
rect 26329 25245 26341 25248
rect 26375 25245 26387 25279
rect 28718 25276 28724 25288
rect 26329 25239 26387 25245
rect 28184 25248 28724 25276
rect 22695 25180 23244 25208
rect 22695 25177 22707 25180
rect 22649 25171 22707 25177
rect 17218 25140 17224 25152
rect 5684 25112 6914 25140
rect 17179 25112 17224 25140
rect 5684 25100 5690 25112
rect 17218 25100 17224 25112
rect 17276 25100 17282 25152
rect 23569 25143 23627 25149
rect 23569 25109 23581 25143
rect 23615 25140 23627 25143
rect 26234 25140 26240 25152
rect 23615 25112 26240 25140
rect 23615 25109 23627 25112
rect 23569 25103 23627 25109
rect 26234 25100 26240 25112
rect 26292 25100 26298 25152
rect 26510 25140 26516 25152
rect 26471 25112 26516 25140
rect 26510 25100 26516 25112
rect 26568 25100 26574 25152
rect 27614 25100 27620 25152
rect 27672 25140 27678 25152
rect 28184 25149 28212 25248
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 31478 25276 31484 25288
rect 31439 25248 31484 25276
rect 31478 25236 31484 25248
rect 31536 25236 31542 25288
rect 36538 25276 36544 25288
rect 36499 25248 36544 25276
rect 36538 25236 36544 25248
rect 36596 25236 36602 25288
rect 37366 25276 37372 25288
rect 37327 25248 37372 25276
rect 37366 25236 37372 25248
rect 37424 25236 37430 25288
rect 37829 25279 37887 25285
rect 37829 25245 37841 25279
rect 37875 25245 37887 25279
rect 37829 25239 37887 25245
rect 37844 25208 37872 25239
rect 35866 25180 37872 25208
rect 28169 25143 28227 25149
rect 28169 25140 28181 25143
rect 27672 25112 28181 25140
rect 27672 25100 27678 25112
rect 28169 25109 28181 25112
rect 28215 25109 28227 25143
rect 28169 25103 28227 25109
rect 28905 25143 28963 25149
rect 28905 25109 28917 25143
rect 28951 25140 28963 25143
rect 30006 25140 30012 25152
rect 28951 25112 30012 25140
rect 28951 25109 28963 25112
rect 28905 25103 28963 25109
rect 30006 25100 30012 25112
rect 30064 25100 30070 25152
rect 31665 25143 31723 25149
rect 31665 25109 31677 25143
rect 31711 25140 31723 25143
rect 35866 25140 35894 25180
rect 31711 25112 35894 25140
rect 31711 25109 31723 25112
rect 31665 25103 31723 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 2130 24896 2136 24948
rect 2188 24936 2194 24948
rect 2501 24939 2559 24945
rect 2501 24936 2513 24939
rect 2188 24908 2513 24936
rect 2188 24896 2194 24908
rect 2501 24905 2513 24908
rect 2547 24905 2559 24939
rect 19334 24936 19340 24948
rect 19295 24908 19340 24936
rect 2501 24899 2559 24905
rect 19334 24896 19340 24908
rect 19392 24896 19398 24948
rect 37366 24936 37372 24948
rect 37327 24908 37372 24936
rect 37366 24896 37372 24908
rect 37424 24896 37430 24948
rect 26510 24828 26516 24880
rect 26568 24868 26574 24880
rect 26568 24840 35894 24868
rect 26568 24828 26574 24840
rect 1854 24800 1860 24812
rect 1815 24772 1860 24800
rect 1854 24760 1860 24772
rect 1912 24800 1918 24812
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 1912 24772 3065 24800
rect 1912 24760 1918 24772
rect 3053 24769 3065 24772
rect 3099 24769 3111 24803
rect 3053 24763 3111 24769
rect 7929 24803 7987 24809
rect 7929 24769 7941 24803
rect 7975 24800 7987 24803
rect 8018 24800 8024 24812
rect 7975 24772 8024 24800
rect 7975 24769 7987 24772
rect 7929 24763 7987 24769
rect 8018 24760 8024 24772
rect 8076 24800 8082 24812
rect 8389 24803 8447 24809
rect 8389 24800 8401 24803
rect 8076 24772 8401 24800
rect 8076 24760 8082 24772
rect 8389 24769 8401 24772
rect 8435 24769 8447 24803
rect 8389 24763 8447 24769
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24800 14979 24803
rect 15378 24800 15384 24812
rect 14967 24772 15384 24800
rect 14967 24769 14979 24772
rect 14921 24763 14979 24769
rect 15378 24760 15384 24772
rect 15436 24760 15442 24812
rect 17218 24760 17224 24812
rect 17276 24800 17282 24812
rect 18213 24803 18271 24809
rect 18213 24800 18225 24803
rect 17276 24772 18225 24800
rect 17276 24760 17282 24772
rect 18213 24769 18225 24772
rect 18259 24769 18271 24803
rect 23382 24800 23388 24812
rect 23343 24772 23388 24800
rect 18213 24763 18271 24769
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 23569 24803 23627 24809
rect 23569 24769 23581 24803
rect 23615 24800 23627 24803
rect 24854 24800 24860 24812
rect 23615 24772 24860 24800
rect 23615 24769 23627 24772
rect 23569 24763 23627 24769
rect 24854 24760 24860 24772
rect 24912 24760 24918 24812
rect 35866 24800 35894 24840
rect 37829 24803 37887 24809
rect 37829 24800 37841 24803
rect 35866 24772 37841 24800
rect 37829 24769 37841 24772
rect 37875 24769 37887 24803
rect 37829 24763 37887 24769
rect 17402 24732 17408 24744
rect 17315 24704 17408 24732
rect 17402 24692 17408 24704
rect 17460 24732 17466 24744
rect 17957 24735 18015 24741
rect 17957 24732 17969 24735
rect 17460 24704 17969 24732
rect 17460 24692 17466 24704
rect 17957 24701 17969 24704
rect 18003 24701 18015 24735
rect 23201 24735 23259 24741
rect 23201 24732 23213 24735
rect 17957 24695 18015 24701
rect 22664 24704 23213 24732
rect 14737 24667 14795 24673
rect 14737 24633 14749 24667
rect 14783 24664 14795 24667
rect 15838 24664 15844 24676
rect 14783 24636 15844 24664
rect 14783 24633 14795 24636
rect 14737 24627 14795 24633
rect 15838 24624 15844 24636
rect 15896 24624 15902 24676
rect 1946 24596 1952 24608
rect 1907 24568 1952 24596
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 7374 24556 7380 24608
rect 7432 24596 7438 24608
rect 7745 24599 7803 24605
rect 7745 24596 7757 24599
rect 7432 24568 7757 24596
rect 7432 24556 7438 24568
rect 7745 24565 7757 24568
rect 7791 24565 7803 24599
rect 7745 24559 7803 24565
rect 17126 24556 17132 24608
rect 17184 24596 17190 24608
rect 17420 24605 17448 24692
rect 22664 24608 22692 24704
rect 23201 24701 23213 24704
rect 23247 24701 23259 24735
rect 23201 24695 23259 24701
rect 17405 24599 17463 24605
rect 17405 24596 17417 24599
rect 17184 24568 17417 24596
rect 17184 24556 17190 24568
rect 17405 24565 17417 24568
rect 17451 24565 17463 24599
rect 22646 24596 22652 24608
rect 22607 24568 22652 24596
rect 17405 24559 17463 24565
rect 22646 24556 22652 24568
rect 22704 24556 22710 24608
rect 38010 24596 38016 24608
rect 37971 24568 38016 24596
rect 38010 24556 38016 24568
rect 38068 24556 38074 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1946 24352 1952 24404
rect 2004 24392 2010 24404
rect 28997 24395 29055 24401
rect 28997 24392 29009 24395
rect 2004 24364 29009 24392
rect 2004 24352 2010 24364
rect 28997 24361 29009 24364
rect 29043 24392 29055 24395
rect 31757 24395 31815 24401
rect 29043 24364 29592 24392
rect 29043 24361 29055 24364
rect 28997 24355 29055 24361
rect 1581 24327 1639 24333
rect 1581 24293 1593 24327
rect 1627 24293 1639 24327
rect 1581 24287 1639 24293
rect 1596 24256 1624 24287
rect 5534 24284 5540 24336
rect 5592 24324 5598 24336
rect 22646 24324 22652 24336
rect 5592 24296 22652 24324
rect 5592 24284 5598 24296
rect 22646 24284 22652 24296
rect 22704 24284 22710 24336
rect 5626 24256 5632 24268
rect 1596 24228 5632 24256
rect 5626 24216 5632 24228
rect 5684 24216 5690 24268
rect 29564 24265 29592 24364
rect 31757 24361 31769 24395
rect 31803 24392 31815 24395
rect 31803 24364 37872 24392
rect 31803 24361 31815 24364
rect 31757 24355 31815 24361
rect 37185 24327 37243 24333
rect 37185 24324 37197 24327
rect 36740 24296 37197 24324
rect 29549 24259 29607 24265
rect 6886 24228 29500 24256
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24188 1458 24200
rect 2041 24191 2099 24197
rect 2041 24188 2053 24191
rect 1452 24160 2053 24188
rect 1452 24148 1458 24160
rect 2041 24157 2053 24160
rect 2087 24157 2099 24191
rect 2682 24188 2688 24200
rect 2595 24160 2688 24188
rect 2041 24151 2099 24157
rect 2682 24148 2688 24160
rect 2740 24188 2746 24200
rect 6886 24188 6914 24228
rect 2740 24160 6914 24188
rect 14369 24191 14427 24197
rect 2740 24148 2746 24160
rect 14369 24157 14381 24191
rect 14415 24188 14427 24191
rect 15378 24188 15384 24200
rect 14415 24160 15384 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 26292 24160 26337 24188
rect 26292 24148 26298 24160
rect 29472 24120 29500 24228
rect 29549 24225 29561 24259
rect 29595 24225 29607 24259
rect 30006 24256 30012 24268
rect 29549 24219 29607 24225
rect 29748 24228 30012 24256
rect 29748 24197 29776 24228
rect 30006 24216 30012 24228
rect 30064 24216 30070 24268
rect 36740 24265 36768 24296
rect 37185 24293 37197 24296
rect 37231 24293 37243 24327
rect 37185 24287 37243 24293
rect 36725 24259 36783 24265
rect 36725 24225 36737 24259
rect 36771 24225 36783 24259
rect 36725 24219 36783 24225
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24188 29975 24191
rect 31573 24191 31631 24197
rect 31573 24188 31585 24191
rect 29963 24160 31585 24188
rect 29963 24157 29975 24160
rect 29917 24151 29975 24157
rect 31573 24157 31585 24160
rect 31619 24157 31631 24191
rect 31573 24151 31631 24157
rect 34977 24191 35035 24197
rect 34977 24157 34989 24191
rect 35023 24157 35035 24191
rect 34977 24151 35035 24157
rect 34992 24120 35020 24151
rect 35342 24148 35348 24200
rect 35400 24188 35406 24200
rect 35529 24191 35587 24197
rect 35529 24188 35541 24191
rect 35400 24160 35541 24188
rect 35400 24148 35406 24160
rect 35529 24157 35541 24160
rect 35575 24157 35587 24191
rect 36538 24188 36544 24200
rect 36451 24160 36544 24188
rect 35529 24151 35587 24157
rect 36538 24148 36544 24160
rect 36596 24148 36602 24200
rect 37366 24188 37372 24200
rect 37327 24160 37372 24188
rect 37366 24148 37372 24160
rect 37424 24148 37430 24200
rect 37844 24197 37872 24364
rect 37829 24191 37887 24197
rect 37829 24157 37841 24191
rect 37875 24157 37887 24191
rect 37829 24151 37887 24157
rect 36357 24123 36415 24129
rect 36357 24120 36369 24123
rect 29472 24092 34836 24120
rect 34992 24092 36369 24120
rect 8018 24012 8024 24064
rect 8076 24052 8082 24064
rect 14185 24055 14243 24061
rect 14185 24052 14197 24055
rect 8076 24024 14197 24052
rect 8076 24012 8082 24024
rect 14185 24021 14197 24024
rect 14231 24021 14243 24055
rect 26418 24052 26424 24064
rect 26379 24024 26424 24052
rect 14185 24015 14243 24021
rect 26418 24012 26424 24024
rect 26476 24012 26482 24064
rect 34808 24061 34836 24092
rect 36357 24089 36369 24092
rect 36403 24089 36415 24123
rect 36357 24083 36415 24089
rect 34793 24055 34851 24061
rect 34793 24021 34805 24055
rect 34839 24021 34851 24055
rect 34793 24015 34851 24021
rect 35713 24055 35771 24061
rect 35713 24021 35725 24055
rect 35759 24052 35771 24055
rect 35894 24052 35900 24064
rect 35759 24024 35900 24052
rect 35759 24021 35771 24024
rect 35713 24015 35771 24021
rect 35894 24012 35900 24024
rect 35952 24052 35958 24064
rect 36556 24052 36584 24148
rect 38010 24052 38016 24064
rect 35952 24024 36584 24052
rect 37971 24024 38016 24052
rect 35952 24012 35958 24024
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 8294 23848 8300 23860
rect 8255 23820 8300 23848
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 37366 23780 37372 23792
rect 37327 23752 37372 23780
rect 37366 23740 37372 23752
rect 37424 23740 37430 23792
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23712 1918 23724
rect 2501 23715 2559 23721
rect 2501 23712 2513 23715
rect 1912 23684 2513 23712
rect 1912 23672 1918 23684
rect 2501 23681 2513 23684
rect 2547 23681 2559 23715
rect 2501 23675 2559 23681
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 10045 23715 10103 23721
rect 10045 23712 10057 23715
rect 9631 23684 10057 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 10045 23681 10057 23684
rect 10091 23712 10103 23715
rect 15654 23712 15660 23724
rect 10091 23684 15660 23712
rect 10091 23681 10103 23684
rect 10045 23675 10103 23681
rect 15654 23672 15660 23684
rect 15712 23672 15718 23724
rect 26418 23672 26424 23724
rect 26476 23712 26482 23724
rect 37829 23715 37887 23721
rect 37829 23712 37841 23715
rect 26476 23684 37841 23712
rect 26476 23672 26482 23684
rect 37829 23681 37841 23684
rect 37875 23681 37887 23715
rect 37829 23675 37887 23681
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 29641 23579 29699 23585
rect 29641 23576 29653 23579
rect 2087 23548 29653 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 29641 23545 29653 23548
rect 29687 23576 29699 23579
rect 29822 23576 29828 23588
rect 29687 23548 29828 23576
rect 29687 23545 29699 23548
rect 29641 23539 29699 23545
rect 29822 23536 29828 23548
rect 29880 23536 29886 23588
rect 3142 23508 3148 23520
rect 3103 23480 3148 23508
rect 3142 23468 3148 23480
rect 3200 23468 3206 23520
rect 35342 23508 35348 23520
rect 35303 23480 35348 23508
rect 35342 23468 35348 23480
rect 35400 23468 35406 23520
rect 38010 23508 38016 23520
rect 37971 23480 38016 23508
rect 38010 23468 38016 23480
rect 38068 23468 38074 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1486 23304 1492 23316
rect 1447 23276 1492 23304
rect 1486 23264 1492 23276
rect 1544 23264 1550 23316
rect 3142 23264 3148 23316
rect 3200 23304 3206 23316
rect 34793 23307 34851 23313
rect 34793 23304 34805 23307
rect 3200 23276 34805 23304
rect 3200 23264 3206 23276
rect 34793 23273 34805 23276
rect 34839 23273 34851 23307
rect 34793 23267 34851 23273
rect 3160 23168 3188 23264
rect 8205 23239 8263 23245
rect 8205 23205 8217 23239
rect 8251 23205 8263 23239
rect 37185 23239 37243 23245
rect 37185 23236 37197 23239
rect 8205 23199 8263 23205
rect 36556 23208 37197 23236
rect 1688 23140 3188 23168
rect 1688 23109 1716 23140
rect 7374 23128 7380 23180
rect 7432 23168 7438 23180
rect 7561 23171 7619 23177
rect 7561 23168 7573 23171
rect 7432 23140 7573 23168
rect 7432 23128 7438 23140
rect 7561 23137 7573 23140
rect 7607 23137 7619 23171
rect 7561 23131 7619 23137
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23069 1731 23103
rect 2130 23100 2136 23112
rect 2091 23072 2136 23100
rect 1673 23063 1731 23069
rect 2130 23060 2136 23072
rect 2188 23100 2194 23112
rect 2777 23103 2835 23109
rect 2777 23100 2789 23103
rect 2188 23072 2789 23100
rect 2188 23060 2194 23072
rect 2777 23069 2789 23072
rect 2823 23069 2835 23103
rect 8220 23100 8248 23199
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 9490 23168 9496 23180
rect 8352 23140 9496 23168
rect 8352 23128 8358 23140
rect 9490 23128 9496 23140
rect 9548 23168 9554 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9548 23140 9689 23168
rect 9548 23128 9554 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 29822 23168 29828 23180
rect 29783 23140 29828 23168
rect 9677 23131 9735 23137
rect 29822 23128 29828 23140
rect 29880 23128 29886 23180
rect 35894 23128 35900 23180
rect 35952 23168 35958 23180
rect 36556 23177 36584 23208
rect 37185 23205 37197 23208
rect 37231 23205 37243 23239
rect 37185 23199 37243 23205
rect 36541 23171 36599 23177
rect 35952 23140 36400 23168
rect 35952 23128 35958 23140
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8220 23072 8953 23100
rect 2777 23063 2835 23069
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 23201 23103 23259 23109
rect 23201 23100 23213 23103
rect 8941 23063 8999 23069
rect 9048 23072 11100 23100
rect 7745 23035 7803 23041
rect 7745 23032 7757 23035
rect 2332 23004 7757 23032
rect 2332 22973 2360 23004
rect 7745 23001 7757 23004
rect 7791 23001 7803 23035
rect 7745 22995 7803 23001
rect 7837 23035 7895 23041
rect 7837 23001 7849 23035
rect 7883 23032 7895 23035
rect 9048 23032 9076 23072
rect 9922 23035 9980 23041
rect 9922 23032 9934 23035
rect 7883 23004 9076 23032
rect 9140 23004 9934 23032
rect 7883 23001 7895 23004
rect 7837 22995 7895 23001
rect 9140 22973 9168 23004
rect 9922 23001 9934 23004
rect 9968 23001 9980 23035
rect 9922 22995 9980 23001
rect 11072 22973 11100 23072
rect 16546 23072 23213 23100
rect 2317 22967 2375 22973
rect 2317 22933 2329 22967
rect 2363 22933 2375 22967
rect 2317 22927 2375 22933
rect 9125 22967 9183 22973
rect 9125 22933 9137 22967
rect 9171 22933 9183 22967
rect 9125 22927 9183 22933
rect 11057 22967 11115 22973
rect 11057 22933 11069 22967
rect 11103 22964 11115 22967
rect 16546 22964 16574 23072
rect 23201 23069 23213 23072
rect 23247 23069 23259 23103
rect 23382 23100 23388 23112
rect 23343 23072 23388 23100
rect 23201 23063 23259 23069
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 30006 23100 30012 23112
rect 29967 23072 30012 23100
rect 30006 23060 30012 23072
rect 30064 23060 30070 23112
rect 36372 23109 36400 23140
rect 36541 23137 36553 23171
rect 36587 23137 36599 23171
rect 36541 23131 36599 23137
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23100 30251 23103
rect 31757 23103 31815 23109
rect 31757 23100 31769 23103
rect 30239 23072 31769 23100
rect 30239 23069 30251 23072
rect 30193 23063 30251 23069
rect 31757 23069 31769 23072
rect 31803 23069 31815 23103
rect 31757 23063 31815 23069
rect 34977 23103 35035 23109
rect 34977 23069 34989 23103
rect 35023 23100 35035 23103
rect 36173 23103 36231 23109
rect 36173 23100 36185 23103
rect 35023 23072 36185 23100
rect 35023 23069 35035 23072
rect 34977 23063 35035 23069
rect 36173 23069 36185 23072
rect 36219 23069 36231 23103
rect 36173 23063 36231 23069
rect 36357 23103 36415 23109
rect 36357 23069 36369 23103
rect 36403 23069 36415 23103
rect 37366 23100 37372 23112
rect 37327 23072 37372 23100
rect 36357 23063 36415 23069
rect 37366 23060 37372 23072
rect 37424 23060 37430 23112
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23069 37887 23103
rect 37829 23063 37887 23069
rect 21269 23035 21327 23041
rect 21269 23001 21281 23035
rect 21315 23001 21327 23035
rect 21450 23032 21456 23044
rect 21411 23004 21456 23032
rect 21269 22995 21327 23001
rect 11103 22936 16574 22964
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 21284 22964 21312 22995
rect 21450 22992 21456 23004
rect 21508 22992 21514 23044
rect 37844 23032 37872 23063
rect 31956 23004 37872 23032
rect 22002 22964 22008 22976
rect 21140 22936 22008 22964
rect 21140 22924 21146 22936
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 23569 22967 23627 22973
rect 23569 22933 23581 22967
rect 23615 22964 23627 22967
rect 24946 22964 24952 22976
rect 23615 22936 24952 22964
rect 23615 22933 23627 22936
rect 23569 22927 23627 22933
rect 24946 22924 24952 22936
rect 25004 22924 25010 22976
rect 31956 22973 31984 23004
rect 31941 22967 31999 22973
rect 31941 22933 31953 22967
rect 31987 22933 31999 22967
rect 38010 22964 38016 22976
rect 37971 22936 38016 22964
rect 31941 22927 31999 22933
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 9490 22760 9496 22772
rect 9451 22732 9496 22760
rect 9490 22720 9496 22732
rect 9548 22720 9554 22772
rect 23293 22763 23351 22769
rect 23293 22729 23305 22763
rect 23339 22760 23351 22763
rect 23382 22760 23388 22772
rect 23339 22732 23388 22760
rect 23339 22729 23351 22732
rect 23293 22723 23351 22729
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 1719 22596 3372 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 3344 22497 3372 22596
rect 22002 22584 22008 22636
rect 22060 22624 22066 22636
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 22060 22596 23121 22624
rect 22060 22584 22066 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 24946 22624 24952 22636
rect 24907 22596 24952 22624
rect 23109 22587 23167 22593
rect 23124 22556 23152 22587
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 30006 22584 30012 22636
rect 30064 22624 30070 22636
rect 30285 22627 30343 22633
rect 30285 22624 30297 22627
rect 30064 22596 30297 22624
rect 30064 22584 30070 22596
rect 30285 22593 30297 22596
rect 30331 22593 30343 22627
rect 34514 22624 34520 22636
rect 34475 22596 34520 22624
rect 30285 22587 30343 22593
rect 34514 22584 34520 22596
rect 34572 22584 34578 22636
rect 37274 22584 37280 22636
rect 37332 22624 37338 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37332 22596 37841 22624
rect 37332 22584 37338 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23124 22528 23857 22556
rect 23845 22525 23857 22528
rect 23891 22556 23903 22559
rect 26326 22556 26332 22568
rect 23891 22528 26332 22556
rect 23891 22525 23903 22528
rect 23845 22519 23903 22525
rect 26326 22516 26332 22528
rect 26384 22516 26390 22568
rect 29546 22516 29552 22568
rect 29604 22556 29610 22568
rect 30101 22559 30159 22565
rect 30101 22556 30113 22559
rect 29604 22528 30113 22556
rect 29604 22516 29610 22528
rect 30101 22525 30113 22528
rect 30147 22525 30159 22559
rect 37366 22556 37372 22568
rect 37327 22528 37372 22556
rect 30101 22519 30159 22525
rect 37366 22516 37372 22528
rect 37424 22516 37430 22568
rect 3329 22491 3387 22497
rect 3329 22457 3341 22491
rect 3375 22488 3387 22491
rect 34333 22491 34391 22497
rect 34333 22488 34345 22491
rect 3375 22460 34345 22488
rect 3375 22457 3387 22460
rect 3329 22451 3387 22457
rect 34333 22457 34345 22460
rect 34379 22457 34391 22491
rect 34333 22451 34391 22457
rect 1486 22420 1492 22432
rect 1447 22392 1492 22420
rect 1486 22380 1492 22392
rect 1544 22380 1550 22432
rect 1854 22380 1860 22432
rect 1912 22420 1918 22432
rect 2133 22423 2191 22429
rect 2133 22420 2145 22423
rect 1912 22392 2145 22420
rect 1912 22380 1918 22392
rect 2133 22389 2145 22392
rect 2179 22389 2191 22423
rect 2133 22383 2191 22389
rect 2777 22423 2835 22429
rect 2777 22389 2789 22423
rect 2823 22420 2835 22423
rect 3878 22420 3884 22432
rect 2823 22392 3884 22420
rect 2823 22389 2835 22392
rect 2777 22383 2835 22389
rect 3878 22380 3884 22392
rect 3936 22380 3942 22432
rect 25130 22420 25136 22432
rect 25091 22392 25136 22420
rect 25130 22380 25136 22392
rect 25188 22380 25194 22432
rect 29546 22420 29552 22432
rect 29507 22392 29552 22420
rect 29546 22380 29552 22392
rect 29604 22380 29610 22432
rect 30466 22420 30472 22432
rect 30427 22392 30472 22420
rect 30466 22380 30472 22392
rect 30524 22380 30530 22432
rect 38013 22423 38071 22429
rect 38013 22389 38025 22423
rect 38059 22420 38071 22423
rect 38102 22420 38108 22432
rect 38059 22392 38108 22420
rect 38059 22389 38071 22392
rect 38013 22383 38071 22389
rect 38102 22380 38108 22392
rect 38160 22380 38166 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 21082 22216 21088 22228
rect 21043 22188 21088 22216
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 25188 22188 26234 22216
rect 25188 22176 25194 22188
rect 26206 22148 26234 22188
rect 34514 22176 34520 22228
rect 34572 22216 34578 22228
rect 35713 22219 35771 22225
rect 35713 22216 35725 22219
rect 34572 22188 35725 22216
rect 34572 22176 34578 22188
rect 35713 22185 35725 22188
rect 35759 22185 35771 22219
rect 35713 22179 35771 22185
rect 26206 22120 37872 22148
rect 29546 22080 29552 22092
rect 16316 22052 29552 22080
rect 1854 22012 1860 22024
rect 1815 21984 1860 22012
rect 1854 21972 1860 21984
rect 1912 21972 1918 22024
rect 2501 22015 2559 22021
rect 2501 21981 2513 22015
rect 2547 22012 2559 22015
rect 2774 22012 2780 22024
rect 2547 21984 2780 22012
rect 2547 21981 2559 21984
rect 2501 21975 2559 21981
rect 2774 21972 2780 21984
rect 2832 22012 2838 22024
rect 3145 22015 3203 22021
rect 3145 22012 3157 22015
rect 2832 21984 3157 22012
rect 2832 21972 2838 21984
rect 3145 21981 3157 21984
rect 3191 21981 3203 22015
rect 16316 22012 16344 22052
rect 29546 22040 29552 22052
rect 29604 22040 29610 22092
rect 37274 22080 37280 22092
rect 36280 22052 37280 22080
rect 3145 21975 3203 21981
rect 6886 21984 16344 22012
rect 16393 22015 16451 22021
rect 2041 21947 2099 21953
rect 2041 21913 2053 21947
rect 2087 21944 2099 21947
rect 6886 21944 6914 21984
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 20349 22015 20407 22021
rect 16439 21984 16574 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 2087 21916 6914 21944
rect 2087 21913 2099 21916
rect 2041 21907 2099 21913
rect 15102 21904 15108 21956
rect 15160 21944 15166 21956
rect 16126 21947 16184 21953
rect 16126 21944 16138 21947
rect 15160 21916 16138 21944
rect 15160 21904 15166 21916
rect 16126 21913 16138 21916
rect 16172 21913 16184 21947
rect 16126 21907 16184 21913
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21876 2743 21879
rect 3970 21876 3976 21888
rect 2731 21848 3976 21876
rect 2731 21845 2743 21848
rect 2685 21839 2743 21845
rect 3970 21836 3976 21848
rect 4028 21836 4034 21888
rect 15013 21879 15071 21885
rect 15013 21845 15025 21879
rect 15059 21876 15071 21879
rect 15194 21876 15200 21888
rect 15059 21848 15200 21876
rect 15059 21845 15071 21848
rect 15013 21839 15071 21845
rect 15194 21836 15200 21848
rect 15252 21836 15258 21888
rect 16546 21876 16574 21984
rect 20349 21981 20361 22015
rect 20395 22012 20407 22015
rect 21082 22012 21088 22024
rect 20395 21984 21088 22012
rect 20395 21981 20407 21984
rect 20349 21975 20407 21981
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 30466 21972 30472 22024
rect 30524 22012 30530 22024
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 30524 21984 32229 22012
rect 30524 21972 30530 21984
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 32217 21975 32275 21981
rect 35894 21972 35900 22024
rect 35952 22012 35958 22024
rect 35952 21984 35997 22012
rect 35952 21972 35958 21984
rect 36078 21972 36084 22024
rect 36136 22012 36142 22024
rect 36136 21984 36181 22012
rect 36136 21972 36142 21984
rect 36280 21944 36308 22052
rect 37274 22040 37280 22052
rect 37332 22040 37338 22092
rect 37366 22012 37372 22024
rect 37292 21984 37372 22012
rect 35866 21916 36308 21944
rect 36725 21947 36783 21953
rect 16945 21879 17003 21885
rect 16945 21876 16957 21879
rect 16546 21848 16957 21876
rect 16945 21845 16957 21848
rect 16991 21876 17003 21879
rect 17126 21876 17132 21888
rect 16991 21848 17132 21876
rect 16991 21845 17003 21848
rect 16945 21839 17003 21845
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 20533 21879 20591 21885
rect 20533 21845 20545 21879
rect 20579 21876 20591 21879
rect 20714 21876 20720 21888
rect 20579 21848 20720 21876
rect 20579 21845 20591 21848
rect 20533 21839 20591 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 32401 21879 32459 21885
rect 32401 21845 32413 21879
rect 32447 21876 32459 21879
rect 35866 21876 35894 21916
rect 36725 21913 36737 21947
rect 36771 21944 36783 21947
rect 37292 21944 37320 21984
rect 37366 21972 37372 21984
rect 37424 21972 37430 22024
rect 37844 22021 37872 22120
rect 37829 22015 37887 22021
rect 37829 21981 37841 22015
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 36771 21916 37320 21944
rect 36771 21913 36783 21916
rect 36725 21907 36783 21913
rect 32447 21848 35894 21876
rect 32447 21845 32459 21848
rect 32401 21839 32459 21845
rect 36078 21836 36084 21888
rect 36136 21876 36142 21888
rect 37185 21879 37243 21885
rect 37185 21876 37197 21879
rect 36136 21848 37197 21876
rect 36136 21836 36142 21848
rect 37185 21845 37197 21848
rect 37231 21845 37243 21879
rect 38010 21876 38016 21888
rect 37971 21848 38016 21876
rect 37185 21839 37243 21845
rect 38010 21836 38016 21848
rect 38068 21836 38074 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 3878 21672 3884 21684
rect 1688 21644 3884 21672
rect 1688 21545 1716 21644
rect 3878 21632 3884 21644
rect 3936 21632 3942 21684
rect 4617 21675 4675 21681
rect 4617 21641 4629 21675
rect 4663 21672 4675 21675
rect 8294 21672 8300 21684
rect 4663 21644 8300 21672
rect 4663 21641 4675 21644
rect 4617 21635 4675 21641
rect 4632 21604 4660 21635
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 15013 21675 15071 21681
rect 15013 21641 15025 21675
rect 15059 21672 15071 21675
rect 15102 21672 15108 21684
rect 15059 21644 15108 21672
rect 15059 21641 15071 21644
rect 15013 21635 15071 21641
rect 15102 21632 15108 21644
rect 15160 21632 15166 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 20530 21672 20536 21684
rect 15252 21644 20536 21672
rect 15252 21632 15258 21644
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 21910 21632 21916 21684
rect 21968 21672 21974 21684
rect 24946 21672 24952 21684
rect 21968 21644 24952 21672
rect 21968 21632 21974 21644
rect 24946 21632 24952 21644
rect 25004 21672 25010 21684
rect 25225 21675 25283 21681
rect 25225 21672 25237 21675
rect 25004 21644 25237 21672
rect 25004 21632 25010 21644
rect 25225 21641 25237 21644
rect 25271 21641 25283 21675
rect 25225 21635 25283 21641
rect 25498 21632 25504 21684
rect 25556 21672 25562 21684
rect 25958 21672 25964 21684
rect 25556 21644 25964 21672
rect 25556 21632 25562 21644
rect 25958 21632 25964 21644
rect 26016 21672 26022 21684
rect 26237 21675 26295 21681
rect 26237 21672 26249 21675
rect 26016 21644 26249 21672
rect 26016 21632 26022 21644
rect 26237 21641 26249 21644
rect 26283 21641 26295 21675
rect 26237 21635 26295 21641
rect 2700 21576 4660 21604
rect 2700 21545 2728 21576
rect 2958 21545 2964 21548
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 2685 21539 2743 21545
rect 2685 21505 2697 21539
rect 2731 21505 2743 21539
rect 2685 21499 2743 21505
rect 2952 21499 2964 21545
rect 3016 21536 3022 21548
rect 14829 21539 14887 21545
rect 3016 21508 3052 21536
rect 2958 21496 2964 21499
rect 3016 21496 3022 21508
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15194 21536 15200 21548
rect 14875 21508 15200 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21536 20591 21539
rect 20622 21536 20628 21548
rect 20579 21508 20628 21536
rect 20579 21505 20591 21508
rect 20533 21499 20591 21505
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 25406 21536 25412 21548
rect 25367 21508 25412 21536
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 26418 21536 26424 21548
rect 26379 21508 26424 21536
rect 26418 21496 26424 21508
rect 26476 21536 26482 21548
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 26476 21508 26985 21536
rect 26476 21496 26482 21508
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 28442 21536 28448 21548
rect 28403 21508 28448 21536
rect 26973 21499 27031 21505
rect 28442 21496 28448 21508
rect 28500 21496 28506 21548
rect 37826 21536 37832 21548
rect 37787 21508 37832 21536
rect 37826 21496 37832 21508
rect 37884 21496 37890 21548
rect 20346 21468 20352 21480
rect 20307 21440 20352 21468
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 20717 21471 20775 21477
rect 20717 21437 20729 21471
rect 20763 21468 20775 21471
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 20763 21440 21833 21468
rect 20763 21437 20775 21440
rect 20717 21431 20775 21437
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 22097 21471 22155 21477
rect 22097 21437 22109 21471
rect 22143 21468 22155 21471
rect 37458 21468 37464 21480
rect 22143 21440 37464 21468
rect 22143 21437 22155 21440
rect 22097 21431 22155 21437
rect 37458 21428 37464 21440
rect 37516 21428 37522 21480
rect 1486 21332 1492 21344
rect 1447 21304 1492 21332
rect 1486 21292 1492 21304
rect 1544 21292 1550 21344
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 2133 21335 2191 21341
rect 2133 21332 2145 21335
rect 1912 21304 2145 21332
rect 1912 21292 1918 21304
rect 2133 21301 2145 21304
rect 2179 21301 2191 21335
rect 2133 21295 2191 21301
rect 4065 21335 4123 21341
rect 4065 21301 4077 21335
rect 4111 21332 4123 21335
rect 4614 21332 4620 21344
rect 4111 21304 4620 21332
rect 4111 21301 4123 21304
rect 4065 21295 4123 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 27157 21335 27215 21341
rect 27157 21301 27169 21335
rect 27203 21332 27215 21335
rect 27614 21332 27620 21344
rect 27203 21304 27620 21332
rect 27203 21301 27215 21304
rect 27157 21295 27215 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 28721 21335 28779 21341
rect 28721 21301 28733 21335
rect 28767 21332 28779 21335
rect 30098 21332 30104 21344
rect 28767 21304 30104 21332
rect 28767 21301 28779 21304
rect 28721 21295 28779 21301
rect 30098 21292 30104 21304
rect 30156 21292 30162 21344
rect 38013 21335 38071 21341
rect 38013 21301 38025 21335
rect 38059 21332 38071 21335
rect 38102 21332 38108 21344
rect 38059 21304 38108 21332
rect 38059 21301 38071 21304
rect 38013 21295 38071 21301
rect 38102 21292 38108 21304
rect 38160 21292 38166 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 2958 21128 2964 21140
rect 2919 21100 2964 21128
rect 2958 21088 2964 21100
rect 3016 21088 3022 21140
rect 4614 21088 4620 21140
rect 4672 21128 4678 21140
rect 20346 21128 20352 21140
rect 4672 21100 20352 21128
rect 4672 21088 4678 21100
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 25406 21088 25412 21140
rect 25464 21128 25470 21140
rect 26513 21131 26571 21137
rect 26513 21128 26525 21131
rect 25464 21100 26525 21128
rect 25464 21088 25470 21100
rect 26513 21097 26525 21100
rect 26559 21128 26571 21131
rect 28442 21128 28448 21140
rect 26559 21100 28448 21128
rect 26559 21097 26571 21100
rect 26513 21091 26571 21097
rect 28442 21088 28448 21100
rect 28500 21088 28506 21140
rect 3789 21063 3847 21069
rect 3789 21029 3801 21063
rect 3835 21029 3847 21063
rect 3789 21023 3847 21029
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20924 3203 20927
rect 3804 20924 3832 21023
rect 3878 21020 3884 21072
rect 3936 21060 3942 21072
rect 15194 21060 15200 21072
rect 3936 21032 14688 21060
rect 15155 21032 15200 21060
rect 3936 21020 3942 21032
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 4249 20995 4307 21001
rect 4249 20992 4261 20995
rect 4028 20964 4261 20992
rect 4028 20952 4034 20964
rect 4249 20961 4261 20964
rect 4295 20961 4307 20995
rect 4249 20955 4307 20961
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20992 4491 20995
rect 7374 20992 7380 21004
rect 4479 20964 7380 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 12894 20952 12900 21004
rect 12952 20992 12958 21004
rect 14553 20995 14611 21001
rect 14553 20992 14565 20995
rect 12952 20964 14565 20992
rect 12952 20952 12958 20964
rect 14553 20961 14565 20964
rect 14599 20961 14611 20995
rect 14660 20992 14688 21032
rect 15194 21020 15200 21032
rect 15252 21020 15258 21072
rect 25590 21020 25596 21072
rect 25648 21060 25654 21072
rect 26329 21063 26387 21069
rect 26329 21060 26341 21063
rect 25648 21032 26341 21060
rect 25648 21020 25654 21032
rect 26329 21029 26341 21032
rect 26375 21029 26387 21063
rect 26329 21023 26387 21029
rect 35529 21063 35587 21069
rect 35529 21029 35541 21063
rect 35575 21029 35587 21063
rect 35529 21023 35587 21029
rect 35544 20992 35572 21023
rect 14660 20964 35572 20992
rect 14553 20955 14611 20961
rect 3191 20896 3832 20924
rect 4157 20927 4215 20933
rect 3191 20893 3203 20896
rect 3145 20887 3203 20893
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 4614 20924 4620 20936
rect 4203 20896 4620 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 7006 20924 7012 20936
rect 6967 20896 7012 20924
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 15286 20924 15292 20936
rect 14875 20896 15292 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 15654 20924 15660 20936
rect 15615 20896 15660 20924
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 20530 20924 20536 20936
rect 20491 20896 20536 20924
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 35713 20927 35771 20933
rect 35713 20893 35725 20927
rect 35759 20924 35771 20927
rect 36906 20924 36912 20936
rect 35759 20896 36912 20924
rect 35759 20893 35771 20896
rect 35713 20887 35771 20893
rect 36906 20884 36912 20896
rect 36964 20884 36970 20936
rect 37090 20884 37096 20936
rect 37148 20924 37154 20936
rect 37369 20927 37427 20933
rect 37369 20924 37381 20927
rect 37148 20896 37381 20924
rect 37148 20884 37154 20896
rect 37369 20893 37381 20896
rect 37415 20893 37427 20927
rect 37369 20887 37427 20893
rect 37458 20884 37464 20936
rect 37516 20924 37522 20936
rect 37829 20927 37887 20933
rect 37829 20924 37841 20927
rect 37516 20896 37841 20924
rect 37516 20884 37522 20896
rect 37829 20893 37841 20896
rect 37875 20893 37887 20927
rect 37829 20887 37887 20893
rect 1854 20856 1860 20868
rect 1815 20828 1860 20856
rect 1854 20816 1860 20828
rect 1912 20816 1918 20868
rect 2038 20856 2044 20868
rect 1999 20828 2044 20856
rect 2038 20816 2044 20828
rect 2096 20816 2102 20868
rect 26053 20859 26111 20865
rect 26053 20825 26065 20859
rect 26099 20856 26111 20859
rect 26142 20856 26148 20868
rect 26099 20828 26148 20856
rect 26099 20825 26111 20828
rect 26053 20819 26111 20825
rect 26142 20816 26148 20828
rect 26200 20816 26206 20868
rect 36725 20859 36783 20865
rect 36725 20825 36737 20859
rect 36771 20856 36783 20859
rect 37108 20856 37136 20884
rect 36771 20828 37136 20856
rect 36771 20825 36783 20828
rect 36725 20819 36783 20825
rect 7190 20788 7196 20800
rect 7151 20760 7196 20788
rect 7190 20748 7196 20760
rect 7248 20748 7254 20800
rect 12526 20748 12532 20800
rect 12584 20788 12590 20800
rect 14737 20791 14795 20797
rect 14737 20788 14749 20791
rect 12584 20760 14749 20788
rect 12584 20748 12590 20760
rect 14737 20757 14749 20760
rect 14783 20757 14795 20791
rect 17126 20788 17132 20800
rect 17087 20760 17132 20788
rect 14737 20751 14795 20757
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 20901 20791 20959 20797
rect 20901 20757 20913 20791
rect 20947 20788 20959 20791
rect 22002 20788 22008 20800
rect 20947 20760 22008 20788
rect 20947 20757 20959 20760
rect 20901 20751 20959 20757
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 25590 20788 25596 20800
rect 25551 20760 25596 20788
rect 25590 20748 25596 20760
rect 25648 20748 25654 20800
rect 37185 20791 37243 20797
rect 37185 20757 37197 20791
rect 37231 20788 37243 20791
rect 37274 20788 37280 20800
rect 37231 20760 37280 20788
rect 37231 20757 37243 20760
rect 37185 20751 37243 20757
rect 37274 20748 37280 20760
rect 37332 20748 37338 20800
rect 38010 20788 38016 20800
rect 37971 20760 38016 20788
rect 38010 20748 38016 20760
rect 38068 20748 38074 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6825 20587 6883 20593
rect 6825 20553 6837 20587
rect 6871 20584 6883 20587
rect 7006 20584 7012 20596
rect 6871 20556 7012 20584
rect 6871 20553 6883 20556
rect 6825 20547 6883 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 15565 20587 15623 20593
rect 15565 20553 15577 20587
rect 15611 20584 15623 20587
rect 15654 20584 15660 20596
rect 15611 20556 15660 20584
rect 15611 20553 15623 20556
rect 15565 20547 15623 20553
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 26418 20584 26424 20596
rect 26379 20556 26424 20584
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 32585 20587 32643 20593
rect 32585 20553 32597 20587
rect 32631 20584 32643 20587
rect 37826 20584 37832 20596
rect 32631 20556 37832 20584
rect 32631 20553 32643 20556
rect 32585 20547 32643 20553
rect 37826 20544 37832 20556
rect 37884 20544 37890 20596
rect 2038 20476 2044 20528
rect 2096 20516 2102 20528
rect 2096 20488 16574 20516
rect 2096 20476 2102 20488
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20417 1731 20451
rect 2130 20448 2136 20460
rect 2091 20420 2136 20448
rect 1673 20411 1731 20417
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 1688 20244 1716 20411
rect 2130 20408 2136 20420
rect 2188 20448 2194 20460
rect 2777 20451 2835 20457
rect 2777 20448 2789 20451
rect 2188 20420 2789 20448
rect 2188 20408 2194 20420
rect 2777 20417 2789 20420
rect 2823 20417 2835 20451
rect 2777 20411 2835 20417
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20448 7251 20451
rect 7466 20448 7472 20460
rect 7239 20420 7472 20448
rect 7239 20417 7251 20420
rect 7193 20411 7251 20417
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 7285 20383 7343 20389
rect 7285 20380 7297 20383
rect 6886 20352 7297 20380
rect 2317 20315 2375 20321
rect 2317 20281 2329 20315
rect 2363 20312 2375 20315
rect 6886 20312 6914 20352
rect 7285 20349 7297 20352
rect 7331 20349 7343 20383
rect 7285 20343 7343 20349
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 7432 20352 7477 20380
rect 7432 20340 7438 20352
rect 2363 20284 6914 20312
rect 16546 20312 16574 20488
rect 20714 20448 20720 20460
rect 20627 20420 20720 20448
rect 20714 20408 20720 20420
rect 20772 20448 20778 20460
rect 21082 20448 21088 20460
rect 20772 20420 21088 20448
rect 20772 20408 20778 20420
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 30282 20408 30288 20460
rect 30340 20448 30346 20460
rect 30377 20451 30435 20457
rect 30377 20448 30389 20451
rect 30340 20420 30389 20448
rect 30340 20408 30346 20420
rect 30377 20417 30389 20420
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 32401 20451 32459 20457
rect 32401 20448 32413 20451
rect 30607 20420 32413 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 32401 20417 32413 20420
rect 32447 20417 32459 20451
rect 32401 20411 32459 20417
rect 32582 20408 32588 20460
rect 32640 20448 32646 20460
rect 37829 20451 37887 20457
rect 37829 20448 37841 20451
rect 32640 20420 37841 20448
rect 32640 20408 32646 20420
rect 37829 20417 37841 20420
rect 37875 20417 37887 20451
rect 37829 20411 37887 20417
rect 20530 20380 20536 20392
rect 20491 20352 20536 20380
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 25590 20340 25596 20392
rect 25648 20380 25654 20392
rect 25961 20383 26019 20389
rect 25961 20380 25973 20383
rect 25648 20352 25973 20380
rect 25648 20340 25654 20352
rect 25961 20349 25973 20352
rect 26007 20349 26019 20383
rect 29641 20383 29699 20389
rect 29641 20380 29653 20383
rect 25961 20343 26019 20349
rect 26068 20352 29653 20380
rect 26068 20312 26096 20352
rect 29641 20349 29653 20352
rect 29687 20380 29699 20383
rect 30193 20383 30251 20389
rect 30193 20380 30205 20383
rect 29687 20352 30205 20380
rect 29687 20349 29699 20352
rect 29641 20343 29699 20349
rect 30193 20349 30205 20352
rect 30239 20349 30251 20383
rect 30193 20343 30251 20349
rect 16546 20284 26096 20312
rect 2363 20281 2375 20284
rect 2317 20275 2375 20281
rect 26142 20272 26148 20324
rect 26200 20312 26206 20324
rect 26237 20315 26295 20321
rect 26237 20312 26249 20315
rect 26200 20284 26249 20312
rect 26200 20272 26206 20284
rect 26237 20281 26249 20284
rect 26283 20281 26295 20315
rect 26237 20275 26295 20281
rect 3421 20247 3479 20253
rect 3421 20244 3433 20247
rect 1688 20216 3433 20244
rect 3421 20213 3433 20216
rect 3467 20244 3479 20247
rect 11698 20244 11704 20256
rect 3467 20216 11704 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 25501 20247 25559 20253
rect 25501 20213 25513 20247
rect 25547 20244 25559 20247
rect 25590 20244 25596 20256
rect 25547 20216 25596 20244
rect 25547 20213 25559 20216
rect 25501 20207 25559 20213
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 37182 20204 37188 20256
rect 37240 20244 37246 20256
rect 38013 20247 38071 20253
rect 38013 20244 38025 20247
rect 37240 20216 38025 20244
rect 37240 20204 37246 20216
rect 38013 20213 38025 20216
rect 38059 20213 38071 20247
rect 38013 20207 38071 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 8294 20040 8300 20052
rect 6932 20012 8300 20040
rect 6932 19913 6960 20012
rect 8294 20000 8300 20012
rect 8352 20040 8358 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8352 20012 8953 20040
rect 8352 20000 8358 20012
rect 8941 20009 8953 20012
rect 8987 20040 8999 20043
rect 10505 20043 10563 20049
rect 10505 20040 10517 20043
rect 8987 20012 10517 20040
rect 8987 20009 8999 20012
rect 8941 20003 8999 20009
rect 10505 20009 10517 20012
rect 10551 20009 10563 20043
rect 10505 20003 10563 20009
rect 6917 19907 6975 19913
rect 6917 19873 6929 19907
rect 6963 19873 6975 19907
rect 10520 19904 10548 20003
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 35161 20043 35219 20049
rect 35161 20040 35173 20043
rect 11756 20012 35173 20040
rect 11756 20000 11762 20012
rect 35161 20009 35173 20012
rect 35207 20009 35219 20043
rect 36906 20040 36912 20052
rect 36867 20012 36912 20040
rect 35161 20003 35219 20009
rect 36906 20000 36912 20012
rect 36964 20000 36970 20052
rect 11057 19907 11115 19913
rect 11057 19904 11069 19907
rect 10520 19876 11069 19904
rect 6917 19867 6975 19873
rect 11057 19873 11069 19876
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 22002 19864 22008 19916
rect 22060 19904 22066 19916
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 22060 19876 22293 19904
rect 22060 19864 22066 19876
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 37274 19904 37280 19916
rect 37235 19876 37280 19904
rect 22281 19867 22339 19873
rect 37274 19864 37280 19876
rect 37332 19864 37338 19916
rect 7190 19845 7196 19848
rect 7184 19836 7196 19845
rect 7151 19808 7196 19836
rect 7184 19799 7196 19808
rect 7190 19796 7196 19799
rect 7248 19796 7254 19848
rect 7466 19796 7472 19848
rect 7524 19836 7530 19848
rect 20530 19836 20536 19848
rect 7524 19808 20536 19836
rect 7524 19796 7530 19808
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19768 1918 19780
rect 2501 19771 2559 19777
rect 2501 19768 2513 19771
rect 1912 19740 2513 19768
rect 1912 19728 1918 19740
rect 2501 19737 2513 19740
rect 2547 19737 2559 19771
rect 2501 19731 2559 19737
rect 1946 19700 1952 19712
rect 1907 19672 1952 19700
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 8312 19709 8340 19808
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19836 22615 19839
rect 34514 19836 34520 19848
rect 22603 19808 34520 19836
rect 22603 19805 22615 19808
rect 22557 19799 22615 19805
rect 34514 19796 34520 19808
rect 34572 19796 34578 19848
rect 36262 19796 36268 19848
rect 36320 19836 36326 19848
rect 37093 19839 37151 19845
rect 37093 19836 37105 19839
rect 36320 19808 37105 19836
rect 36320 19796 36326 19808
rect 37093 19805 37105 19808
rect 37139 19805 37151 19839
rect 37093 19799 37151 19805
rect 37829 19839 37887 19845
rect 37829 19805 37841 19839
rect 37875 19805 37887 19839
rect 37829 19799 37887 19805
rect 11324 19771 11382 19777
rect 11324 19737 11336 19771
rect 11370 19768 11382 19771
rect 11514 19768 11520 19780
rect 11370 19740 11520 19768
rect 11370 19737 11382 19740
rect 11324 19731 11382 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 35253 19771 35311 19777
rect 35253 19737 35265 19771
rect 35299 19768 35311 19771
rect 36538 19768 36544 19780
rect 35299 19740 36544 19768
rect 35299 19737 35311 19740
rect 35253 19731 35311 19737
rect 36538 19728 36544 19740
rect 36596 19728 36602 19780
rect 37844 19768 37872 19799
rect 36740 19740 37872 19768
rect 8297 19703 8355 19709
rect 8297 19669 8309 19703
rect 8343 19669 8355 19703
rect 12434 19700 12440 19712
rect 12395 19672 12440 19700
rect 8297 19663 8355 19669
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 30190 19660 30196 19712
rect 30248 19700 30254 19712
rect 36740 19700 36768 19740
rect 38010 19700 38016 19712
rect 30248 19672 36768 19700
rect 37971 19672 38016 19700
rect 30248 19660 30254 19672
rect 38010 19660 38016 19672
rect 38068 19660 38074 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 32582 19496 32588 19508
rect 32543 19468 32588 19496
rect 32582 19456 32588 19468
rect 32640 19456 32646 19508
rect 35713 19499 35771 19505
rect 35713 19465 35725 19499
rect 35759 19496 35771 19499
rect 36262 19496 36268 19508
rect 35759 19468 36268 19496
rect 35759 19465 35771 19468
rect 35713 19459 35771 19465
rect 36262 19456 36268 19468
rect 36320 19456 36326 19508
rect 36538 19456 36544 19508
rect 36596 19496 36602 19508
rect 37277 19499 37335 19505
rect 37277 19496 37289 19499
rect 36596 19468 37289 19496
rect 36596 19456 36602 19468
rect 37277 19465 37289 19468
rect 37323 19465 37335 19499
rect 37277 19459 37335 19465
rect 12526 19428 12532 19440
rect 6886 19400 12532 19428
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19360 2007 19363
rect 6886 19360 6914 19400
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 30098 19388 30104 19440
rect 30156 19428 30162 19440
rect 35342 19428 35348 19440
rect 30156 19400 35348 19428
rect 30156 19388 30162 19400
rect 35342 19388 35348 19400
rect 35400 19428 35406 19440
rect 35400 19400 35572 19428
rect 35400 19388 35406 19400
rect 11698 19360 11704 19372
rect 1995 19332 6914 19360
rect 11659 19332 11704 19360
rect 1995 19329 2007 19332
rect 1949 19323 2007 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19360 22523 19363
rect 30190 19360 30196 19372
rect 22511 19332 30196 19360
rect 22511 19329 22523 19332
rect 22465 19323 22523 19329
rect 30190 19320 30196 19332
rect 30248 19320 30254 19372
rect 30282 19320 30288 19372
rect 30340 19360 30346 19372
rect 35544 19369 35572 19400
rect 30469 19363 30527 19369
rect 30340 19332 30385 19360
rect 30340 19320 30346 19332
rect 30469 19329 30481 19363
rect 30515 19360 30527 19363
rect 32401 19363 32459 19369
rect 32401 19360 32413 19363
rect 30515 19332 32413 19360
rect 30515 19329 30527 19332
rect 30469 19323 30527 19329
rect 32401 19329 32413 19332
rect 32447 19329 32459 19363
rect 32401 19323 32459 19329
rect 35529 19363 35587 19369
rect 35529 19329 35541 19363
rect 35575 19360 35587 19363
rect 35575 19332 35894 19360
rect 35575 19329 35587 19332
rect 35529 19323 35587 19329
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19292 2286 19304
rect 2685 19295 2743 19301
rect 2685 19292 2697 19295
rect 2280 19264 2697 19292
rect 2280 19252 2286 19264
rect 2685 19261 2697 19264
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 20956 19264 22201 19292
rect 20956 19252 20962 19264
rect 22189 19261 22201 19264
rect 22235 19261 22247 19295
rect 22189 19255 22247 19261
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19261 30159 19295
rect 30101 19255 30159 19261
rect 1946 19184 1952 19236
rect 2004 19224 2010 19236
rect 29549 19227 29607 19233
rect 29549 19224 29561 19227
rect 2004 19196 29561 19224
rect 2004 19184 2010 19196
rect 29549 19193 29561 19196
rect 29595 19224 29607 19227
rect 30116 19224 30144 19255
rect 29595 19196 30144 19224
rect 29595 19193 29607 19196
rect 29549 19187 29607 19193
rect 35866 19156 35894 19332
rect 36262 19320 36268 19372
rect 36320 19360 36326 19372
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 36320 19332 37473 19360
rect 36320 19320 36326 19332
rect 37461 19329 37473 19332
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 37366 19252 37372 19304
rect 37424 19292 37430 19304
rect 37645 19295 37703 19301
rect 37645 19292 37657 19295
rect 37424 19264 37657 19292
rect 37424 19252 37430 19264
rect 37645 19261 37657 19264
rect 37691 19261 37703 19295
rect 37645 19255 37703 19261
rect 36173 19159 36231 19165
rect 36173 19156 36185 19159
rect 35866 19128 36185 19156
rect 36173 19125 36185 19128
rect 36219 19125 36231 19159
rect 36173 19119 36231 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 11425 18955 11483 18961
rect 11425 18921 11437 18955
rect 11471 18952 11483 18955
rect 11698 18952 11704 18964
rect 11471 18924 11704 18952
rect 11471 18921 11483 18924
rect 11425 18915 11483 18921
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 26326 18912 26332 18964
rect 26384 18952 26390 18964
rect 26421 18955 26479 18961
rect 26421 18952 26433 18955
rect 26384 18924 26433 18952
rect 26384 18912 26390 18924
rect 26421 18921 26433 18924
rect 26467 18952 26479 18955
rect 26878 18952 26884 18964
rect 26467 18924 26884 18952
rect 26467 18921 26479 18924
rect 26421 18915 26479 18921
rect 26878 18912 26884 18924
rect 26936 18912 26942 18964
rect 37366 18952 37372 18964
rect 37327 18924 37372 18952
rect 37366 18912 37372 18924
rect 37424 18912 37430 18964
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18816 12127 18819
rect 12894 18816 12900 18828
rect 12115 18788 12900 18816
rect 12115 18785 12127 18788
rect 12069 18779 12127 18785
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 34514 18776 34520 18828
rect 34572 18816 34578 18828
rect 34572 18788 37872 18816
rect 34572 18776 34578 18788
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 17126 18748 17132 18760
rect 16623 18720 17132 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 17126 18708 17132 18720
rect 17184 18748 17190 18760
rect 26329 18751 26387 18757
rect 26329 18748 26341 18751
rect 17184 18720 18552 18748
rect 17184 18708 17190 18720
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18680 1918 18692
rect 2501 18683 2559 18689
rect 2501 18680 2513 18683
rect 1912 18652 2513 18680
rect 1912 18640 1918 18652
rect 2501 18649 2513 18652
rect 2547 18649 2559 18683
rect 2501 18643 2559 18649
rect 11793 18683 11851 18689
rect 11793 18649 11805 18683
rect 11839 18680 11851 18683
rect 12434 18680 12440 18692
rect 11839 18652 12440 18680
rect 11839 18649 11851 18652
rect 11793 18643 11851 18649
rect 12434 18640 12440 18652
rect 12492 18640 12498 18692
rect 16850 18689 16856 18692
rect 16844 18643 16856 18689
rect 16908 18680 16914 18692
rect 16908 18652 16944 18680
rect 16850 18640 16856 18643
rect 16908 18640 16914 18652
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 11882 18572 11888 18624
rect 11940 18612 11946 18624
rect 17954 18612 17960 18624
rect 11940 18584 11985 18612
rect 17915 18584 17960 18612
rect 11940 18572 11946 18584
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18524 18621 18552 18720
rect 25608 18720 26341 18748
rect 25608 18624 25636 18720
rect 26329 18717 26341 18720
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 36725 18751 36783 18757
rect 36725 18717 36737 18751
rect 36771 18748 36783 18751
rect 37182 18748 37188 18760
rect 36771 18720 37188 18748
rect 36771 18717 36783 18720
rect 36725 18711 36783 18717
rect 37182 18708 37188 18720
rect 37240 18708 37246 18760
rect 37844 18757 37872 18788
rect 37829 18751 37887 18757
rect 37829 18717 37841 18751
rect 37875 18717 37887 18751
rect 37829 18711 37887 18717
rect 25774 18640 25780 18692
rect 25832 18680 25838 18692
rect 26142 18680 26148 18692
rect 25832 18652 26148 18680
rect 25832 18640 25838 18652
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 18509 18615 18567 18621
rect 18509 18581 18521 18615
rect 18555 18612 18567 18615
rect 24302 18612 24308 18624
rect 18555 18584 24308 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 24302 18572 24308 18584
rect 24360 18572 24366 18624
rect 25590 18612 25596 18624
rect 25551 18584 25596 18612
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 38010 18612 38016 18624
rect 37971 18584 38016 18612
rect 38010 18572 38016 18584
rect 38068 18572 38074 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1486 18408 1492 18420
rect 1447 18380 1492 18408
rect 1486 18368 1492 18380
rect 1544 18368 1550 18420
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 32309 18411 32367 18417
rect 2004 18380 29868 18408
rect 2004 18368 2010 18380
rect 3421 18343 3479 18349
rect 3421 18340 3433 18343
rect 1688 18312 3433 18340
rect 1688 18281 1716 18312
rect 3421 18309 3433 18312
rect 3467 18340 3479 18343
rect 3467 18312 26234 18340
rect 3467 18309 3479 18312
rect 3421 18303 3479 18309
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 2130 18272 2136 18284
rect 2091 18244 2136 18272
rect 1673 18235 1731 18241
rect 2130 18232 2136 18244
rect 2188 18272 2194 18284
rect 2777 18275 2835 18281
rect 2777 18272 2789 18275
rect 2188 18244 2789 18272
rect 2188 18232 2194 18244
rect 2777 18241 2789 18244
rect 2823 18241 2835 18275
rect 16666 18272 16672 18284
rect 16627 18244 16672 18272
rect 2777 18235 2835 18241
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21140 18244 22017 18272
rect 21140 18232 21146 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 21821 18207 21879 18213
rect 21821 18204 21833 18207
rect 12492 18176 21833 18204
rect 12492 18164 12498 18176
rect 21821 18173 21833 18176
rect 21867 18173 21879 18207
rect 26206 18204 26234 18312
rect 27614 18232 27620 18284
rect 27672 18272 27678 18284
rect 28445 18275 28503 18281
rect 28445 18272 28457 18275
rect 27672 18244 28457 18272
rect 27672 18232 27678 18244
rect 28445 18241 28457 18244
rect 28491 18272 28503 18275
rect 28902 18272 28908 18284
rect 28491 18244 28908 18272
rect 28491 18241 28503 18244
rect 28445 18235 28503 18241
rect 28902 18232 28908 18244
rect 28960 18232 28966 18284
rect 29730 18232 29736 18284
rect 29788 18272 29794 18284
rect 29840 18281 29868 18380
rect 32309 18377 32321 18411
rect 32355 18408 32367 18411
rect 32355 18380 35894 18408
rect 32355 18377 32367 18380
rect 32309 18371 32367 18377
rect 30282 18340 30288 18352
rect 30024 18312 30288 18340
rect 30024 18281 30052 18312
rect 30282 18300 30288 18312
rect 30340 18300 30346 18352
rect 35866 18340 35894 18380
rect 35866 18312 37872 18340
rect 29825 18275 29883 18281
rect 29825 18272 29837 18275
rect 29788 18244 29837 18272
rect 29788 18232 29794 18244
rect 29825 18241 29837 18244
rect 29871 18241 29883 18275
rect 29825 18235 29883 18241
rect 30009 18275 30067 18281
rect 30009 18241 30021 18275
rect 30055 18241 30067 18275
rect 30009 18235 30067 18241
rect 30193 18275 30251 18281
rect 30193 18241 30205 18275
rect 30239 18272 30251 18275
rect 32125 18275 32183 18281
rect 32125 18272 32137 18275
rect 30239 18244 32137 18272
rect 30239 18241 30251 18244
rect 30193 18235 30251 18241
rect 32125 18241 32137 18244
rect 32171 18241 32183 18275
rect 32125 18235 32183 18241
rect 34241 18275 34299 18281
rect 34241 18241 34253 18275
rect 34287 18272 34299 18275
rect 35713 18275 35771 18281
rect 35713 18272 35725 18275
rect 34287 18244 35725 18272
rect 34287 18241 34299 18244
rect 34241 18235 34299 18241
rect 35713 18241 35725 18244
rect 35759 18241 35771 18275
rect 35713 18235 35771 18241
rect 35897 18275 35955 18281
rect 35897 18241 35909 18275
rect 35943 18272 35955 18275
rect 36262 18272 36268 18284
rect 35943 18244 36268 18272
rect 35943 18241 35955 18244
rect 35897 18235 35955 18241
rect 36262 18232 36268 18244
rect 36320 18232 36326 18284
rect 37844 18281 37872 18312
rect 37829 18275 37887 18281
rect 37829 18241 37841 18275
rect 37875 18241 37887 18275
rect 37829 18235 37887 18241
rect 34057 18207 34115 18213
rect 34057 18204 34069 18207
rect 26206 18176 34069 18204
rect 21821 18167 21879 18173
rect 34057 18173 34069 18176
rect 34103 18173 34115 18207
rect 34057 18167 34115 18173
rect 36081 18207 36139 18213
rect 36081 18173 36093 18207
rect 36127 18204 36139 18207
rect 37918 18204 37924 18216
rect 36127 18176 37924 18204
rect 36127 18173 36139 18176
rect 36081 18167 36139 18173
rect 37918 18164 37924 18176
rect 37976 18164 37982 18216
rect 2317 18139 2375 18145
rect 2317 18105 2329 18139
rect 2363 18136 2375 18139
rect 11882 18136 11888 18148
rect 2363 18108 11888 18136
rect 2363 18105 2375 18108
rect 2317 18099 2375 18105
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 16850 18136 16856 18148
rect 16811 18108 16856 18136
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 29089 18139 29147 18145
rect 29089 18105 29101 18139
rect 29135 18136 29147 18139
rect 29454 18136 29460 18148
rect 29135 18108 29460 18136
rect 29135 18105 29147 18108
rect 29089 18099 29147 18105
rect 29454 18096 29460 18108
rect 29512 18136 29518 18148
rect 30282 18136 30288 18148
rect 29512 18108 30288 18136
rect 29512 18096 29518 18108
rect 30282 18096 30288 18108
rect 30340 18096 30346 18148
rect 22186 18068 22192 18080
rect 22147 18040 22192 18068
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 38010 18068 38016 18080
rect 37971 18040 38016 18068
rect 38010 18028 38016 18040
rect 38068 18028 38074 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 15712 17836 15761 17864
rect 15712 17824 15718 17836
rect 15749 17833 15761 17836
rect 15795 17833 15807 17867
rect 16666 17864 16672 17876
rect 16627 17836 16672 17864
rect 15749 17827 15807 17833
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 25774 17864 25780 17876
rect 25735 17836 25780 17864
rect 25774 17824 25780 17836
rect 25832 17824 25838 17876
rect 29730 17864 29736 17876
rect 29691 17836 29736 17864
rect 29730 17824 29736 17836
rect 29788 17824 29794 17876
rect 37918 17864 37924 17876
rect 37879 17836 37924 17864
rect 37918 17824 37924 17836
rect 37976 17824 37982 17876
rect 16206 17688 16212 17740
rect 16264 17728 16270 17740
rect 17221 17731 17279 17737
rect 17221 17728 17233 17731
rect 16264 17700 17233 17728
rect 16264 17688 16270 17700
rect 17221 17697 17233 17700
rect 17267 17697 17279 17731
rect 17221 17691 17279 17697
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 18012 17700 20913 17728
rect 18012 17688 18018 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 22186 17688 22192 17740
rect 22244 17728 22250 17740
rect 22649 17731 22707 17737
rect 22649 17728 22661 17731
rect 22244 17700 22661 17728
rect 22244 17688 22250 17700
rect 22649 17697 22661 17700
rect 22695 17697 22707 17731
rect 22649 17691 22707 17697
rect 22925 17731 22983 17737
rect 22925 17697 22937 17731
rect 22971 17728 22983 17731
rect 22971 17700 24532 17728
rect 22971 17697 22983 17700
rect 22925 17691 22983 17697
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 17037 17663 17095 17669
rect 1719 17632 3924 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2222 17524 2228 17536
rect 2183 17496 2228 17524
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 2777 17527 2835 17533
rect 2777 17493 2789 17527
rect 2823 17524 2835 17527
rect 2866 17524 2872 17536
rect 2823 17496 2872 17524
rect 2823 17493 2835 17496
rect 2777 17487 2835 17493
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 3896 17533 3924 17632
rect 17037 17629 17049 17663
rect 17083 17660 17095 17663
rect 17972 17660 18000 17688
rect 21082 17660 21088 17672
rect 17083 17632 18000 17660
rect 21043 17632 21088 17660
rect 17083 17629 17095 17632
rect 17037 17623 17095 17629
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 24302 17620 24308 17672
rect 24360 17660 24366 17672
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 24360 17632 24409 17660
rect 24360 17620 24366 17632
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 24504 17660 24532 17700
rect 36814 17660 36820 17672
rect 24504 17632 36820 17660
rect 24397 17623 24455 17629
rect 36814 17620 36820 17632
rect 36872 17620 36878 17672
rect 37461 17663 37519 17669
rect 37461 17629 37473 17663
rect 37507 17660 37519 17663
rect 38102 17660 38108 17672
rect 37507 17632 38108 17660
rect 37507 17629 37519 17632
rect 37461 17623 37519 17629
rect 38102 17620 38108 17632
rect 38160 17620 38166 17672
rect 14458 17592 14464 17604
rect 14419 17564 14464 17592
rect 14458 17552 14464 17564
rect 14516 17552 14522 17604
rect 24118 17552 24124 17604
rect 24176 17592 24182 17604
rect 24642 17595 24700 17601
rect 24642 17592 24654 17595
rect 24176 17564 24654 17592
rect 24176 17552 24182 17564
rect 24642 17561 24654 17564
rect 24688 17561 24700 17595
rect 24642 17555 24700 17561
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17524 3939 17527
rect 11698 17524 11704 17536
rect 3927 17496 11704 17524
rect 3927 17493 3939 17496
rect 3881 17487 3939 17493
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 21269 17527 21327 17533
rect 17184 17496 17229 17524
rect 17184 17484 17190 17496
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 22554 17524 22560 17536
rect 21315 17496 22560 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8018 17320 8024 17332
rect 1964 17292 7420 17320
rect 7979 17292 8024 17320
rect 1964 17193 1992 17292
rect 4062 17252 4068 17264
rect 2792 17224 4068 17252
rect 2792 17193 2820 17224
rect 4062 17212 4068 17224
rect 4120 17252 4126 17264
rect 4801 17255 4859 17261
rect 4801 17252 4813 17255
rect 4120 17224 4813 17252
rect 4120 17212 4126 17224
rect 4801 17221 4813 17224
rect 4847 17252 4859 17255
rect 6914 17252 6920 17264
rect 4847 17224 6920 17252
rect 4847 17221 4859 17224
rect 4801 17215 4859 17221
rect 6914 17212 6920 17224
rect 6972 17212 6978 17264
rect 7392 17252 7420 17292
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 24302 17320 24308 17332
rect 11756 17292 18184 17320
rect 24263 17292 24308 17320
rect 11756 17280 11762 17292
rect 17126 17252 17132 17264
rect 7392 17224 17132 17252
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 18156 17252 18184 17292
rect 24302 17280 24308 17292
rect 24360 17280 24366 17332
rect 34333 17255 34391 17261
rect 34333 17252 34345 17255
rect 18156 17224 34345 17252
rect 34333 17221 34345 17224
rect 34379 17221 34391 17255
rect 34333 17215 34391 17221
rect 3050 17193 3056 17196
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17153 2007 17187
rect 1949 17147 2007 17153
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 3044 17147 3056 17193
rect 3108 17184 3114 17196
rect 3108 17156 3144 17184
rect 3050 17144 3056 17147
rect 3108 17144 3114 17156
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 8076 17156 12817 17184
rect 8076 17144 8082 17156
rect 12805 17153 12817 17156
rect 12851 17184 12863 17187
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 12851 17156 13553 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 29178 17144 29184 17196
rect 29236 17184 29242 17196
rect 29454 17184 29460 17196
rect 29236 17156 29460 17184
rect 29236 17144 29242 17156
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 34517 17187 34575 17193
rect 34517 17153 34529 17187
rect 34563 17184 34575 17187
rect 36078 17184 36084 17196
rect 34563 17156 36084 17184
rect 34563 17153 34575 17156
rect 34517 17147 34575 17153
rect 36078 17144 36084 17156
rect 36136 17144 36142 17196
rect 36814 17144 36820 17196
rect 36872 17184 36878 17196
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 36872 17156 37841 17184
rect 36872 17144 36878 17156
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 2222 17116 2228 17128
rect 2183 17088 2228 17116
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 29273 17119 29331 17125
rect 29273 17116 29285 17119
rect 28736 17088 29285 17116
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 5074 16980 5080 16992
rect 4203 16952 5080 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 12952 16952 13001 16980
rect 12952 16940 12958 16952
rect 12989 16949 13001 16952
rect 13035 16949 13047 16983
rect 12989 16943 13047 16949
rect 14369 16983 14427 16989
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 14458 16980 14464 16992
rect 14415 16952 14464 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 14458 16940 14464 16952
rect 14516 16940 14522 16992
rect 21358 16940 21364 16992
rect 21416 16980 21422 16992
rect 28736 16989 28764 17088
rect 29273 17085 29285 17088
rect 29319 17085 29331 17119
rect 29273 17079 29331 17085
rect 28721 16983 28779 16989
rect 28721 16980 28733 16983
rect 21416 16952 28733 16980
rect 21416 16940 21422 16952
rect 28721 16949 28733 16952
rect 28767 16949 28779 16983
rect 29638 16980 29644 16992
rect 29599 16952 29644 16980
rect 28721 16943 28779 16949
rect 29638 16940 29644 16952
rect 29696 16940 29702 16992
rect 37366 16980 37372 16992
rect 37327 16952 37372 16980
rect 37366 16940 37372 16952
rect 37424 16940 37430 16992
rect 38010 16980 38016 16992
rect 37971 16952 38016 16980
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 21358 16776 21364 16788
rect 1995 16748 21364 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 36078 16776 36084 16788
rect 36039 16748 36084 16776
rect 36078 16736 36084 16748
rect 36136 16736 36142 16788
rect 37826 16776 37832 16788
rect 36372 16748 37832 16776
rect 4614 16708 4620 16720
rect 4264 16680 4620 16708
rect 4264 16649 4292 16680
rect 4614 16668 4620 16680
rect 4672 16668 4678 16720
rect 36372 16708 36400 16748
rect 37826 16736 37832 16748
rect 37884 16736 37890 16788
rect 37185 16711 37243 16717
rect 37185 16708 37197 16711
rect 26206 16680 36400 16708
rect 36464 16680 37197 16708
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 7466 16640 7472 16652
rect 4479 16612 7472 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 7466 16600 7472 16612
rect 7524 16600 7530 16652
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 16206 16640 16212 16652
rect 12952 16612 16212 16640
rect 12952 16600 12958 16612
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 22554 16640 22560 16652
rect 22515 16612 22560 16640
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 22833 16643 22891 16649
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 26206 16640 26234 16680
rect 36464 16649 36492 16680
rect 37185 16677 37197 16680
rect 37231 16677 37243 16711
rect 37185 16671 37243 16677
rect 22879 16612 26234 16640
rect 36449 16643 36507 16649
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 36449 16609 36461 16643
rect 36495 16609 36507 16643
rect 36449 16603 36507 16609
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16572 2835 16575
rect 4522 16572 4528 16584
rect 2823 16544 4528 16572
rect 2823 16541 2835 16544
rect 2777 16535 2835 16541
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8018 16572 8024 16584
rect 7975 16544 8024 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 29638 16532 29644 16584
rect 29696 16572 29702 16584
rect 30745 16575 30803 16581
rect 30745 16572 30757 16575
rect 29696 16544 30757 16572
rect 29696 16532 29702 16544
rect 30745 16541 30757 16544
rect 30791 16541 30803 16575
rect 36262 16572 36268 16584
rect 36223 16544 36268 16572
rect 30745 16535 30803 16541
rect 36262 16532 36268 16544
rect 36320 16532 36326 16584
rect 37366 16572 37372 16584
rect 37327 16544 37372 16572
rect 37366 16532 37372 16544
rect 37424 16532 37430 16584
rect 37829 16575 37887 16581
rect 37829 16541 37841 16575
rect 37875 16541 37887 16575
rect 37829 16535 37887 16541
rect 1857 16507 1915 16513
rect 1857 16473 1869 16507
rect 1903 16504 1915 16507
rect 2866 16504 2872 16516
rect 1903 16476 2872 16504
rect 1903 16473 1915 16476
rect 1857 16467 1915 16473
rect 2866 16464 2872 16476
rect 2924 16464 2930 16516
rect 37844 16504 37872 16535
rect 30944 16476 37872 16504
rect 2593 16439 2651 16445
rect 2593 16405 2605 16439
rect 2639 16436 2651 16439
rect 2774 16436 2780 16448
rect 2639 16408 2780 16436
rect 2639 16405 2651 16408
rect 2593 16399 2651 16405
rect 2774 16396 2780 16408
rect 2832 16396 2838 16448
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16436 4215 16439
rect 5074 16436 5080 16448
rect 4203 16408 5080 16436
rect 4203 16405 4215 16408
rect 4157 16399 4215 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 7466 16396 7472 16448
rect 7524 16436 7530 16448
rect 30944 16445 30972 16476
rect 7745 16439 7803 16445
rect 7745 16436 7757 16439
rect 7524 16408 7757 16436
rect 7524 16396 7530 16408
rect 7745 16405 7757 16408
rect 7791 16405 7803 16439
rect 7745 16399 7803 16405
rect 30929 16439 30987 16445
rect 30929 16405 30941 16439
rect 30975 16405 30987 16439
rect 38010 16436 38016 16448
rect 37971 16408 38016 16436
rect 30929 16399 30987 16405
rect 38010 16396 38016 16408
rect 38068 16396 38074 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 3050 16232 3056 16244
rect 3007 16204 3056 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 8018 16124 8024 16176
rect 8076 16164 8082 16176
rect 8205 16167 8263 16173
rect 8205 16164 8217 16167
rect 8076 16136 8217 16164
rect 8076 16124 8082 16136
rect 8205 16133 8217 16136
rect 8251 16164 8263 16167
rect 8757 16167 8815 16173
rect 8757 16164 8769 16167
rect 8251 16136 8769 16164
rect 8251 16133 8263 16136
rect 8205 16127 8263 16133
rect 8757 16133 8769 16136
rect 8803 16133 8815 16167
rect 8757 16127 8815 16133
rect 36262 16124 36268 16176
rect 36320 16164 36326 16176
rect 36320 16136 37504 16164
rect 36320 16124 36326 16136
rect 1854 16096 1860 16108
rect 1815 16068 1860 16096
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 3145 16099 3203 16105
rect 3145 16065 3157 16099
rect 3191 16096 3203 16099
rect 3786 16096 3792 16108
rect 3191 16068 3792 16096
rect 3191 16065 3203 16068
rect 3145 16059 3203 16065
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 29178 16096 29184 16108
rect 29139 16068 29184 16096
rect 29178 16056 29184 16068
rect 29236 16056 29242 16108
rect 37476 16105 37504 16136
rect 29365 16099 29423 16105
rect 29365 16065 29377 16099
rect 29411 16096 29423 16099
rect 30377 16099 30435 16105
rect 30377 16096 30389 16099
rect 29411 16068 30389 16096
rect 29411 16065 29423 16068
rect 29365 16059 29423 16065
rect 30377 16065 30389 16068
rect 30423 16065 30435 16099
rect 30377 16059 30435 16065
rect 36357 16099 36415 16105
rect 36357 16065 36369 16099
rect 36403 16096 36415 16099
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 36403 16068 37289 16096
rect 36403 16065 36415 16068
rect 36357 16059 36415 16065
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37277 16059 37335 16065
rect 37461 16099 37519 16105
rect 37461 16065 37473 16099
rect 37507 16065 37519 16099
rect 37461 16059 37519 16065
rect 1872 16028 1900 16056
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 1872 16000 3617 16028
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 28997 16031 29055 16037
rect 28997 15997 29009 16031
rect 29043 15997 29055 16031
rect 28997 15991 29055 15997
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15960 2099 15963
rect 28445 15963 28503 15969
rect 28445 15960 28457 15963
rect 2087 15932 28457 15960
rect 2087 15929 2099 15932
rect 2041 15923 2099 15929
rect 28445 15929 28457 15932
rect 28491 15960 28503 15963
rect 29012 15960 29040 15991
rect 36078 15988 36084 16040
rect 36136 16028 36142 16040
rect 37645 16031 37703 16037
rect 37645 16028 37657 16031
rect 36136 16000 37657 16028
rect 36136 15988 36142 16000
rect 37645 15997 37657 16000
rect 37691 15997 37703 16031
rect 37645 15991 37703 15997
rect 28491 15932 29040 15960
rect 28491 15929 28503 15932
rect 28445 15923 28503 15929
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 4614 15892 4620 15904
rect 4295 15864 4620 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 7926 15892 7932 15904
rect 7887 15864 7932 15892
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 30558 15892 30564 15904
rect 30519 15864 30564 15892
rect 30558 15852 30564 15864
rect 30616 15852 30622 15904
rect 36170 15892 36176 15904
rect 36131 15864 36176 15892
rect 36170 15852 36176 15864
rect 36228 15852 36234 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 36170 15688 36176 15700
rect 4672 15660 36176 15688
rect 4672 15648 4678 15660
rect 36170 15648 36176 15660
rect 36228 15648 36234 15700
rect 38010 15688 38016 15700
rect 37971 15660 38016 15688
rect 38010 15648 38016 15660
rect 38068 15648 38074 15700
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 16206 15552 16212 15564
rect 6972 15524 7017 15552
rect 16167 15524 16212 15552
rect 6972 15512 6978 15524
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15453 2007 15487
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 1949 15447 2007 15453
rect 1964 15416 1992 15447
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3878 15484 3884 15496
rect 3007 15456 3884 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 6932 15484 6960 15512
rect 8938 15484 8944 15496
rect 6932 15456 8944 15484
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 11698 15484 11704 15496
rect 11659 15456 11704 15484
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 30558 15444 30564 15496
rect 30616 15484 30622 15496
rect 37093 15487 37151 15493
rect 37093 15484 37105 15487
rect 30616 15456 37105 15484
rect 30616 15444 30622 15456
rect 37093 15453 37105 15456
rect 37139 15453 37151 15487
rect 37826 15484 37832 15496
rect 37787 15456 37832 15484
rect 37093 15447 37151 15453
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 7184 15419 7242 15425
rect 1964 15388 6914 15416
rect 2774 15348 2780 15360
rect 2735 15320 2780 15348
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 3878 15348 3884 15360
rect 3839 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 6886 15348 6914 15388
rect 7184 15385 7196 15419
rect 7230 15416 7242 15419
rect 7282 15416 7288 15428
rect 7230 15388 7288 15416
rect 7230 15385 7242 15388
rect 7184 15379 7242 15385
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 16393 15419 16451 15425
rect 16393 15416 16405 15419
rect 7392 15388 16405 15416
rect 7392 15348 7420 15388
rect 16393 15385 16405 15388
rect 16439 15385 16451 15419
rect 16393 15379 16451 15385
rect 16485 15419 16543 15425
rect 16485 15385 16497 15419
rect 16531 15416 16543 15419
rect 19242 15416 19248 15428
rect 16531 15388 19248 15416
rect 16531 15385 16543 15388
rect 16485 15379 16543 15385
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 8294 15348 8300 15360
rect 6886 15320 7420 15348
rect 8255 15320 8300 15348
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 11885 15351 11943 15357
rect 11885 15317 11897 15351
rect 11931 15348 11943 15351
rect 11974 15348 11980 15360
rect 11931 15320 11980 15348
rect 11931 15317 11943 15320
rect 11885 15311 11943 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 16853 15351 16911 15357
rect 16853 15317 16865 15351
rect 16899 15348 16911 15351
rect 17310 15348 17316 15360
rect 16899 15320 17316 15348
rect 16899 15317 16911 15320
rect 16853 15311 16911 15317
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 36262 15348 36268 15360
rect 36223 15320 36268 15348
rect 36262 15308 36268 15320
rect 36320 15308 36326 15360
rect 37274 15348 37280 15360
rect 37235 15320 37280 15348
rect 37274 15308 37280 15320
rect 37332 15308 37338 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 2501 15147 2559 15153
rect 2501 15144 2513 15147
rect 2280 15116 2513 15144
rect 2280 15104 2286 15116
rect 2501 15113 2513 15116
rect 2547 15113 2559 15147
rect 7282 15144 7288 15156
rect 7243 15116 7288 15144
rect 2501 15107 2559 15113
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 8996 15116 10885 15144
rect 8996 15104 9002 15116
rect 10873 15113 10885 15116
rect 10919 15144 10931 15147
rect 17497 15147 17555 15153
rect 10919 15116 11744 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 3878 15036 3884 15088
rect 3936 15076 3942 15088
rect 3936 15048 10824 15076
rect 3936 15036 3942 15048
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 15008 1918 15020
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 1912 14980 3065 15008
rect 1912 14968 1918 14980
rect 3053 14977 3065 14980
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 6972 14980 7113 15008
rect 6972 14968 6978 14980
rect 7101 14977 7113 14980
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 10796 14940 10824 15048
rect 11716 15017 11744 15116
rect 16546 15116 17448 15144
rect 16546 15076 16574 15116
rect 11808 15048 16574 15076
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11808 14940 11836 15048
rect 11974 15017 11980 15020
rect 11968 15008 11980 15017
rect 11935 14980 11980 15008
rect 11968 14971 11980 14980
rect 11974 14968 11980 14971
rect 12032 14968 12038 15020
rect 17310 15008 17316 15020
rect 17271 14980 17316 15008
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 17420 15008 17448 15116
rect 17497 15113 17509 15147
rect 17543 15113 17555 15147
rect 24946 15144 24952 15156
rect 24907 15116 24952 15144
rect 17497 15107 17555 15113
rect 17512 15076 17540 15107
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 36078 15144 36084 15156
rect 36039 15116 36084 15144
rect 36078 15104 36084 15116
rect 36136 15104 36142 15156
rect 18662 15079 18720 15085
rect 18662 15076 18674 15079
rect 17512 15048 18674 15076
rect 18662 15045 18674 15048
rect 18708 15045 18720 15079
rect 18662 15039 18720 15045
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 17420 14980 23489 15008
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 23658 15008 23664 15020
rect 23619 14980 23664 15008
rect 23477 14971 23535 14977
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 24305 15011 24363 15017
rect 24305 14977 24317 15011
rect 24351 15008 24363 15011
rect 24964 15008 24992 15104
rect 24351 14980 24992 15008
rect 24351 14977 24363 14980
rect 24305 14971 24363 14977
rect 33226 14968 33232 15020
rect 33284 15008 33290 15020
rect 33321 15011 33379 15017
rect 33321 15008 33333 15011
rect 33284 14980 33333 15008
rect 33284 14968 33290 14980
rect 33321 14977 33333 14980
rect 33367 14977 33379 15011
rect 33321 14971 33379 14977
rect 35897 15011 35955 15017
rect 35897 14977 35909 15011
rect 35943 15008 35955 15011
rect 36262 15008 36268 15020
rect 35943 14980 36268 15008
rect 35943 14977 35955 14980
rect 35897 14971 35955 14977
rect 36262 14968 36268 14980
rect 36320 14968 36326 15020
rect 36541 15011 36599 15017
rect 36541 14977 36553 15011
rect 36587 14977 36599 15011
rect 37829 15011 37887 15017
rect 37829 15008 37841 15011
rect 36541 14971 36599 14977
rect 36740 14980 37841 15008
rect 10796 14912 11836 14940
rect 18417 14943 18475 14949
rect 18417 14909 18429 14943
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 13078 14804 13084 14816
rect 13039 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 18432 14804 18460 14903
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 33137 14943 33195 14949
rect 33137 14940 33149 14943
rect 19484 14912 33149 14940
rect 19484 14900 19490 14912
rect 19812 14881 19840 14912
rect 33137 14909 33149 14912
rect 33183 14909 33195 14943
rect 33137 14903 33195 14909
rect 33505 14943 33563 14949
rect 33505 14909 33517 14943
rect 33551 14940 33563 14943
rect 36556 14940 36584 14971
rect 33551 14912 36584 14940
rect 33551 14909 33563 14912
rect 33505 14903 33563 14909
rect 19797 14875 19855 14881
rect 19797 14841 19809 14875
rect 19843 14841 19855 14875
rect 19797 14835 19855 14841
rect 24762 14832 24768 14884
rect 24820 14872 24826 14884
rect 36630 14872 36636 14884
rect 24820 14844 36636 14872
rect 24820 14832 24826 14844
rect 36630 14832 36636 14844
rect 36688 14832 36694 14884
rect 36740 14881 36768 14980
rect 37829 14977 37841 14980
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 36725 14875 36783 14881
rect 36725 14841 36737 14875
rect 36771 14841 36783 14875
rect 36725 14835 36783 14841
rect 19334 14804 19340 14816
rect 18432 14776 19340 14804
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 24302 14764 24308 14816
rect 24360 14804 24366 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 24360 14776 24501 14804
rect 24360 14764 24366 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 38010 14804 38016 14816
rect 37971 14776 38016 14804
rect 24489 14767 24547 14773
rect 38010 14764 38016 14776
rect 38068 14764 38074 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 21358 14600 21364 14612
rect 2004 14572 21364 14600
rect 2004 14560 2010 14572
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 23658 14560 23664 14612
rect 23716 14600 23722 14612
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 23716 14572 24409 14600
rect 23716 14560 23722 14572
rect 24397 14569 24409 14572
rect 24443 14569 24455 14603
rect 24397 14563 24455 14569
rect 26142 14560 26148 14612
rect 26200 14600 26206 14612
rect 26513 14603 26571 14609
rect 26513 14600 26525 14603
rect 26200 14572 26525 14600
rect 26200 14560 26206 14572
rect 26513 14569 26525 14572
rect 26559 14569 26571 14603
rect 26513 14563 26571 14569
rect 36630 14560 36636 14612
rect 36688 14600 36694 14612
rect 37185 14603 37243 14609
rect 37185 14600 37197 14603
rect 36688 14572 37197 14600
rect 36688 14560 36694 14572
rect 37185 14569 37197 14572
rect 37231 14569 37243 14603
rect 37185 14563 37243 14569
rect 5074 14492 5080 14544
rect 5132 14532 5138 14544
rect 32585 14535 32643 14541
rect 32585 14532 32597 14535
rect 5132 14504 32597 14532
rect 5132 14492 5138 14504
rect 32585 14501 32597 14504
rect 32631 14532 32643 14535
rect 32631 14504 33180 14532
rect 32631 14501 32643 14504
rect 32585 14495 32643 14501
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14464 12403 14467
rect 12894 14464 12900 14476
rect 12391 14436 12900 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 13078 14464 13084 14476
rect 13035 14436 13084 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14396 1458 14408
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1452 14368 2053 14396
rect 1452 14356 1458 14368
rect 2041 14365 2053 14368
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 13004 14396 13032 14427
rect 13078 14424 13084 14436
rect 13136 14464 13142 14476
rect 32490 14464 32496 14476
rect 13136 14436 32496 14464
rect 13136 14424 13142 14436
rect 32490 14424 32496 14436
rect 32548 14424 32554 14476
rect 33152 14473 33180 14504
rect 33137 14467 33195 14473
rect 33137 14433 33149 14467
rect 33183 14433 33195 14467
rect 33137 14427 33195 14433
rect 12115 14368 13032 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 24302 14356 24308 14408
rect 24360 14396 24366 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24360 14368 24593 14396
rect 24360 14356 24366 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24762 14396 24768 14408
rect 24723 14368 24768 14396
rect 24581 14359 24639 14365
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 24854 14356 24860 14408
rect 24912 14396 24918 14408
rect 26142 14396 26148 14408
rect 24912 14368 26148 14396
rect 24912 14356 24918 14368
rect 26142 14356 26148 14368
rect 26200 14396 26206 14408
rect 27065 14399 27123 14405
rect 27065 14396 27077 14399
rect 26200 14368 27077 14396
rect 26200 14356 26206 14368
rect 27065 14365 27077 14368
rect 27111 14365 27123 14399
rect 27065 14359 27123 14365
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28537 14399 28595 14405
rect 28537 14365 28549 14399
rect 28583 14396 28595 14399
rect 29641 14399 29699 14405
rect 29641 14396 29653 14399
rect 28583 14368 29653 14396
rect 28583 14365 28595 14368
rect 28537 14359 28595 14365
rect 29641 14365 29653 14368
rect 29687 14365 29699 14399
rect 29641 14359 29699 14365
rect 12161 14331 12219 14337
rect 12161 14328 12173 14331
rect 1596 14300 12173 14328
rect 1596 14269 1624 14300
rect 12161 14297 12173 14300
rect 12207 14297 12219 14331
rect 12161 14291 12219 14297
rect 21358 14288 21364 14340
rect 21416 14328 21422 14340
rect 27982 14328 27988 14340
rect 21416 14300 27988 14328
rect 21416 14288 21422 14300
rect 27982 14288 27988 14300
rect 28040 14328 28046 14340
rect 28184 14328 28212 14359
rect 28040 14300 28212 14328
rect 28040 14288 28046 14300
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14229 1639 14263
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 1581 14223 1639 14229
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 11698 14260 11704 14272
rect 11659 14232 11704 14260
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 18325 14263 18383 14269
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 19334 14260 19340 14272
rect 18371 14232 19340 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 27249 14263 27307 14269
rect 27249 14229 27261 14263
rect 27295 14260 27307 14263
rect 28368 14260 28396 14359
rect 33226 14356 33232 14408
rect 33284 14396 33290 14408
rect 33321 14399 33379 14405
rect 33321 14396 33333 14399
rect 33284 14368 33333 14396
rect 33284 14356 33290 14368
rect 33321 14365 33333 14368
rect 33367 14365 33379 14399
rect 33321 14359 33379 14365
rect 36725 14399 36783 14405
rect 36725 14365 36737 14399
rect 36771 14396 36783 14399
rect 37182 14396 37188 14408
rect 36771 14368 37188 14396
rect 36771 14365 36783 14368
rect 36725 14359 36783 14365
rect 37182 14356 37188 14368
rect 37240 14396 37246 14408
rect 37369 14399 37427 14405
rect 37369 14396 37381 14399
rect 37240 14368 37381 14396
rect 37240 14356 37246 14368
rect 37369 14365 37381 14368
rect 37415 14365 37427 14399
rect 37369 14359 37427 14365
rect 37829 14399 37887 14405
rect 37829 14365 37841 14399
rect 37875 14365 37887 14399
rect 37829 14359 37887 14365
rect 37844 14328 37872 14359
rect 29840 14300 37872 14328
rect 28442 14260 28448 14272
rect 27295 14232 28448 14260
rect 27295 14229 27307 14232
rect 27249 14223 27307 14229
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 29840 14269 29868 14300
rect 29825 14263 29883 14269
rect 29825 14229 29837 14263
rect 29871 14229 29883 14263
rect 29825 14223 29883 14229
rect 33505 14263 33563 14269
rect 33505 14229 33517 14263
rect 33551 14260 33563 14263
rect 36262 14260 36268 14272
rect 33551 14232 36268 14260
rect 33551 14229 33563 14232
rect 33505 14223 33563 14229
rect 36262 14220 36268 14232
rect 36320 14220 36326 14272
rect 38010 14260 38016 14272
rect 37971 14232 38016 14260
rect 38010 14220 38016 14232
rect 38068 14220 38074 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 24305 14059 24363 14065
rect 24305 14056 24317 14059
rect 6972 14028 7017 14056
rect 16546 14028 24317 14056
rect 6972 14016 6978 14028
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 16546 13988 16574 14028
rect 24305 14025 24317 14028
rect 24351 14025 24363 14059
rect 27982 14056 27988 14068
rect 27943 14028 27988 14056
rect 24305 14019 24363 14025
rect 27982 14016 27988 14028
rect 28040 14016 28046 14068
rect 32490 14056 32496 14068
rect 32451 14028 32496 14056
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 34514 14016 34520 14068
rect 34572 14056 34578 14068
rect 37921 14059 37979 14065
rect 37921 14056 37933 14059
rect 34572 14028 37933 14056
rect 34572 14016 34578 14028
rect 37921 14025 37933 14028
rect 37967 14025 37979 14059
rect 37921 14019 37979 14025
rect 2740 13960 16574 13988
rect 23017 13991 23075 13997
rect 2740 13948 2746 13960
rect 23017 13957 23029 13991
rect 23063 13988 23075 13991
rect 24946 13988 24952 14000
rect 23063 13960 24952 13988
rect 23063 13957 23075 13960
rect 23017 13951 23075 13957
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13920 1918 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 1912 13892 3065 13920
rect 1912 13880 1918 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13920 7343 13923
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 7331 13892 8248 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 7374 13852 7380 13864
rect 7335 13824 7380 13852
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 8220 13861 8248 13892
rect 21376 13892 22017 13920
rect 21376 13864 21404 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13889 22339 13923
rect 22281 13883 22339 13889
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13920 22523 13923
rect 23032 13920 23060 13951
rect 24946 13948 24952 13960
rect 25004 13948 25010 14000
rect 24394 13920 24400 13932
rect 22511 13892 23060 13920
rect 24355 13892 24400 13920
rect 22511 13889 22523 13892
rect 22465 13883 22523 13889
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13852 8263 13855
rect 8294 13852 8300 13864
rect 8251 13824 8300 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 2038 13784 2044 13796
rect 1999 13756 2044 13784
rect 2038 13744 2044 13756
rect 2096 13744 2102 13796
rect 7466 13744 7472 13796
rect 7524 13784 7530 13796
rect 7576 13784 7604 13815
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21358 13852 21364 13864
rect 21315 13824 21364 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 21818 13852 21824 13864
rect 21779 13824 21824 13852
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22296 13852 22324 13883
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 32508 13920 32536 14016
rect 33045 13923 33103 13929
rect 33045 13920 33057 13923
rect 32508 13892 33057 13920
rect 33045 13889 33057 13892
rect 33091 13889 33103 13923
rect 33045 13883 33103 13889
rect 33134 13880 33140 13932
rect 33192 13920 33198 13932
rect 33229 13923 33287 13929
rect 33229 13920 33241 13923
rect 33192 13892 33241 13920
rect 33192 13880 33198 13892
rect 33229 13889 33241 13892
rect 33275 13889 33287 13923
rect 33229 13883 33287 13889
rect 33413 13923 33471 13929
rect 33413 13889 33425 13923
rect 33459 13920 33471 13923
rect 37277 13923 37335 13929
rect 37277 13920 37289 13923
rect 33459 13892 37289 13920
rect 33459 13889 33471 13892
rect 33413 13883 33471 13889
rect 37277 13889 37289 13892
rect 37323 13889 37335 13923
rect 38102 13920 38108 13932
rect 38063 13892 38108 13920
rect 37277 13883 37335 13889
rect 38102 13880 38108 13892
rect 38160 13880 38166 13932
rect 23477 13855 23535 13861
rect 23477 13852 23489 13855
rect 22296 13824 23489 13852
rect 23477 13821 23489 13824
rect 23523 13852 23535 13855
rect 24854 13852 24860 13864
rect 23523 13824 24860 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 36725 13855 36783 13861
rect 36725 13821 36737 13855
rect 36771 13852 36783 13855
rect 38120 13852 38148 13880
rect 36771 13824 38148 13852
rect 36771 13821 36783 13824
rect 36725 13815 36783 13821
rect 7524 13756 7604 13784
rect 7524 13744 7530 13756
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 2501 13719 2559 13725
rect 2501 13716 2513 13719
rect 2004 13688 2513 13716
rect 2004 13676 2010 13688
rect 2501 13685 2513 13688
rect 2547 13685 2559 13719
rect 2501 13679 2559 13685
rect 37461 13719 37519 13725
rect 37461 13685 37473 13719
rect 37507 13716 37519 13719
rect 37826 13716 37832 13728
rect 37507 13688 37832 13716
rect 37507 13685 37519 13688
rect 37461 13679 37519 13685
rect 37826 13676 37832 13688
rect 37884 13676 37890 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1486 13512 1492 13524
rect 1447 13484 1492 13512
rect 1486 13472 1492 13484
rect 1544 13472 1550 13524
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 4706 13512 4712 13524
rect 2363 13484 4712 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 24857 13515 24915 13521
rect 24857 13512 24869 13515
rect 24452 13484 24869 13512
rect 24452 13472 24458 13484
rect 24857 13481 24869 13484
rect 24903 13481 24915 13515
rect 24857 13475 24915 13481
rect 2682 13376 2688 13388
rect 1688 13348 2688 13376
rect 1688 13317 1716 13348
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 25225 13379 25283 13385
rect 25225 13345 25237 13379
rect 25271 13376 25283 13379
rect 34514 13376 34520 13388
rect 25271 13348 34520 13376
rect 25271 13345 25283 13348
rect 25225 13339 25283 13345
rect 34514 13336 34520 13348
rect 34572 13336 34578 13388
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 2130 13308 2136 13320
rect 2091 13280 2136 13308
rect 1673 13271 1731 13277
rect 2130 13268 2136 13280
rect 2188 13308 2194 13320
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2188 13280 2789 13308
rect 2188 13268 2194 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 24302 13268 24308 13320
rect 24360 13308 24366 13320
rect 25041 13311 25099 13317
rect 25041 13308 25053 13311
rect 24360 13280 25053 13308
rect 24360 13268 24366 13280
rect 25041 13277 25053 13280
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 28261 13311 28319 13317
rect 28261 13277 28273 13311
rect 28307 13277 28319 13311
rect 28442 13308 28448 13320
rect 28403 13280 28448 13308
rect 28261 13271 28319 13277
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 27709 13243 27767 13249
rect 27709 13240 27721 13243
rect 2096 13212 27721 13240
rect 2096 13200 2102 13212
rect 27709 13209 27721 13212
rect 27755 13240 27767 13243
rect 28276 13240 28304 13271
rect 28442 13268 28448 13280
rect 28500 13268 28506 13320
rect 36078 13308 36084 13320
rect 36039 13280 36084 13308
rect 36078 13268 36084 13280
rect 36136 13268 36142 13320
rect 36262 13268 36268 13320
rect 36320 13308 36326 13320
rect 36725 13311 36783 13317
rect 36725 13308 36737 13311
rect 36320 13280 36737 13308
rect 36320 13268 36326 13280
rect 36725 13277 36737 13280
rect 36771 13277 36783 13311
rect 37826 13308 37832 13320
rect 37787 13280 37832 13308
rect 36725 13271 36783 13277
rect 37826 13268 37832 13280
rect 37884 13268 37890 13320
rect 27755 13212 28304 13240
rect 27755 13209 27767 13212
rect 27709 13203 27767 13209
rect 28626 13172 28632 13184
rect 28587 13144 28632 13172
rect 28626 13132 28632 13144
rect 28684 13132 28690 13184
rect 36262 13172 36268 13184
rect 36223 13144 36268 13172
rect 36262 13132 36268 13144
rect 36320 13132 36326 13184
rect 36909 13175 36967 13181
rect 36909 13141 36921 13175
rect 36955 13172 36967 13175
rect 37826 13172 37832 13184
rect 36955 13144 37832 13172
rect 36955 13141 36967 13144
rect 36909 13135 36967 13141
rect 37826 13132 37832 13144
rect 37884 13132 37890 13184
rect 38010 13172 38016 13184
rect 37971 13144 38016 13172
rect 38010 13132 38016 13144
rect 38068 13132 38074 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4120 12940 4813 12968
rect 4120 12928 4126 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 15105 12971 15163 12977
rect 15105 12937 15117 12971
rect 15151 12968 15163 12971
rect 15378 12968 15384 12980
rect 15151 12940 15384 12968
rect 15151 12937 15163 12940
rect 15105 12931 15163 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 28626 12928 28632 12980
rect 28684 12968 28690 12980
rect 36078 12968 36084 12980
rect 28684 12940 36084 12968
rect 28684 12928 28690 12940
rect 36078 12928 36084 12940
rect 36136 12928 36142 12980
rect 4080 12900 4108 12928
rect 2884 12872 4108 12900
rect 15120 12872 15976 12900
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 2884 12841 2912 12872
rect 3142 12841 3148 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 3136 12795 3148 12841
rect 3200 12832 3206 12844
rect 3200 12804 3236 12832
rect 3142 12792 3148 12795
rect 3200 12792 3206 12804
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 15120 12841 15148 12872
rect 15948 12841 15976 12872
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14608 12804 14933 12832
rect 14608 12792 14614 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 26878 12832 26884 12844
rect 15979 12804 26884 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 15304 12764 15332 12795
rect 26878 12792 26884 12804
rect 26936 12792 26942 12844
rect 33134 12832 33140 12844
rect 33095 12804 33140 12832
rect 33134 12792 33140 12804
rect 33192 12792 33198 12844
rect 36262 12792 36268 12844
rect 36320 12832 36326 12844
rect 37829 12835 37887 12841
rect 37829 12832 37841 12835
rect 36320 12804 37841 12832
rect 36320 12792 36326 12804
rect 37829 12801 37841 12804
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 21358 12764 21364 12776
rect 14323 12736 21364 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 21358 12724 21364 12736
rect 21416 12724 21422 12776
rect 32953 12767 33011 12773
rect 32953 12733 32965 12767
rect 32999 12733 33011 12767
rect 32953 12727 33011 12733
rect 2038 12696 2044 12708
rect 1999 12668 2044 12696
rect 2038 12656 2044 12668
rect 2096 12656 2102 12708
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 32401 12699 32459 12705
rect 32401 12696 32413 12699
rect 8352 12668 32413 12696
rect 8352 12656 8358 12668
rect 32401 12665 32413 12668
rect 32447 12696 32459 12699
rect 32968 12696 32996 12727
rect 38010 12696 38016 12708
rect 32447 12668 32996 12696
rect 37971 12668 38016 12696
rect 32447 12665 32459 12668
rect 32401 12659 32459 12665
rect 38010 12656 38016 12668
rect 38068 12656 38074 12708
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 4614 12628 4620 12640
rect 4295 12600 4620 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 33321 12631 33379 12637
rect 33321 12597 33333 12631
rect 33367 12628 33379 12631
rect 36630 12628 36636 12640
rect 33367 12600 36636 12628
rect 33367 12597 33379 12600
rect 33321 12591 33379 12597
rect 36630 12588 36636 12600
rect 36688 12588 36694 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1486 12424 1492 12436
rect 1447 12396 1492 12424
rect 1486 12384 1492 12396
rect 1544 12384 1550 12436
rect 3053 12427 3111 12433
rect 3053 12393 3065 12427
rect 3099 12424 3111 12427
rect 3142 12424 3148 12436
rect 3099 12396 3148 12424
rect 3099 12393 3111 12396
rect 3053 12387 3111 12393
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 26878 12384 26884 12436
rect 26936 12424 26942 12436
rect 29825 12427 29883 12433
rect 29825 12424 29837 12427
rect 26936 12396 29837 12424
rect 26936 12384 26942 12396
rect 29825 12393 29837 12396
rect 29871 12424 29883 12427
rect 30374 12424 30380 12436
rect 29871 12396 30380 12424
rect 29871 12393 29883 12396
rect 29825 12387 29883 12393
rect 30374 12384 30380 12396
rect 30432 12384 30438 12436
rect 2317 12359 2375 12365
rect 2317 12325 2329 12359
rect 2363 12356 2375 12359
rect 7374 12356 7380 12368
rect 2363 12328 7380 12356
rect 2363 12325 2375 12328
rect 2317 12319 2375 12325
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 32309 12359 32367 12365
rect 32309 12325 32321 12359
rect 32355 12356 32367 12359
rect 33134 12356 33140 12368
rect 32355 12328 33140 12356
rect 32355 12325 32367 12328
rect 32309 12319 32367 12325
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 2746 12260 4261 12288
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2746 12164 2774 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 4338 12248 4344 12300
rect 4396 12288 4402 12300
rect 4396 12260 4441 12288
rect 4396 12248 4402 12260
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4672 12260 5089 12288
rect 4672 12248 4678 12260
rect 5077 12257 5089 12260
rect 5123 12288 5135 12291
rect 32582 12288 32588 12300
rect 5123 12260 32588 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 32582 12248 32588 12260
rect 32640 12288 32646 12300
rect 32769 12291 32827 12297
rect 32769 12288 32781 12291
rect 32640 12260 32781 12288
rect 32640 12248 32646 12260
rect 32769 12257 32781 12260
rect 32815 12257 32827 12291
rect 32769 12251 32827 12257
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12220 3295 12223
rect 4157 12223 4215 12229
rect 3283 12192 3832 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 2682 12112 2688 12164
rect 2740 12124 2774 12164
rect 2740 12112 2746 12124
rect 3804 12093 3832 12192
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4632 12220 4660 12248
rect 4203 12192 4660 12220
rect 28353 12223 28411 12229
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 28353 12189 28365 12223
rect 28399 12189 28411 12223
rect 28353 12183 28411 12189
rect 23201 12155 23259 12161
rect 23201 12121 23213 12155
rect 23247 12152 23259 12155
rect 24210 12152 24216 12164
rect 23247 12124 24216 12152
rect 23247 12121 23259 12124
rect 23201 12115 23259 12121
rect 24210 12112 24216 12124
rect 24268 12112 24274 12164
rect 27798 12152 27804 12164
rect 27759 12124 27804 12152
rect 27798 12112 27804 12124
rect 27856 12152 27862 12164
rect 28368 12152 28396 12183
rect 28442 12180 28448 12232
rect 28500 12220 28506 12232
rect 28537 12223 28595 12229
rect 28537 12220 28549 12223
rect 28500 12192 28549 12220
rect 28500 12180 28506 12192
rect 28537 12189 28549 12192
rect 28583 12189 28595 12223
rect 30374 12220 30380 12232
rect 30335 12192 30380 12220
rect 28537 12183 28595 12189
rect 30374 12180 30380 12192
rect 30432 12180 30438 12232
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12220 30711 12223
rect 32125 12223 32183 12229
rect 32125 12220 32137 12223
rect 30699 12192 32137 12220
rect 30699 12189 30711 12192
rect 30653 12183 30711 12189
rect 32125 12189 32137 12192
rect 32171 12220 32183 12223
rect 32306 12220 32312 12232
rect 32171 12192 32312 12220
rect 32171 12189 32183 12192
rect 32125 12183 32183 12189
rect 32306 12180 32312 12192
rect 32364 12180 32370 12232
rect 32968 12229 32996 12328
rect 33134 12316 33140 12328
rect 33192 12316 33198 12368
rect 32953 12223 33011 12229
rect 32953 12189 32965 12223
rect 32999 12189 33011 12223
rect 36630 12220 36636 12232
rect 36591 12192 36636 12220
rect 32953 12183 33011 12189
rect 36630 12180 36636 12192
rect 36688 12180 36694 12232
rect 37826 12220 37832 12232
rect 37787 12192 37832 12220
rect 37826 12180 37832 12192
rect 37884 12180 37890 12232
rect 27856 12124 28396 12152
rect 27856 12112 27862 12124
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12053 3847 12087
rect 14550 12084 14556 12096
rect 14511 12056 14556 12084
rect 3789 12047 3847 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 23106 12084 23112 12096
rect 23067 12056 23112 12084
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 28718 12084 28724 12096
rect 28679 12056 28724 12084
rect 28718 12044 28724 12056
rect 28776 12044 28782 12096
rect 33137 12087 33195 12093
rect 33137 12053 33149 12087
rect 33183 12084 33195 12087
rect 34698 12084 34704 12096
rect 33183 12056 34704 12084
rect 33183 12053 33195 12056
rect 33137 12047 33195 12053
rect 34698 12044 34704 12056
rect 34756 12044 34762 12096
rect 36817 12087 36875 12093
rect 36817 12053 36829 12087
rect 36863 12084 36875 12087
rect 37826 12084 37832 12096
rect 36863 12056 37832 12084
rect 36863 12053 36875 12056
rect 36817 12047 36875 12053
rect 37826 12044 37832 12056
rect 37884 12044 37890 12096
rect 38010 12084 38016 12096
rect 37971 12056 38016 12084
rect 38010 12044 38016 12056
rect 38068 12044 38074 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 2130 11880 2136 11892
rect 2091 11852 2136 11880
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 24210 11880 24216 11892
rect 24171 11852 24216 11880
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 32582 11880 32588 11892
rect 32543 11852 32588 11880
rect 32582 11840 32588 11852
rect 32640 11840 32646 11892
rect 2777 11815 2835 11821
rect 2777 11781 2789 11815
rect 2823 11812 2835 11815
rect 2823 11784 2857 11812
rect 2823 11781 2835 11784
rect 2777 11775 2835 11781
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2792 11744 2820 11775
rect 1719 11716 12434 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 12406 11676 12434 11716
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15436 11716 15853 11744
rect 15436 11704 15442 11716
rect 15841 11713 15853 11716
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 24302 11704 24308 11756
rect 24360 11744 24366 11756
rect 24397 11747 24455 11753
rect 24397 11744 24409 11747
rect 24360 11716 24409 11744
rect 24360 11704 24366 11716
rect 24397 11713 24409 11716
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 28718 11704 28724 11756
rect 28776 11744 28782 11756
rect 36541 11747 36599 11753
rect 36541 11744 36553 11747
rect 28776 11716 36553 11744
rect 28776 11704 28782 11716
rect 36541 11713 36553 11716
rect 36587 11713 36599 11747
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 36541 11707 36599 11713
rect 36740 11716 37841 11744
rect 23382 11676 23388 11688
rect 12406 11648 23388 11676
rect 23382 11636 23388 11648
rect 23440 11636 23446 11688
rect 24581 11679 24639 11685
rect 24581 11645 24593 11679
rect 24627 11676 24639 11679
rect 36630 11676 36636 11688
rect 24627 11648 36636 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 36630 11636 36636 11648
rect 36688 11636 36694 11688
rect 1670 11568 1676 11620
rect 1728 11608 1734 11620
rect 3329 11611 3387 11617
rect 3329 11608 3341 11611
rect 1728 11580 3341 11608
rect 1728 11568 1734 11580
rect 3329 11577 3341 11580
rect 3375 11608 3387 11611
rect 23106 11608 23112 11620
rect 3375 11580 23112 11608
rect 3375 11577 3387 11580
rect 3329 11571 3387 11577
rect 23106 11568 23112 11580
rect 23164 11568 23170 11620
rect 36740 11617 36768 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 36725 11611 36783 11617
rect 36725 11577 36737 11611
rect 36771 11577 36783 11611
rect 36725 11571 36783 11577
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 8754 11540 8760 11552
rect 8715 11512 8760 11540
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 17954 11540 17960 11552
rect 16071 11512 17960 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 17954 11500 17960 11512
rect 18012 11500 18018 11552
rect 38010 11540 38016 11552
rect 37971 11512 38016 11540
rect 38010 11500 38016 11512
rect 38068 11500 38074 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 36630 11296 36636 11348
rect 36688 11336 36694 11348
rect 37185 11339 37243 11345
rect 37185 11336 37197 11339
rect 36688 11308 37197 11336
rect 36688 11296 36694 11308
rect 37185 11305 37197 11308
rect 37231 11305 37243 11339
rect 37185 11299 37243 11305
rect 8205 11271 8263 11277
rect 8205 11237 8217 11271
rect 8251 11237 8263 11271
rect 23382 11268 23388 11280
rect 23343 11240 23388 11268
rect 8205 11231 8263 11237
rect 8220 11200 8248 11231
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 34885 11271 34943 11277
rect 34885 11237 34897 11271
rect 34931 11268 34943 11271
rect 35342 11268 35348 11280
rect 34931 11240 35348 11268
rect 34931 11237 34943 11240
rect 34885 11231 34943 11237
rect 35342 11228 35348 11240
rect 35400 11228 35406 11280
rect 38010 11268 38016 11280
rect 37971 11240 38016 11268
rect 38010 11228 38016 11240
rect 38068 11228 38074 11280
rect 22097 11203 22155 11209
rect 22097 11200 22109 11203
rect 8220 11172 9076 11200
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 2774 11132 2780 11144
rect 2547 11104 2780 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 2832 11104 3157 11132
rect 2832 11092 2838 11104
rect 3145 11101 3157 11104
rect 3191 11101 3203 11135
rect 8018 11132 8024 11144
rect 7979 11104 8024 11132
rect 3145 11095 3203 11101
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8754 11132 8760 11144
rect 8352 11104 8760 11132
rect 8352 11092 8358 11104
rect 8754 11092 8760 11104
rect 8812 11132 8818 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8812 11104 8953 11132
rect 8812 11092 8818 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 9048 11132 9076 11172
rect 21468 11172 22109 11200
rect 21468 11144 21496 11172
rect 22097 11169 22109 11172
rect 22143 11169 22155 11203
rect 28629 11203 28687 11209
rect 22097 11163 22155 11169
rect 26206 11172 28580 11200
rect 9197 11135 9255 11141
rect 9197 11132 9209 11135
rect 9048 11104 9209 11132
rect 8941 11095 8999 11101
rect 9197 11101 9209 11104
rect 9243 11101 9255 11135
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 9197 11095 9255 11101
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 19484 11104 21281 11132
rect 19484 11092 19490 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21450 11132 21456 11144
rect 21411 11104 21456 11132
rect 21269 11095 21327 11101
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11132 21695 11135
rect 26206 11132 26234 11172
rect 21683 11104 26234 11132
rect 28261 11135 28319 11141
rect 21683 11101 21695 11104
rect 21637 11095 21695 11101
rect 28261 11101 28273 11135
rect 28307 11101 28319 11135
rect 28442 11132 28448 11144
rect 28403 11104 28448 11132
rect 28261 11095 28319 11101
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2038 11064 2044 11076
rect 1999 11036 2044 11064
rect 2038 11024 2044 11036
rect 2096 11024 2102 11076
rect 23566 11064 23572 11076
rect 23527 11036 23572 11064
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 27706 11064 27712 11076
rect 27667 11036 27712 11064
rect 27706 11024 27712 11036
rect 27764 11064 27770 11076
rect 28276 11064 28304 11095
rect 28442 11092 28448 11104
rect 28500 11092 28506 11144
rect 28552 11132 28580 11172
rect 28629 11169 28641 11203
rect 28675 11200 28687 11203
rect 36998 11200 37004 11212
rect 28675 11172 37004 11200
rect 28675 11169 28687 11172
rect 28629 11163 28687 11169
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 34514 11132 34520 11144
rect 28552 11104 34520 11132
rect 34514 11092 34520 11104
rect 34572 11092 34578 11144
rect 34698 11132 34704 11144
rect 34659 11104 34704 11132
rect 34698 11092 34704 11104
rect 34756 11092 34762 11144
rect 36725 11135 36783 11141
rect 36725 11101 36737 11135
rect 36771 11132 36783 11135
rect 37366 11132 37372 11144
rect 36771 11104 37372 11132
rect 36771 11101 36783 11104
rect 36725 11095 36783 11101
rect 37366 11092 37372 11104
rect 37424 11092 37430 11144
rect 37826 11132 37832 11144
rect 37787 11104 37832 11132
rect 37826 11092 37832 11104
rect 37884 11092 37890 11144
rect 27764 11036 28304 11064
rect 27764 11024 27770 11036
rect 10318 10996 10324 11008
rect 10279 10968 10324 10996
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 18233 10999 18291 11005
rect 18233 10965 18245 10999
rect 18279 10996 18291 10999
rect 18322 10996 18328 11008
rect 18279 10968 18328 10996
rect 18279 10965 18291 10968
rect 18233 10959 18291 10965
rect 18322 10956 18328 10968
rect 18380 10956 18386 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 2133 10795 2191 10801
rect 2133 10792 2145 10795
rect 1912 10764 2145 10792
rect 1912 10752 1918 10764
rect 2133 10761 2145 10764
rect 2179 10761 2191 10795
rect 2133 10755 2191 10761
rect 10137 10795 10195 10801
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 10183 10764 15301 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 9585 10727 9643 10733
rect 1688 10696 2820 10724
rect 1688 10665 1716 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 2792 10597 2820 10696
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 10152 10724 10180 10755
rect 13004 10733 13032 10764
rect 15289 10761 15301 10764
rect 15335 10792 15347 10795
rect 15654 10792 15660 10804
rect 15335 10764 15660 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 19426 10792 19432 10804
rect 19387 10764 19432 10792
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 23566 10752 23572 10804
rect 23624 10792 23630 10804
rect 24397 10795 24455 10801
rect 24397 10792 24409 10795
rect 23624 10764 24409 10792
rect 23624 10752 23630 10764
rect 24397 10761 24409 10764
rect 24443 10761 24455 10795
rect 24397 10755 24455 10761
rect 9631 10696 10180 10724
rect 12989 10727 13047 10733
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 12989 10693 13001 10727
rect 13035 10693 13047 10727
rect 19334 10724 19340 10736
rect 12989 10687 13047 10693
rect 18064 10696 19340 10724
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12308 10628 12357 10656
rect 12308 10616 12314 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 14826 10656 14832 10668
rect 14783 10628 14832 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 14826 10616 14832 10628
rect 14884 10656 14890 10668
rect 18064 10665 18092 10696
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 18322 10665 18328 10668
rect 17589 10659 17647 10665
rect 17589 10656 17601 10659
rect 14884 10628 17601 10656
rect 14884 10616 14890 10628
rect 17589 10625 17601 10628
rect 17635 10656 17647 10659
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17635 10628 18061 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18316 10656 18328 10665
rect 18283 10628 18328 10656
rect 18049 10619 18107 10625
rect 18316 10619 18328 10628
rect 18322 10616 18328 10619
rect 18380 10616 18386 10668
rect 24302 10616 24308 10668
rect 24360 10656 24366 10668
rect 24581 10659 24639 10665
rect 24581 10656 24593 10659
rect 24360 10628 24593 10656
rect 24360 10616 24366 10628
rect 24581 10625 24593 10628
rect 24627 10625 24639 10659
rect 24581 10619 24639 10625
rect 34514 10616 34520 10668
rect 34572 10656 34578 10668
rect 36541 10659 36599 10665
rect 36541 10656 36553 10659
rect 34572 10628 36553 10656
rect 34572 10616 34578 10628
rect 36541 10625 36553 10628
rect 36587 10625 36599 10659
rect 36541 10619 36599 10625
rect 37182 10616 37188 10668
rect 37240 10656 37246 10668
rect 37829 10659 37887 10665
rect 37829 10656 37841 10659
rect 37240 10628 37841 10656
rect 37240 10616 37246 10628
rect 37829 10625 37841 10628
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 24765 10591 24823 10597
rect 2823 10560 12388 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 12360 10532 12388 10560
rect 24765 10557 24777 10591
rect 24811 10588 24823 10591
rect 36354 10588 36360 10600
rect 24811 10560 36360 10588
rect 24811 10557 24823 10560
rect 24765 10551 24823 10557
rect 36354 10548 36360 10560
rect 36412 10548 36418 10600
rect 12342 10480 12348 10532
rect 12400 10480 12406 10532
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 8294 10452 8300 10464
rect 8255 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 36725 10455 36783 10461
rect 36725 10421 36737 10455
rect 36771 10452 36783 10455
rect 37734 10452 37740 10464
rect 36771 10424 37740 10452
rect 36771 10421 36783 10424
rect 36725 10415 36783 10421
rect 37734 10412 37740 10424
rect 37792 10412 37798 10464
rect 38010 10452 38016 10464
rect 37971 10424 38016 10452
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 8076 10220 8125 10248
rect 8076 10208 8082 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 12250 10248 12256 10260
rect 12211 10220 12256 10248
rect 8113 10211 8171 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 17865 10251 17923 10257
rect 12400 10220 17264 10248
rect 12400 10208 12406 10220
rect 2746 10152 11100 10180
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 2746 10044 2774 10152
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 7466 10112 7472 10124
rect 4120 10084 7472 10112
rect 4120 10072 4126 10084
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 7760 10084 9045 10112
rect 2087 10016 2774 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 1854 9976 1860 9988
rect 1815 9948 1860 9976
rect 1854 9936 1860 9948
rect 1912 9976 1918 9988
rect 7760 9985 7788 10084
rect 9033 10081 9045 10084
rect 9079 10112 9091 10115
rect 10318 10112 10324 10124
rect 9079 10084 10324 10112
rect 9079 10081 9091 10084
rect 9033 10075 9091 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 11072 10044 11100 10152
rect 11698 10140 11704 10192
rect 11756 10180 11762 10192
rect 17236 10180 17264 10220
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 18046 10248 18052 10260
rect 17911 10220 18052 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 36354 10248 36360 10260
rect 36315 10220 36360 10248
rect 36354 10208 36360 10220
rect 36412 10208 36418 10260
rect 37182 10248 37188 10260
rect 37143 10220 37188 10248
rect 37182 10208 37188 10220
rect 37240 10208 37246 10260
rect 23017 10183 23075 10189
rect 23017 10180 23029 10183
rect 11756 10152 12848 10180
rect 17236 10152 23029 10180
rect 11756 10140 11762 10152
rect 12710 10112 12716 10124
rect 12671 10084 12716 10112
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 12820 10121 12848 10152
rect 23017 10149 23029 10152
rect 23063 10149 23075 10183
rect 23017 10143 23075 10149
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10112 14427 10115
rect 14826 10112 14832 10124
rect 14415 10084 14832 10112
rect 14415 10081 14427 10084
rect 14369 10075 14427 10081
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 18012 10084 18429 10112
rect 18012 10072 18018 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 18417 10075 18475 10081
rect 28629 10115 28687 10121
rect 28629 10081 28641 10115
rect 28675 10112 28687 10115
rect 36170 10112 36176 10124
rect 28675 10084 36176 10112
rect 28675 10081 28687 10084
rect 28629 10075 28687 10081
rect 36170 10072 36176 10084
rect 36228 10072 36234 10124
rect 27709 10047 27767 10053
rect 27709 10044 27721 10047
rect 11072 10016 27721 10044
rect 27709 10013 27721 10016
rect 27755 10044 27767 10047
rect 28261 10047 28319 10053
rect 28261 10044 28273 10047
rect 27755 10016 28273 10044
rect 27755 10013 27767 10016
rect 27709 10007 27767 10013
rect 28261 10013 28273 10016
rect 28307 10013 28319 10047
rect 28442 10044 28448 10056
rect 28403 10016 28448 10044
rect 28261 10007 28319 10013
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 30098 10044 30104 10056
rect 30059 10016 30104 10044
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 35897 10047 35955 10053
rect 35897 10013 35909 10047
rect 35943 10044 35955 10047
rect 36538 10044 36544 10056
rect 35943 10016 36544 10044
rect 35943 10013 35955 10016
rect 35897 10007 35955 10013
rect 36538 10004 36544 10016
rect 36596 10004 36602 10056
rect 36998 10044 37004 10056
rect 36959 10016 37004 10044
rect 36998 10004 37004 10016
rect 37056 10004 37062 10056
rect 37090 10004 37096 10056
rect 37148 10044 37154 10056
rect 37829 10047 37887 10053
rect 37829 10044 37841 10047
rect 37148 10016 37841 10044
rect 37148 10004 37154 10016
rect 37829 10013 37841 10016
rect 37875 10013 37887 10047
rect 37829 10007 37887 10013
rect 2501 9979 2559 9985
rect 2501 9976 2513 9979
rect 1912 9948 2513 9976
rect 1912 9936 1918 9948
rect 2501 9945 2513 9948
rect 2547 9945 2559 9979
rect 2501 9939 2559 9945
rect 7745 9979 7803 9985
rect 7745 9945 7757 9979
rect 7791 9945 7803 9979
rect 7745 9939 7803 9945
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 15074 9979 15132 9985
rect 15074 9976 15086 9979
rect 12584 9948 15086 9976
rect 12584 9936 12590 9948
rect 15074 9945 15086 9948
rect 15120 9945 15132 9979
rect 15074 9939 15132 9945
rect 15194 9936 15200 9988
rect 15252 9976 15258 9988
rect 17313 9979 17371 9985
rect 17313 9976 17325 9979
rect 15252 9948 17325 9976
rect 15252 9936 15258 9948
rect 17313 9945 17325 9948
rect 17359 9945 17371 9979
rect 17313 9939 17371 9945
rect 18233 9979 18291 9985
rect 18233 9945 18245 9979
rect 18279 9976 18291 9979
rect 19426 9976 19432 9988
rect 18279 9948 19432 9976
rect 18279 9945 18291 9948
rect 18233 9939 18291 9945
rect 3050 9908 3056 9920
rect 3011 9880 3056 9908
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 5592 9880 7665 9908
rect 5592 9868 5598 9880
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 11698 9908 11704 9920
rect 7984 9880 11704 9908
rect 7984 9868 7990 9880
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 12667 9880 13553 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 13541 9877 13553 9880
rect 13587 9908 13599 9911
rect 16206 9908 16212 9920
rect 13587 9880 16212 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 17328 9908 17356 9939
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 23198 9976 23204 9988
rect 23159 9948 23204 9976
rect 23198 9936 23204 9948
rect 23256 9936 23262 9988
rect 29822 9936 29828 9988
rect 29880 9976 29886 9988
rect 29917 9979 29975 9985
rect 29917 9976 29929 9979
rect 29880 9948 29929 9976
rect 29880 9936 29886 9948
rect 29917 9945 29929 9948
rect 29963 9945 29975 9979
rect 29917 9939 29975 9945
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 17328 9880 18337 9908
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 38013 9911 38071 9917
rect 38013 9877 38025 9911
rect 38059 9908 38071 9911
rect 38102 9908 38108 9920
rect 38059 9880 38108 9908
rect 38059 9877 38071 9880
rect 38013 9871 38071 9877
rect 38102 9868 38108 9880
rect 38160 9868 38166 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9673 1639 9707
rect 1581 9667 1639 9673
rect 1596 9636 1624 9667
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 29825 9707 29883 9713
rect 16264 9676 29776 9704
rect 16264 9664 16270 9676
rect 5534 9636 5540 9648
rect 1596 9608 5540 9636
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 24121 9639 24179 9645
rect 24121 9636 24133 9639
rect 23256 9608 24133 9636
rect 23256 9596 23262 9608
rect 24121 9605 24133 9608
rect 24167 9605 24179 9639
rect 24121 9599 24179 9605
rect 27614 9596 27620 9648
rect 27672 9636 27678 9648
rect 28902 9636 28908 9648
rect 27672 9608 28908 9636
rect 27672 9596 27678 9608
rect 28902 9596 28908 9608
rect 28960 9596 28966 9648
rect 29748 9636 29776 9676
rect 29825 9673 29837 9707
rect 29871 9704 29883 9707
rect 30098 9704 30104 9716
rect 29871 9676 30104 9704
rect 29871 9673 29883 9676
rect 29825 9667 29883 9673
rect 30098 9664 30104 9676
rect 30156 9664 30162 9716
rect 36725 9707 36783 9713
rect 36725 9673 36737 9707
rect 36771 9704 36783 9707
rect 37090 9704 37096 9716
rect 36771 9676 37096 9704
rect 36771 9673 36783 9676
rect 36725 9667 36783 9673
rect 37090 9664 37096 9676
rect 37148 9664 37154 9716
rect 31481 9639 31539 9645
rect 31481 9636 31493 9639
rect 29748 9608 31493 9636
rect 31481 9605 31493 9608
rect 31527 9636 31539 9639
rect 31527 9608 32168 9636
rect 31527 9605 31539 9608
rect 31481 9599 31539 9605
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9568 2102 9580
rect 3050 9568 3056 9580
rect 2096 9540 3056 9568
rect 2096 9528 2102 9540
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 24302 9568 24308 9580
rect 24263 9540 24308 9568
rect 24302 9528 24308 9540
rect 24360 9528 24366 9580
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9568 24547 9571
rect 31018 9568 31024 9580
rect 24535 9540 31024 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 32140 9577 32168 9608
rect 35342 9596 35348 9648
rect 35400 9636 35406 9648
rect 35400 9608 37872 9636
rect 35400 9596 35406 9608
rect 32125 9571 32183 9577
rect 32125 9537 32137 9571
rect 32171 9537 32183 9571
rect 32306 9568 32312 9580
rect 32267 9540 32312 9568
rect 32125 9531 32183 9537
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 34333 9571 34391 9577
rect 34333 9537 34345 9571
rect 34379 9568 34391 9571
rect 34790 9568 34796 9580
rect 34379 9540 34796 9568
rect 34379 9537 34391 9540
rect 34333 9531 34391 9537
rect 34790 9528 34796 9540
rect 34848 9528 34854 9580
rect 36170 9528 36176 9580
rect 36228 9568 36234 9580
rect 37844 9577 37872 9608
rect 36541 9571 36599 9577
rect 36541 9568 36553 9571
rect 36228 9540 36553 9568
rect 36228 9528 36234 9540
rect 36541 9537 36553 9540
rect 36587 9537 36599 9571
rect 36541 9531 36599 9537
rect 37829 9571 37887 9577
rect 37829 9537 37841 9571
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 1412 9500 1440 9528
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 1412 9472 2697 9500
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 10318 9460 10324 9512
rect 10376 9500 10382 9512
rect 27065 9503 27123 9509
rect 10376 9472 22094 9500
rect 10376 9460 10382 9472
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 12710 9432 12716 9444
rect 2271 9404 12716 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 22066 9432 22094 9472
rect 27065 9469 27077 9503
rect 27111 9500 27123 9503
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27111 9472 27537 9500
rect 27111 9469 27123 9472
rect 27065 9463 27123 9469
rect 27525 9469 27537 9472
rect 27571 9500 27583 9503
rect 27614 9500 27620 9512
rect 27571 9472 27620 9500
rect 27571 9469 27583 9472
rect 27525 9463 27583 9469
rect 27614 9460 27620 9472
rect 27672 9460 27678 9512
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9500 27859 9503
rect 27890 9500 27896 9512
rect 27847 9472 27896 9500
rect 27847 9469 27859 9472
rect 27801 9463 27859 9469
rect 27890 9460 27896 9472
rect 27948 9460 27954 9512
rect 34149 9503 34207 9509
rect 34149 9469 34161 9503
rect 34195 9469 34207 9503
rect 34149 9463 34207 9469
rect 32493 9435 32551 9441
rect 22066 9404 31340 9432
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 31312 9364 31340 9404
rect 32493 9401 32505 9435
rect 32539 9432 32551 9435
rect 34054 9432 34060 9444
rect 32539 9404 34060 9432
rect 32539 9401 32551 9404
rect 32493 9395 32551 9401
rect 34054 9392 34060 9404
rect 34112 9392 34118 9444
rect 33597 9367 33655 9373
rect 33597 9364 33609 9367
rect 31312 9336 33609 9364
rect 33597 9333 33609 9336
rect 33643 9364 33655 9367
rect 34164 9364 34192 9463
rect 38010 9432 38016 9444
rect 37971 9404 38016 9432
rect 38010 9392 38016 9404
rect 38068 9392 38074 9444
rect 33643 9336 34192 9364
rect 34517 9367 34575 9373
rect 33643 9333 33655 9336
rect 33597 9327 33655 9333
rect 34517 9333 34529 9367
rect 34563 9364 34575 9367
rect 36630 9364 36636 9376
rect 34563 9336 36636 9364
rect 34563 9333 34575 9336
rect 34517 9327 34575 9333
rect 36630 9324 36636 9336
rect 36688 9324 36694 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 4062 9160 4068 9172
rect 3804 9132 4068 9160
rect 3804 9092 3832 9132
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 5166 9092 5172 9104
rect 2746 9064 3832 9092
rect 5079 9064 5172 9092
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 2746 9024 2774 9064
rect 5166 9052 5172 9064
rect 5224 9092 5230 9104
rect 5224 9064 12434 9092
rect 5224 9052 5230 9064
rect 2639 8996 2774 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2682 8956 2688 8968
rect 1719 8928 2688 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 3835 8928 5856 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 2866 8888 2872 8900
rect 2827 8860 2872 8888
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 3418 8848 3424 8900
rect 3476 8888 3482 8900
rect 4034 8891 4092 8897
rect 4034 8888 4046 8891
rect 3476 8860 4046 8888
rect 3476 8848 3482 8860
rect 4034 8857 4046 8860
rect 4080 8857 4092 8891
rect 4034 8851 4092 8857
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 5828 8829 5856 8928
rect 12406 8888 12434 9064
rect 31018 9052 31024 9104
rect 31076 9092 31082 9104
rect 31076 9064 35894 9092
rect 31076 9052 31082 9064
rect 32306 8984 32312 9036
rect 32364 9024 32370 9036
rect 32769 9027 32827 9033
rect 32769 9024 32781 9027
rect 32364 8996 32781 9024
rect 32364 8984 32370 8996
rect 32769 8993 32781 8996
rect 32815 8993 32827 9027
rect 35866 9024 35894 9064
rect 37553 9027 37611 9033
rect 37553 9024 37565 9027
rect 35866 8996 37565 9024
rect 32769 8987 32827 8993
rect 37553 8993 37565 8996
rect 37599 8993 37611 9027
rect 37553 8987 37611 8993
rect 33045 8959 33103 8965
rect 33045 8925 33057 8959
rect 33091 8956 33103 8959
rect 34790 8956 34796 8968
rect 33091 8928 34796 8956
rect 33091 8925 33103 8928
rect 33045 8919 33103 8925
rect 34790 8916 34796 8928
rect 34848 8916 34854 8968
rect 36630 8956 36636 8968
rect 36591 8928 36636 8956
rect 36630 8916 36636 8928
rect 36688 8916 36694 8968
rect 37277 8959 37335 8965
rect 37277 8925 37289 8959
rect 37323 8956 37335 8959
rect 37366 8956 37372 8968
rect 37323 8928 37372 8956
rect 37323 8925 37335 8928
rect 37277 8919 37335 8925
rect 37366 8916 37372 8928
rect 37424 8916 37430 8968
rect 33778 8888 33784 8900
rect 12406 8860 33784 8888
rect 33778 8848 33784 8860
rect 33836 8848 33842 8900
rect 5813 8823 5871 8829
rect 2832 8792 2877 8820
rect 2832 8780 2838 8792
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 8294 8820 8300 8832
rect 5859 8792 8300 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 36817 8823 36875 8829
rect 36817 8789 36829 8823
rect 36863 8820 36875 8823
rect 37826 8820 37832 8832
rect 36863 8792 37832 8820
rect 36863 8789 36875 8792
rect 36817 8783 36875 8789
rect 37826 8780 37832 8792
rect 37884 8780 37890 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 2924 8588 3985 8616
rect 2924 8576 2930 8588
rect 3973 8585 3985 8588
rect 4019 8616 4031 8619
rect 5166 8616 5172 8628
rect 4019 8588 5172 8616
rect 4019 8585 4031 8588
rect 3973 8579 4031 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 33778 8616 33784 8628
rect 33739 8588 33784 8616
rect 33778 8576 33784 8588
rect 33836 8576 33842 8628
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 27157 8483 27215 8489
rect 2915 8452 3464 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3436 8424 3464 8452
rect 27157 8449 27169 8483
rect 27203 8480 27215 8483
rect 27890 8480 27896 8492
rect 27203 8452 27896 8480
rect 27203 8449 27215 8452
rect 27157 8443 27215 8449
rect 27890 8440 27896 8452
rect 27948 8440 27954 8492
rect 33796 8480 33824 8576
rect 34054 8508 34060 8560
rect 34112 8548 34118 8560
rect 37366 8548 37372 8560
rect 34112 8520 35894 8548
rect 37327 8520 37372 8548
rect 34112 8508 34118 8520
rect 34333 8483 34391 8489
rect 34333 8480 34345 8483
rect 33796 8452 34345 8480
rect 34333 8449 34345 8452
rect 34379 8449 34391 8483
rect 34333 8443 34391 8449
rect 34517 8483 34575 8489
rect 34517 8449 34529 8483
rect 34563 8449 34575 8483
rect 35866 8480 35894 8520
rect 37366 8508 37372 8520
rect 37424 8508 37430 8560
rect 36541 8483 36599 8489
rect 36541 8480 36553 8483
rect 35866 8452 36553 8480
rect 34517 8443 34575 8449
rect 36541 8449 36553 8452
rect 36587 8449 36599 8483
rect 37826 8480 37832 8492
rect 37787 8452 37832 8480
rect 36541 8443 36599 8449
rect 3418 8412 3424 8424
rect 3379 8384 3424 8412
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 26421 8415 26479 8421
rect 26421 8412 26433 8415
rect 26206 8384 26433 8412
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 26206 8344 26234 8384
rect 26421 8381 26433 8384
rect 26467 8412 26479 8415
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26467 8384 26985 8412
rect 26467 8381 26479 8384
rect 26421 8375 26479 8381
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 34532 8412 34560 8443
rect 37826 8440 37832 8452
rect 37884 8440 37890 8492
rect 34790 8412 34796 8424
rect 34532 8384 34796 8412
rect 26973 8375 27031 8381
rect 34790 8372 34796 8384
rect 34848 8372 34854 8424
rect 36998 8412 37004 8424
rect 35866 8384 37004 8412
rect 2087 8316 26234 8344
rect 27341 8347 27399 8353
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 27341 8313 27353 8347
rect 27387 8344 27399 8347
rect 35866 8344 35894 8384
rect 36998 8372 37004 8384
rect 37056 8372 37062 8424
rect 27387 8316 35894 8344
rect 36725 8347 36783 8353
rect 27387 8313 27399 8316
rect 27341 8307 27399 8313
rect 36725 8313 36737 8347
rect 36771 8344 36783 8347
rect 37826 8344 37832 8356
rect 36771 8316 37832 8344
rect 36771 8313 36783 8316
rect 36725 8307 36783 8313
rect 37826 8304 37832 8316
rect 37884 8304 37890 8356
rect 38010 8344 38016 8356
rect 37971 8316 38016 8344
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 34698 8276 34704 8288
rect 34659 8248 34704 8276
rect 34698 8236 34704 8248
rect 34756 8236 34762 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2774 8072 2780 8084
rect 1627 8044 2780 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19978 7936 19984 7948
rect 19392 7908 19984 7936
rect 19392 7896 19398 7908
rect 19978 7896 19984 7908
rect 20036 7936 20042 7948
rect 20073 7939 20131 7945
rect 20073 7936 20085 7939
rect 20036 7908 20085 7936
rect 20036 7896 20042 7908
rect 20073 7905 20085 7908
rect 20119 7905 20131 7939
rect 20073 7899 20131 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18656 7840 19257 7868
rect 18656 7828 18662 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 29641 7871 29699 7877
rect 29641 7868 29653 7871
rect 19245 7831 19303 7837
rect 19352 7840 29653 7868
rect 1412 7800 1440 7828
rect 2685 7803 2743 7809
rect 2685 7800 2697 7803
rect 1412 7772 2697 7800
rect 2685 7769 2697 7772
rect 2731 7769 2743 7803
rect 2685 7763 2743 7769
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 19352 7800 19380 7840
rect 29641 7837 29653 7840
rect 29687 7837 29699 7871
rect 29822 7868 29828 7880
rect 29783 7840 29828 7868
rect 29641 7831 29699 7837
rect 29822 7828 29828 7840
rect 29880 7828 29886 7880
rect 30009 7871 30067 7877
rect 30009 7837 30021 7871
rect 30055 7868 30067 7871
rect 36814 7868 36820 7880
rect 30055 7840 36820 7868
rect 30055 7837 30067 7840
rect 30009 7831 30067 7837
rect 36814 7828 36820 7840
rect 36872 7828 36878 7880
rect 36998 7868 37004 7880
rect 36959 7840 37004 7868
rect 36998 7828 37004 7840
rect 37056 7828 37062 7880
rect 37829 7871 37887 7877
rect 37829 7868 37841 7871
rect 37200 7840 37841 7868
rect 20318 7803 20376 7809
rect 20318 7800 20330 7803
rect 3476 7772 19380 7800
rect 19444 7772 20330 7800
rect 3476 7760 3482 7772
rect 2222 7732 2228 7744
rect 2183 7704 2228 7732
rect 2222 7692 2228 7704
rect 2280 7692 2286 7744
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 8113 7735 8171 7741
rect 8113 7732 8125 7735
rect 7432 7704 8125 7732
rect 7432 7692 7438 7704
rect 8113 7701 8125 7704
rect 8159 7732 8171 7735
rect 9674 7732 9680 7744
rect 8159 7704 9680 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 19444 7741 19472 7772
rect 20318 7769 20330 7772
rect 20364 7769 20376 7803
rect 32122 7800 32128 7812
rect 20318 7763 20376 7769
rect 22066 7772 32128 7800
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7701 19487 7735
rect 21450 7732 21456 7744
rect 21411 7704 21456 7732
rect 19429 7695 19487 7701
rect 21450 7692 21456 7704
rect 21508 7732 21514 7744
rect 22066 7732 22094 7772
rect 32122 7760 32128 7772
rect 32180 7760 32186 7812
rect 37200 7741 37228 7840
rect 37829 7837 37841 7840
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 21508 7704 22094 7732
rect 37185 7735 37243 7741
rect 21508 7692 21514 7704
rect 37185 7701 37197 7735
rect 37231 7701 37243 7735
rect 38010 7732 38016 7744
rect 37971 7704 38016 7732
rect 37185 7695 37243 7701
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1854 7488 1860 7540
rect 1912 7528 1918 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1912 7500 2145 7528
rect 1912 7488 1918 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 7285 7531 7343 7537
rect 7285 7528 7297 7531
rect 2280 7500 7297 7528
rect 2280 7488 2286 7500
rect 7285 7497 7297 7500
rect 7331 7497 7343 7531
rect 7285 7491 7343 7497
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 18598 7528 18604 7540
rect 7432 7500 7477 7528
rect 18559 7500 18604 7528
rect 7432 7488 7438 7500
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 19978 7528 19984 7540
rect 19939 7500 19984 7528
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 2038 7420 2044 7472
rect 2096 7460 2102 7472
rect 2777 7463 2835 7469
rect 2777 7460 2789 7463
rect 2096 7432 2789 7460
rect 2096 7420 2102 7432
rect 2777 7429 2789 7432
rect 2823 7429 2835 7463
rect 8294 7460 8300 7472
rect 8207 7432 8300 7460
rect 2777 7423 2835 7429
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2682 7392 2688 7404
rect 1719 7364 2688 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 8220 7401 8248 7432
rect 8294 7420 8300 7432
rect 8352 7460 8358 7472
rect 18233 7463 18291 7469
rect 8352 7432 9628 7460
rect 8352 7420 8358 7432
rect 8478 7401 8484 7404
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8472 7355 8484 7401
rect 8536 7392 8542 7404
rect 8536 7364 8572 7392
rect 8478 7352 8484 7355
rect 8536 7352 8542 7364
rect 9600 7336 9628 7432
rect 18233 7429 18245 7463
rect 18279 7460 18291 7463
rect 21450 7460 21456 7472
rect 18279 7432 21456 7460
rect 18279 7429 18291 7432
rect 18233 7423 18291 7429
rect 21450 7420 21456 7432
rect 21508 7420 21514 7472
rect 31404 7432 32352 7460
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 31404 7401 31432 7432
rect 32324 7404 32352 7432
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 15344 7364 18153 7392
rect 15344 7352 15350 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7361 31447 7395
rect 32122 7392 32128 7404
rect 32083 7364 32128 7392
rect 31389 7355 31447 7361
rect 32122 7352 32128 7364
rect 32180 7352 32186 7404
rect 32306 7392 32312 7404
rect 32267 7364 32312 7392
rect 32306 7352 32312 7364
rect 32364 7352 32370 7404
rect 34698 7352 34704 7404
rect 34756 7392 34762 7404
rect 36541 7395 36599 7401
rect 36541 7392 36553 7395
rect 34756 7364 36553 7392
rect 34756 7352 34762 7364
rect 36541 7361 36553 7364
rect 36587 7361 36599 7395
rect 37826 7392 37832 7404
rect 37787 7364 37832 7392
rect 36541 7355 36599 7361
rect 37826 7352 37832 7364
rect 37884 7352 37890 7404
rect 7190 7324 7196 7336
rect 7103 7296 7196 7324
rect 7190 7284 7196 7296
rect 7248 7324 7254 7336
rect 7926 7324 7932 7336
rect 7248 7296 7932 7324
rect 7248 7284 7254 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9640 7296 10057 7324
rect 9640 7284 9646 7296
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 17954 7324 17960 7336
rect 17915 7296 17960 7324
rect 10045 7287 10103 7293
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 31205 7327 31263 7333
rect 31205 7293 31217 7327
rect 31251 7293 31263 7327
rect 31205 7287 31263 7293
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 7745 7191 7803 7197
rect 7745 7157 7757 7191
rect 7791 7188 7803 7191
rect 8110 7188 8116 7200
rect 7791 7160 8116 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7188 9643 7191
rect 9674 7188 9680 7200
rect 9631 7160 9680 7188
rect 9631 7157 9643 7160
rect 9585 7151 9643 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 30650 7188 30656 7200
rect 30611 7160 30656 7188
rect 30650 7148 30656 7160
rect 30708 7188 30714 7200
rect 31220 7188 31248 7287
rect 31573 7259 31631 7265
rect 31573 7225 31585 7259
rect 31619 7256 31631 7259
rect 33318 7256 33324 7268
rect 31619 7228 33324 7256
rect 31619 7225 31631 7228
rect 31573 7219 31631 7225
rect 33318 7216 33324 7228
rect 33376 7216 33382 7268
rect 30708 7160 31248 7188
rect 32493 7191 32551 7197
rect 30708 7148 30714 7160
rect 32493 7157 32505 7191
rect 32539 7188 32551 7191
rect 32858 7188 32864 7200
rect 32539 7160 32864 7188
rect 32539 7157 32551 7160
rect 32493 7151 32551 7157
rect 32858 7148 32864 7160
rect 32916 7148 32922 7200
rect 36725 7191 36783 7197
rect 36725 7157 36737 7191
rect 36771 7188 36783 7191
rect 37826 7188 37832 7200
rect 36771 7160 37832 7188
rect 36771 7157 36783 7160
rect 36725 7151 36783 7157
rect 37826 7148 37832 7160
rect 37884 7148 37890 7200
rect 38010 7188 38016 7200
rect 37971 7160 38016 7188
rect 38010 7148 38016 7160
rect 38068 7148 38074 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 7926 6984 7932 6996
rect 7699 6956 7932 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 8297 6987 8355 6993
rect 8297 6953 8309 6987
rect 8343 6984 8355 6987
rect 8478 6984 8484 6996
rect 8343 6956 8484 6984
rect 8343 6953 8355 6956
rect 8297 6947 8355 6953
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 30650 6984 30656 6996
rect 9732 6956 30656 6984
rect 9732 6944 9738 6956
rect 30650 6944 30656 6956
rect 30708 6944 30714 6996
rect 36814 6944 36820 6996
rect 36872 6984 36878 6996
rect 37185 6987 37243 6993
rect 37185 6984 37197 6987
rect 36872 6956 37197 6984
rect 36872 6944 36878 6956
rect 37185 6953 37197 6956
rect 37231 6953 37243 6987
rect 37185 6947 37243 6953
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 19334 6848 19340 6860
rect 16071 6820 19340 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 8110 6780 8116 6792
rect 8071 6752 8116 6780
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6780 13047 6783
rect 13262 6780 13268 6792
rect 13035 6752 13268 6780
rect 13035 6749 13047 6752
rect 12989 6743 13047 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 15102 6780 15108 6792
rect 14139 6752 15108 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 16040 6780 16068 6811
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 34054 6848 34060 6860
rect 22066 6820 34060 6848
rect 15160 6752 16068 6780
rect 15160 6740 15166 6752
rect 1854 6712 1860 6724
rect 1815 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 2041 6715 2099 6721
rect 2041 6681 2053 6715
rect 2087 6712 2099 6715
rect 12066 6712 12072 6724
rect 2087 6684 12072 6712
rect 2087 6681 2099 6684
rect 2041 6675 2099 6681
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 13188 6684 14350 6712
rect 1872 6644 1900 6672
rect 13188 6653 13216 6684
rect 14338 6681 14350 6684
rect 14384 6681 14396 6715
rect 22066 6712 22094 6820
rect 34054 6808 34060 6820
rect 34112 6808 34118 6860
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6749 27767 6783
rect 27890 6780 27896 6792
rect 27851 6752 27896 6780
rect 27709 6743 27767 6749
rect 14338 6675 14396 6681
rect 15488 6684 22094 6712
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 1872 6616 2513 6644
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 13173 6647 13231 6653
rect 13173 6613 13185 6647
rect 13219 6613 13231 6647
rect 13173 6607 13231 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 15488 6653 15516 6684
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 13872 6616 15485 6644
rect 13872 6604 13878 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 27157 6647 27215 6653
rect 27157 6644 27169 6647
rect 17276 6616 27169 6644
rect 17276 6604 17282 6616
rect 27157 6613 27169 6616
rect 27203 6644 27215 6647
rect 27724 6644 27752 6743
rect 27890 6740 27896 6752
rect 27948 6740 27954 6792
rect 28077 6783 28135 6789
rect 28077 6749 28089 6783
rect 28123 6780 28135 6783
rect 36538 6780 36544 6792
rect 28123 6752 36544 6780
rect 28123 6749 28135 6752
rect 28077 6743 28135 6749
rect 36538 6740 36544 6752
rect 36596 6740 36602 6792
rect 36725 6783 36783 6789
rect 36725 6749 36737 6783
rect 36771 6780 36783 6783
rect 37366 6780 37372 6792
rect 36771 6752 37372 6780
rect 36771 6749 36783 6752
rect 36725 6743 36783 6749
rect 37366 6740 37372 6752
rect 37424 6740 37430 6792
rect 37826 6780 37832 6792
rect 37787 6752 37832 6780
rect 37826 6740 37832 6752
rect 37884 6740 37890 6792
rect 38010 6644 38016 6656
rect 27203 6616 27752 6644
rect 37971 6616 38016 6644
rect 27203 6613 27215 6616
rect 27157 6607 27215 6613
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2682 6440 2688 6452
rect 2643 6412 2688 6440
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 7984 6412 11989 6440
rect 7984 6400 7990 6412
rect 11977 6409 11989 6412
rect 12023 6409 12035 6443
rect 13262 6440 13268 6452
rect 13223 6412 13268 6440
rect 11977 6403 12035 6409
rect 1964 6344 4660 6372
rect 1964 6313 1992 6344
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 3418 6304 3424 6316
rect 2915 6276 3424 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 2222 6236 2228 6248
rect 2183 6208 2228 6236
rect 2222 6196 2228 6208
rect 2280 6236 2286 6248
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 2280 6208 3893 6236
rect 2280 6196 2286 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 4632 6168 4660 6344
rect 11992 6236 12020 6403
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13814 6440 13820 6452
rect 13775 6412 13820 6440
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 36725 6443 36783 6449
rect 36725 6409 36737 6443
rect 36771 6409 36783 6443
rect 36725 6403 36783 6409
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 17218 6372 17224 6384
rect 12124 6344 17224 6372
rect 12124 6332 12130 6344
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6304 12955 6307
rect 13814 6304 13820 6316
rect 12943 6276 13820 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 24578 6313 24584 6316
rect 24572 6267 24584 6313
rect 24636 6304 24642 6316
rect 33318 6304 33324 6316
rect 24636 6276 24672 6304
rect 33279 6276 33324 6304
rect 24578 6264 24584 6267
rect 24636 6264 24642 6276
rect 33318 6264 33324 6276
rect 33376 6264 33382 6316
rect 36538 6304 36544 6316
rect 36499 6276 36544 6304
rect 36538 6264 36544 6276
rect 36596 6264 36602 6316
rect 36740 6304 36768 6403
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 36740 6276 37841 6304
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 11992 6208 12633 6236
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12802 6236 12808 6248
rect 12763 6208 12808 6236
rect 12621 6199 12679 6205
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 23845 6239 23903 6245
rect 23845 6236 23857 6239
rect 19392 6208 23857 6236
rect 19392 6196 19398 6208
rect 23845 6205 23857 6208
rect 23891 6236 23903 6239
rect 24305 6239 24363 6245
rect 24305 6236 24317 6239
rect 23891 6208 24317 6236
rect 23891 6205 23903 6208
rect 23845 6199 23903 6205
rect 24305 6205 24317 6208
rect 24351 6205 24363 6239
rect 24305 6199 24363 6205
rect 15286 6168 15292 6180
rect 4632 6140 15292 6168
rect 15286 6128 15292 6140
rect 15344 6128 15350 6180
rect 3418 6100 3424 6112
rect 3379 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 25682 6100 25688 6112
rect 25643 6072 25688 6100
rect 25682 6060 25688 6072
rect 25740 6060 25746 6112
rect 33505 6103 33563 6109
rect 33505 6069 33517 6103
rect 33551 6100 33563 6103
rect 37826 6100 37832 6112
rect 33551 6072 37832 6100
rect 33551 6069 33563 6072
rect 33505 6063 33563 6069
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 38010 6100 38016 6112
rect 37971 6072 38016 6100
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 29641 5899 29699 5905
rect 29641 5896 29653 5899
rect 3476 5868 29653 5896
rect 3476 5856 3482 5868
rect 29641 5865 29653 5868
rect 29687 5865 29699 5899
rect 34054 5896 34060 5908
rect 34015 5868 34060 5896
rect 29641 5859 29699 5865
rect 34054 5856 34060 5868
rect 34112 5856 34118 5908
rect 37185 5831 37243 5837
rect 37185 5828 37197 5831
rect 35866 5800 37197 5828
rect 30009 5763 30067 5769
rect 30009 5729 30021 5763
rect 30055 5760 30067 5763
rect 35866 5760 35894 5800
rect 37185 5797 37197 5800
rect 37231 5797 37243 5831
rect 37185 5791 37243 5797
rect 30055 5732 35894 5760
rect 30055 5729 30067 5732
rect 30009 5723 30067 5729
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 2130 5652 2136 5664
rect 2188 5692 2194 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2188 5664 2789 5692
rect 2188 5652 2194 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 29730 5652 29736 5704
rect 29788 5692 29794 5704
rect 29825 5695 29883 5701
rect 29825 5692 29837 5695
rect 29788 5664 29837 5692
rect 29788 5652 29794 5664
rect 29825 5661 29837 5664
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 34054 5652 34060 5704
rect 34112 5692 34118 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 34112 5664 34713 5692
rect 34112 5652 34118 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 34790 5652 34796 5704
rect 34848 5692 34854 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34848 5664 34897 5692
rect 34848 5652 34854 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 36725 5695 36783 5701
rect 36725 5661 36737 5695
rect 36771 5692 36783 5695
rect 37366 5692 37372 5704
rect 36771 5664 37372 5692
rect 36771 5661 36783 5664
rect 36725 5655 36783 5661
rect 37366 5652 37372 5664
rect 37424 5652 37430 5704
rect 37826 5692 37832 5704
rect 37787 5664 37832 5692
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 12802 5624 12808 5636
rect 2332 5596 12808 5624
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2332 5565 2360 5596
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5525 2375 5559
rect 35066 5556 35072 5568
rect 35027 5528 35072 5556
rect 2317 5519 2375 5525
rect 35066 5516 35072 5528
rect 35124 5516 35130 5568
rect 38010 5556 38016 5568
rect 37971 5528 38016 5556
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 36725 5355 36783 5361
rect 36725 5321 36737 5355
rect 36771 5321 36783 5355
rect 36725 5315 36783 5321
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2774 5216 2780 5228
rect 2547 5188 2780 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2774 5176 2780 5188
rect 2832 5216 2838 5228
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 2832 5188 3157 5216
rect 2832 5176 2838 5188
rect 3145 5185 3157 5188
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 35066 5176 35072 5228
rect 35124 5216 35130 5228
rect 36541 5219 36599 5225
rect 36541 5216 36553 5219
rect 35124 5188 36553 5216
rect 35124 5176 35130 5188
rect 36541 5185 36553 5188
rect 36587 5185 36599 5219
rect 36740 5216 36768 5315
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 36740 5188 37841 5216
rect 36541 5179 36599 5185
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 1872 5148 1900 5176
rect 3697 5151 3755 5157
rect 3697 5148 3709 5151
rect 1872 5120 3709 5148
rect 3697 5117 3709 5120
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 2041 5083 2099 5089
rect 2041 5049 2053 5083
rect 2087 5080 2099 5083
rect 27246 5080 27252 5092
rect 2087 5052 27252 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 27246 5040 27252 5052
rect 27304 5040 27310 5092
rect 2685 5015 2743 5021
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 5810 5012 5816 5024
rect 2731 4984 5816 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 38010 5012 38016 5024
rect 37971 4984 38016 5012
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 2685 4811 2743 4817
rect 2685 4808 2697 4811
rect 1728 4780 2697 4808
rect 1728 4768 1734 4780
rect 2685 4777 2697 4780
rect 2731 4777 2743 4811
rect 2685 4771 2743 4777
rect 24118 4768 24124 4820
rect 24176 4808 24182 4820
rect 24397 4811 24455 4817
rect 24397 4808 24409 4811
rect 24176 4780 24409 4808
rect 24176 4768 24182 4780
rect 24397 4777 24409 4780
rect 24443 4777 24455 4811
rect 27246 4808 27252 4820
rect 27207 4780 27252 4808
rect 24397 4771 24455 4777
rect 27246 4768 27252 4780
rect 27304 4768 27310 4820
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4672 2099 4675
rect 5997 4675 6055 4681
rect 2087 4644 5856 4672
rect 2087 4641 2099 4644
rect 2041 4635 2099 4641
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3878 4604 3884 4616
rect 2915 4576 3884 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 5828 4604 5856 4644
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 7190 4672 7196 4684
rect 6043 4644 7196 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 27264 4672 27292 4768
rect 27801 4675 27859 4681
rect 27801 4672 27813 4675
rect 27264 4644 27813 4672
rect 27801 4641 27813 4644
rect 27847 4641 27859 4675
rect 27801 4635 27859 4641
rect 15010 4604 15016 4616
rect 5828 4576 15016 4604
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 24486 4564 24492 4616
rect 24544 4604 24550 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 24544 4576 24593 4604
rect 24544 4564 24550 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 24949 4607 25007 4613
rect 24949 4573 24961 4607
rect 24995 4604 25007 4607
rect 27890 4604 27896 4616
rect 24995 4576 27896 4604
rect 24995 4573 25007 4576
rect 24949 4567 25007 4573
rect 27890 4564 27896 4576
rect 27948 4604 27954 4616
rect 27985 4607 28043 4613
rect 27985 4604 27997 4607
rect 27948 4576 27997 4604
rect 27948 4564 27954 4576
rect 27985 4573 27997 4576
rect 28031 4573 28043 4607
rect 32858 4604 32864 4616
rect 32819 4576 32864 4604
rect 27985 4567 28043 4573
rect 32858 4564 32864 4576
rect 32916 4564 32922 4616
rect 37182 4604 37188 4616
rect 37143 4576 37188 4604
rect 37182 4564 37188 4576
rect 37240 4564 37246 4616
rect 37826 4604 37832 4616
rect 37787 4576 37832 4604
rect 37826 4564 37832 4576
rect 37884 4564 37890 4616
rect 1854 4536 1860 4548
rect 1767 4508 1860 4536
rect 1854 4496 1860 4508
rect 1912 4536 1918 4548
rect 4341 4539 4399 4545
rect 4341 4536 4353 4539
rect 1912 4508 4353 4536
rect 1912 4496 1918 4508
rect 4341 4505 4353 4508
rect 4387 4505 4399 4539
rect 5810 4536 5816 4548
rect 5771 4508 5816 4536
rect 4341 4499 4399 4505
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 24673 4539 24731 4545
rect 24673 4505 24685 4539
rect 24719 4505 24731 4539
rect 24673 4499 24731 4505
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 5132 4440 5365 4468
rect 5132 4428 5138 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5718 4468 5724 4480
rect 5631 4440 5724 4468
rect 5353 4431 5411 4437
rect 5718 4428 5724 4440
rect 5776 4468 5782 4480
rect 6638 4468 6644 4480
rect 5776 4440 6644 4468
rect 5776 4428 5782 4440
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 23750 4468 23756 4480
rect 23711 4440 23756 4468
rect 23750 4428 23756 4440
rect 23808 4468 23814 4480
rect 24688 4468 24716 4499
rect 24762 4496 24768 4548
rect 24820 4536 24826 4548
rect 24820 4508 24865 4536
rect 24820 4496 24826 4508
rect 28166 4468 28172 4480
rect 23808 4440 24716 4468
rect 28127 4440 28172 4468
rect 23808 4428 23814 4440
rect 28166 4428 28172 4440
rect 28224 4428 28230 4480
rect 33045 4471 33103 4477
rect 33045 4437 33057 4471
rect 33091 4468 33103 4471
rect 34514 4468 34520 4480
rect 33091 4440 34520 4468
rect 33091 4437 33103 4440
rect 33045 4431 33103 4437
rect 34514 4428 34520 4440
rect 34572 4428 34578 4480
rect 36078 4428 36084 4480
rect 36136 4468 36142 4480
rect 36173 4471 36231 4477
rect 36173 4468 36185 4471
rect 36136 4440 36185 4468
rect 36136 4428 36142 4440
rect 36173 4437 36185 4440
rect 36219 4437 36231 4471
rect 36173 4431 36231 4437
rect 36354 4428 36360 4480
rect 36412 4468 36418 4480
rect 37001 4471 37059 4477
rect 37001 4468 37013 4471
rect 36412 4440 37013 4468
rect 36412 4428 36418 4440
rect 37001 4437 37013 4440
rect 37047 4437 37059 4471
rect 38010 4468 38016 4480
rect 37971 4440 38016 4468
rect 37001 4431 37059 4437
rect 38010 4428 38016 4440
rect 38068 4428 38074 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 5718 4264 5724 4276
rect 5679 4236 5724 4264
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 6457 4267 6515 4273
rect 6457 4233 6469 4267
rect 6503 4264 6515 4267
rect 7190 4264 7196 4276
rect 6503 4236 7196 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 28166 4224 28172 4276
rect 28224 4264 28230 4276
rect 28224 4236 36584 4264
rect 28224 4224 28230 4236
rect 24213 4199 24271 4205
rect 24213 4196 24225 4199
rect 4540 4168 5028 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2869 4131 2927 4137
rect 1719 4100 2728 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2700 4001 2728 4100
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 2915 4100 3433 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3421 4097 3433 4100
rect 3467 4128 3479 4131
rect 4540 4128 4568 4168
rect 3467 4100 4568 4128
rect 4608 4131 4666 4137
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 4608 4097 4620 4131
rect 4654 4128 4666 4131
rect 4890 4128 4896 4140
rect 4654 4100 4896 4128
rect 4654 4097 4666 4100
rect 4608 4091 4666 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5000 4128 5028 4168
rect 16960 4168 17264 4196
rect 11422 4128 11428 4140
rect 5000 4100 11428 4128
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 16960 4128 16988 4168
rect 16899 4100 16988 4128
rect 17037 4131 17095 4137
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4097 17187 4131
rect 17236 4128 17264 4168
rect 20456 4168 20760 4196
rect 17954 4128 17960 4140
rect 17236 4100 17960 4128
rect 17129 4091 17187 4097
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 2685 3995 2743 4001
rect 2685 3961 2697 3995
rect 2731 3961 2743 3995
rect 2685 3955 2743 3961
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1854 3884 1860 3936
rect 1912 3924 1918 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1912 3896 2145 3924
rect 1912 3884 1918 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 4356 3924 4384 4023
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 17052 4060 17080 4091
rect 15620 4032 17080 4060
rect 17144 4060 17172 4091
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19334 4128 19340 4140
rect 19015 4100 19340 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19334 4088 19340 4100
rect 19392 4128 19398 4140
rect 20456 4128 20484 4168
rect 19392 4100 20484 4128
rect 19392 4088 19398 4100
rect 20530 4088 20536 4140
rect 20588 4137 20594 4140
rect 20588 4128 20600 4137
rect 20732 4128 20760 4168
rect 23952 4168 24225 4196
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20588 4100 20633 4128
rect 20732 4100 20821 4128
rect 20588 4091 20600 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 20809 4091 20867 4097
rect 22480 4100 23029 4128
rect 20588 4088 20594 4091
rect 17144 4032 19748 4060
rect 15620 4020 15626 4032
rect 7558 3952 7564 4004
rect 7616 3992 7622 4004
rect 14550 3992 14556 4004
rect 7616 3964 14556 3992
rect 7616 3952 7622 3964
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 15194 3952 15200 4004
rect 15252 3992 15258 4004
rect 19429 3995 19487 4001
rect 19429 3992 19441 3995
rect 15252 3964 19441 3992
rect 15252 3952 15258 3964
rect 19429 3961 19441 3964
rect 19475 3992 19487 3995
rect 19610 3992 19616 4004
rect 19475 3964 19616 3992
rect 19475 3961 19487 3964
rect 19429 3955 19487 3961
rect 19610 3952 19616 3964
rect 19668 3952 19674 4004
rect 4614 3924 4620 3936
rect 4356 3896 4620 3924
rect 2133 3887 2191 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 19720 3924 19748 4032
rect 20806 3924 20812 3936
rect 19720 3896 20812 3924
rect 20806 3884 20812 3896
rect 20864 3884 20870 3936
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 22002 3924 22008 3936
rect 21416 3896 22008 3924
rect 21416 3884 21422 3896
rect 22002 3884 22008 3896
rect 22060 3924 22066 3936
rect 22480 3933 22508 4100
rect 23017 4097 23029 4100
rect 23063 4097 23075 4131
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 23017 4091 23075 4097
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23109 4063 23167 4069
rect 23109 4029 23121 4063
rect 23155 4060 23167 4063
rect 23952 4060 23980 4168
rect 24213 4165 24225 4168
rect 24259 4196 24271 4199
rect 24762 4196 24768 4208
rect 24259 4168 24768 4196
rect 24259 4165 24271 4168
rect 24213 4159 24271 4165
rect 24762 4156 24768 4168
rect 24820 4156 24826 4208
rect 34790 4196 34796 4208
rect 34348 4168 34796 4196
rect 24029 4131 24087 4137
rect 24029 4097 24041 4131
rect 24075 4097 24087 4131
rect 24029 4091 24087 4097
rect 23155 4032 23980 4060
rect 24044 4060 24072 4091
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 24305 4131 24363 4137
rect 24305 4128 24317 4131
rect 24176 4100 24317 4128
rect 24176 4088 24182 4100
rect 24305 4097 24317 4100
rect 24351 4097 24363 4131
rect 24305 4091 24363 4097
rect 24397 4131 24455 4137
rect 24397 4097 24409 4131
rect 24443 4128 24455 4131
rect 24486 4128 24492 4140
rect 24443 4100 24492 4128
rect 24443 4097 24455 4100
rect 24397 4091 24455 4097
rect 24486 4088 24492 4100
rect 24544 4088 24550 4140
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 28169 4131 28227 4137
rect 28169 4128 28181 4131
rect 25740 4100 28181 4128
rect 25740 4088 25746 4100
rect 28169 4097 28181 4100
rect 28215 4128 28227 4131
rect 28813 4131 28871 4137
rect 28813 4128 28825 4131
rect 28215 4100 28825 4128
rect 28215 4097 28227 4100
rect 28169 4091 28227 4097
rect 28813 4097 28825 4100
rect 28859 4097 28871 4131
rect 28813 4091 28871 4097
rect 29730 4088 29736 4140
rect 29788 4128 29794 4140
rect 30101 4131 30159 4137
rect 30101 4128 30113 4131
rect 29788 4100 30113 4128
rect 29788 4088 29794 4100
rect 30101 4097 30113 4100
rect 30147 4097 30159 4131
rect 30101 4091 30159 4097
rect 30208 4100 33548 4128
rect 28261 4063 28319 4069
rect 24044 4032 26234 4060
rect 23155 4029 23167 4032
rect 23109 4023 23167 4029
rect 24578 3992 24584 4004
rect 24539 3964 24584 3992
rect 24578 3952 24584 3964
rect 24636 3952 24642 4004
rect 26206 3992 26234 4032
rect 28261 4029 28273 4063
rect 28307 4060 28319 4063
rect 30208 4060 30236 4100
rect 28307 4032 30236 4060
rect 30285 4063 30343 4069
rect 28307 4029 28319 4032
rect 28261 4023 28319 4029
rect 30285 4029 30297 4063
rect 30331 4029 30343 4063
rect 30285 4023 30343 4029
rect 29730 3992 29736 4004
rect 26206 3964 29736 3992
rect 29730 3952 29736 3964
rect 29788 3952 29794 4004
rect 29914 3992 29920 4004
rect 29875 3964 29920 3992
rect 29914 3952 29920 3964
rect 29972 3952 29978 4004
rect 30300 3992 30328 4023
rect 32858 4020 32864 4072
rect 32916 4060 32922 4072
rect 33413 4063 33471 4069
rect 33413 4060 33425 4063
rect 32916 4032 33425 4060
rect 32916 4020 32922 4032
rect 33413 4029 33425 4032
rect 33459 4029 33471 4063
rect 33520 4060 33548 4100
rect 33594 4088 33600 4140
rect 33652 4128 33658 4140
rect 34348 4128 34376 4168
rect 34790 4156 34796 4168
rect 34848 4156 34854 4208
rect 35802 4128 35808 4140
rect 33652 4100 34376 4128
rect 34440 4100 35808 4128
rect 33652 4088 33658 4100
rect 34440 4060 34468 4100
rect 35802 4088 35808 4100
rect 35860 4088 35866 4140
rect 36078 4128 36084 4140
rect 36039 4100 36084 4128
rect 36078 4088 36084 4100
rect 36136 4088 36142 4140
rect 36556 4137 36584 4236
rect 36541 4131 36599 4137
rect 36541 4097 36553 4131
rect 36587 4097 36599 4131
rect 36541 4091 36599 4097
rect 37829 4131 37887 4137
rect 37829 4097 37841 4131
rect 37875 4097 37887 4131
rect 37829 4091 37887 4097
rect 33520 4032 34468 4060
rect 33413 4023 33471 4029
rect 34514 4020 34520 4072
rect 34572 4060 34578 4072
rect 37844 4060 37872 4091
rect 34572 4032 37872 4060
rect 34572 4020 34578 4032
rect 35897 3995 35955 4001
rect 35897 3992 35909 3995
rect 30300 3964 35909 3992
rect 35897 3961 35909 3964
rect 35943 3961 35955 3995
rect 35897 3955 35955 3961
rect 36725 3995 36783 4001
rect 36725 3961 36737 3995
rect 36771 3992 36783 3995
rect 37826 3992 37832 4004
rect 36771 3964 37832 3992
rect 36771 3961 36783 3964
rect 36725 3955 36783 3961
rect 37826 3952 37832 3964
rect 37884 3952 37890 4004
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 22060 3896 22477 3924
rect 22060 3884 22066 3896
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 22465 3887 22523 3893
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 31018 3924 31024 3936
rect 23256 3896 31024 3924
rect 23256 3884 23262 3896
rect 31018 3884 31024 3896
rect 31076 3884 31082 3936
rect 32858 3924 32864 3936
rect 32819 3896 32864 3924
rect 32858 3884 32864 3896
rect 32916 3884 32922 3936
rect 33781 3927 33839 3933
rect 33781 3893 33793 3927
rect 33827 3924 33839 3927
rect 35526 3924 35532 3936
rect 33827 3896 35532 3924
rect 33827 3893 33839 3896
rect 33781 3887 33839 3893
rect 35526 3884 35532 3896
rect 35584 3884 35590 3936
rect 38010 3924 38016 3936
rect 37971 3896 38016 3924
rect 38010 3884 38016 3896
rect 38068 3884 38074 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 4890 3720 4896 3732
rect 4851 3692 4896 3720
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 15102 3720 15108 3732
rect 15063 3692 15108 3720
rect 15102 3680 15108 3692
rect 15160 3720 15166 3732
rect 19610 3720 19616 3732
rect 15160 3692 16988 3720
rect 19571 3692 19616 3720
rect 15160 3680 15166 3692
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 5997 3655 6055 3661
rect 5997 3652 6009 3655
rect 4672 3624 6009 3652
rect 4672 3612 4678 3624
rect 5997 3621 6009 3624
rect 6043 3652 6055 3655
rect 15562 3652 15568 3664
rect 6043 3624 9628 3652
rect 15523 3624 15568 3652
rect 6043 3621 6055 3624
rect 5997 3615 6055 3621
rect 9600 3596 9628 3624
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3584 2651 3587
rect 7558 3584 7564 3596
rect 2639 3556 7564 3584
rect 2639 3553 2651 3556
rect 2593 3547 2651 3553
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2685 3479 2743 3485
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 2700 3448 2728 3479
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3878 3516 3884 3528
rect 3344 3488 3884 3516
rect 3344 3448 3372 3488
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 8202 3516 8208 3528
rect 7248 3488 8208 3516
rect 7248 3476 7254 3488
rect 8202 3476 8208 3488
rect 8260 3516 8266 3528
rect 9140 3516 9168 3547
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 16960 3593 16988 3692
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 20530 3680 20536 3732
rect 20588 3720 20594 3732
rect 20625 3723 20683 3729
rect 20625 3720 20637 3723
rect 20588 3692 20637 3720
rect 20588 3680 20594 3692
rect 20625 3689 20637 3692
rect 20671 3689 20683 3723
rect 20625 3683 20683 3689
rect 24118 3680 24124 3732
rect 24176 3720 24182 3732
rect 24489 3723 24547 3729
rect 24489 3720 24501 3723
rect 24176 3692 24501 3720
rect 24176 3680 24182 3692
rect 24489 3689 24501 3692
rect 24535 3689 24547 3723
rect 24489 3683 24547 3689
rect 35069 3723 35127 3729
rect 35069 3689 35081 3723
rect 35115 3720 35127 3723
rect 37826 3720 37832 3732
rect 35115 3692 37832 3720
rect 35115 3689 35127 3692
rect 35069 3683 35127 3689
rect 37826 3680 37832 3692
rect 37884 3680 37890 3732
rect 20257 3655 20315 3661
rect 20257 3621 20269 3655
rect 20303 3652 20315 3655
rect 23198 3652 23204 3664
rect 20303 3624 23204 3652
rect 20303 3621 20315 3624
rect 20257 3615 20315 3621
rect 23198 3612 23204 3624
rect 23256 3612 23262 3664
rect 35713 3655 35771 3661
rect 35713 3621 35725 3655
rect 35759 3621 35771 3655
rect 35713 3615 35771 3621
rect 16945 3587 17003 3593
rect 9640 3556 11100 3584
rect 9640 3544 9646 3556
rect 11072 3528 11100 3556
rect 16945 3553 16957 3587
rect 16991 3553 17003 3587
rect 29917 3587 29975 3593
rect 29917 3584 29929 3587
rect 16945 3547 17003 3553
rect 17236 3556 29929 3584
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 8260 3488 9168 3516
rect 9784 3488 10241 3516
rect 8260 3476 8266 3488
rect 2700 3420 3372 3448
rect 3418 3408 3424 3460
rect 3476 3448 3482 3460
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 3476 3420 9321 3448
rect 3476 3408 3482 3420
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 3786 3380 3792 3392
rect 3747 3352 3792 3380
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 9398 3380 9404 3392
rect 9359 3352 9404 3380
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 9784 3389 9812 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 10229 3479 10287 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 16666 3476 16672 3528
rect 16724 3525 16730 3528
rect 16724 3516 16736 3525
rect 16724 3488 16769 3516
rect 16724 3479 16736 3488
rect 16724 3476 16730 3479
rect 11302 3451 11360 3457
rect 11302 3448 11314 3451
rect 10428 3420 11314 3448
rect 10428 3389 10456 3420
rect 11302 3417 11314 3420
rect 11348 3417 11360 3451
rect 11302 3411 11360 3417
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 17236 3448 17264 3556
rect 29917 3553 29929 3556
rect 29963 3553 29975 3587
rect 35728 3584 35756 3615
rect 35802 3612 35808 3664
rect 35860 3652 35866 3664
rect 36538 3652 36544 3664
rect 35860 3624 36544 3652
rect 35860 3612 35866 3624
rect 36538 3612 36544 3624
rect 36596 3652 36602 3664
rect 37182 3652 37188 3664
rect 36596 3624 37188 3652
rect 36596 3612 36602 3624
rect 37182 3612 37188 3624
rect 37240 3612 37246 3664
rect 35728 3556 37872 3584
rect 29917 3547 29975 3553
rect 19610 3476 19616 3528
rect 19668 3516 19674 3528
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 19668 3488 20177 3516
rect 19668 3476 19674 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 20441 3519 20499 3525
rect 20441 3485 20453 3519
rect 20487 3516 20499 3519
rect 20806 3516 20812 3528
rect 20487 3488 20812 3516
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 20806 3476 20812 3488
rect 20864 3516 20870 3528
rect 21818 3516 21824 3528
rect 20864 3488 21824 3516
rect 20864 3476 20870 3488
rect 21818 3476 21824 3488
rect 21876 3476 21882 3528
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3516 24642 3528
rect 25041 3519 25099 3525
rect 25041 3516 25053 3519
rect 24636 3488 25053 3516
rect 24636 3476 24642 3488
rect 25041 3485 25053 3488
rect 25087 3485 25099 3519
rect 25041 3479 25099 3485
rect 27154 3476 27160 3528
rect 27212 3516 27218 3528
rect 27709 3519 27767 3525
rect 27709 3516 27721 3519
rect 27212 3488 27721 3516
rect 27212 3476 27218 3488
rect 27709 3485 27721 3488
rect 27755 3485 27767 3519
rect 27890 3516 27896 3528
rect 27851 3488 27896 3516
rect 27709 3479 27767 3485
rect 27890 3476 27896 3488
rect 27948 3476 27954 3528
rect 29730 3476 29736 3528
rect 29788 3516 29794 3528
rect 30101 3519 30159 3525
rect 30101 3516 30113 3519
rect 29788 3488 30113 3516
rect 29788 3476 29794 3488
rect 30101 3485 30113 3488
rect 30147 3485 30159 3519
rect 30101 3479 30159 3485
rect 30285 3519 30343 3525
rect 30285 3485 30297 3519
rect 30331 3516 30343 3519
rect 33042 3516 33048 3528
rect 30331 3488 33048 3516
rect 30331 3485 30343 3488
rect 30285 3479 30343 3485
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33321 3519 33379 3525
rect 33321 3485 33333 3519
rect 33367 3485 33379 3519
rect 33321 3479 33379 3485
rect 33505 3519 33563 3525
rect 33505 3485 33517 3519
rect 33551 3516 33563 3519
rect 33594 3516 33600 3528
rect 33551 3488 33600 3516
rect 33551 3485 33563 3488
rect 33505 3479 33563 3485
rect 32769 3451 32827 3457
rect 32769 3448 32781 3451
rect 11480 3420 17264 3448
rect 17328 3420 32781 3448
rect 11480 3408 11486 3420
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3349 9827 3383
rect 9769 3343 9827 3349
rect 10413 3383 10471 3389
rect 10413 3349 10425 3383
rect 10459 3349 10471 3383
rect 10413 3343 10471 3349
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 12437 3383 12495 3389
rect 12437 3380 12449 3383
rect 10560 3352 12449 3380
rect 10560 3340 10566 3352
rect 12437 3349 12449 3352
rect 12483 3380 12495 3383
rect 17328 3380 17356 3420
rect 32769 3417 32781 3420
rect 32815 3448 32827 3451
rect 33336 3448 33364 3479
rect 33594 3476 33600 3488
rect 33652 3476 33658 3528
rect 33689 3519 33747 3525
rect 33689 3485 33701 3519
rect 33735 3516 33747 3519
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 33735 3488 34897 3516
rect 33735 3485 33747 3488
rect 33689 3479 33747 3485
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 35526 3516 35532 3528
rect 35487 3488 35532 3516
rect 34885 3479 34943 3485
rect 35526 3476 35532 3488
rect 35584 3476 35590 3528
rect 36446 3516 36452 3528
rect 36407 3488 36452 3516
rect 36446 3476 36452 3488
rect 36504 3476 36510 3528
rect 37844 3525 37872 3556
rect 37093 3519 37151 3525
rect 37093 3516 37105 3519
rect 36648 3488 37105 3516
rect 32815 3420 33364 3448
rect 32815 3417 32827 3420
rect 32769 3411 32827 3417
rect 27154 3380 27160 3392
rect 12483 3352 17356 3380
rect 27115 3352 27160 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 28074 3380 28080 3392
rect 28035 3352 28080 3380
rect 28074 3340 28080 3352
rect 28132 3340 28138 3392
rect 36648 3389 36676 3488
rect 37093 3485 37105 3488
rect 37139 3485 37151 3519
rect 37093 3479 37151 3485
rect 37829 3519 37887 3525
rect 37829 3485 37841 3519
rect 37875 3485 37887 3519
rect 37829 3479 37887 3485
rect 36633 3383 36691 3389
rect 36633 3349 36645 3383
rect 36679 3349 36691 3383
rect 37274 3380 37280 3392
rect 37235 3352 37280 3380
rect 36633 3343 36691 3349
rect 37274 3340 37280 3352
rect 37332 3340 37338 3392
rect 38010 3380 38016 3392
rect 37971 3352 38016 3380
rect 38010 3340 38016 3352
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3786 3176 3792 3188
rect 1872 3148 3792 3176
rect 1872 3120 1900 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 6696 3148 9076 3176
rect 6696 3136 6702 3148
rect 1854 3108 1860 3120
rect 1767 3080 1860 3108
rect 1854 3068 1860 3080
rect 1912 3068 1918 3120
rect 8938 3108 8944 3120
rect 2792 3080 8944 3108
rect 2792 3049 2820 3080
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 9048 3108 9076 3148
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9456 3148 9965 3176
rect 9456 3136 9462 3148
rect 9953 3145 9965 3148
rect 9999 3176 10011 3179
rect 10502 3176 10508 3188
rect 9999 3148 10508 3176
rect 9999 3145 10011 3148
rect 9953 3139 10011 3145
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11054 3176 11060 3188
rect 11011 3148 11060 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 28074 3136 28080 3188
rect 28132 3176 28138 3188
rect 36446 3176 36452 3188
rect 28132 3148 36452 3176
rect 28132 3136 28138 3148
rect 36446 3136 36452 3148
rect 36504 3136 36510 3188
rect 32858 3108 32864 3120
rect 9048 3080 32864 3108
rect 32858 3068 32864 3080
rect 32916 3068 32922 3120
rect 36633 3111 36691 3117
rect 36633 3108 36645 3111
rect 32968 3080 36645 3108
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 3234 3040 3240 3052
rect 3195 3012 3240 3040
rect 2777 3003 2835 3009
rect 3234 3000 3240 3012
rect 3292 3040 3298 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3292 3012 3893 3040
rect 3292 3000 3298 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8260 3012 8861 3040
rect 8260 3000 8266 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 24486 3040 24492 3052
rect 18012 3012 24492 3040
rect 18012 3000 18018 3012
rect 24486 3000 24492 3012
rect 24544 3000 24550 3052
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 32968 3040 32996 3080
rect 36633 3077 36645 3080
rect 36679 3077 36691 3111
rect 36633 3071 36691 3077
rect 31076 3012 32996 3040
rect 35437 3043 35495 3049
rect 31076 3000 31082 3012
rect 35437 3009 35449 3043
rect 35483 3040 35495 3043
rect 35618 3040 35624 3052
rect 35483 3012 35624 3040
rect 35483 3009 35495 3012
rect 35437 3003 35495 3009
rect 35618 3000 35624 3012
rect 35676 3040 35682 3052
rect 35897 3043 35955 3049
rect 35897 3040 35909 3043
rect 35676 3012 35909 3040
rect 35676 3000 35682 3012
rect 35897 3009 35909 3012
rect 35943 3009 35955 3043
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 35897 3003 35955 3009
rect 36096 3012 36553 3040
rect 1946 2932 1952 2984
rect 2004 2972 2010 2984
rect 27154 2972 27160 2984
rect 2004 2944 27160 2972
rect 2004 2932 2010 2944
rect 27154 2932 27160 2944
rect 27212 2932 27218 2984
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 23750 2904 23756 2916
rect 2087 2876 23756 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 23750 2864 23756 2876
rect 23808 2904 23814 2916
rect 24578 2904 24584 2916
rect 23808 2876 24584 2904
rect 23808 2864 23814 2876
rect 24578 2864 24584 2876
rect 24636 2864 24642 2916
rect 36096 2913 36124 3012
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 37734 3000 37740 3052
rect 37792 3040 37798 3052
rect 37829 3043 37887 3049
rect 37829 3040 37841 3043
rect 37792 3012 37841 3040
rect 37792 3000 37798 3012
rect 37829 3009 37841 3012
rect 37875 3009 37887 3043
rect 37829 3003 37887 3009
rect 36081 2907 36139 2913
rect 36081 2873 36093 2907
rect 36127 2873 36139 2907
rect 36081 2867 36139 2873
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 2774 2836 2780 2848
rect 2639 2808 2780 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3418 2836 3424 2848
rect 3379 2808 3424 2836
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 3970 2796 3976 2848
rect 4028 2836 4034 2848
rect 4433 2839 4491 2845
rect 4433 2836 4445 2839
rect 4028 2808 4445 2836
rect 4028 2796 4034 2808
rect 4433 2805 4445 2808
rect 4479 2805 4491 2839
rect 4982 2836 4988 2848
rect 4943 2808 4988 2836
rect 4433 2799 4491 2805
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 15562 2836 15568 2848
rect 8996 2808 15568 2836
rect 8996 2796 9002 2808
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 34790 2836 34796 2848
rect 34751 2808 34796 2836
rect 34790 2796 34796 2808
rect 34848 2796 34854 2848
rect 38013 2839 38071 2845
rect 38013 2805 38025 2839
rect 38059 2836 38071 2839
rect 38102 2836 38108 2848
rect 38059 2808 38108 2836
rect 38059 2805 38071 2808
rect 38013 2799 38071 2805
rect 38102 2796 38108 2808
rect 38160 2796 38166 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3016 2604 3801 2632
rect 3016 2592 3022 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 3936 2604 4445 2632
rect 3936 2592 3942 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 33042 2592 33048 2644
rect 33100 2632 33106 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 33100 2604 35081 2632
rect 33100 2592 33106 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 2179 2536 6914 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 3050 2496 3056 2508
rect 1872 2468 3056 2496
rect 1872 2437 1900 2468
rect 3050 2456 3056 2468
rect 3108 2496 3114 2508
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 3108 2468 5089 2496
rect 3108 2456 3114 2468
rect 5077 2465 5089 2468
rect 5123 2465 5135 2499
rect 6886 2496 6914 2536
rect 35710 2524 35716 2576
rect 35768 2564 35774 2576
rect 36633 2567 36691 2573
rect 36633 2564 36645 2567
rect 35768 2536 36645 2564
rect 35768 2524 35774 2536
rect 36633 2533 36645 2536
rect 36679 2533 36691 2567
rect 36633 2527 36691 2533
rect 22002 2496 22008 2508
rect 6886 2468 22008 2496
rect 5077 2459 5135 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2397 3019 2431
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 2961 2391 3019 2397
rect 2976 2360 3004 2391
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4120 2400 4629 2428
rect 4120 2388 4126 2400
rect 4617 2397 4629 2400
rect 4663 2428 4675 2431
rect 4982 2428 4988 2440
rect 4663 2400 4988 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35250 2428 35256 2440
rect 34848 2400 35256 2428
rect 34848 2388 34854 2400
rect 35250 2388 35256 2400
rect 35308 2388 35314 2440
rect 35989 2431 36047 2437
rect 35989 2397 36001 2431
rect 36035 2428 36047 2431
rect 36354 2428 36360 2440
rect 36035 2400 36360 2428
rect 36035 2397 36047 2400
rect 35989 2391 36047 2397
rect 36354 2388 36360 2400
rect 36412 2388 36418 2440
rect 36449 2431 36507 2437
rect 36449 2397 36461 2431
rect 36495 2428 36507 2431
rect 36538 2428 36544 2440
rect 36495 2400 36544 2428
rect 36495 2397 36507 2400
rect 36449 2391 36507 2397
rect 36538 2388 36544 2400
rect 36596 2388 36602 2440
rect 37826 2428 37832 2440
rect 37787 2400 37832 2428
rect 37826 2388 37832 2400
rect 37884 2388 37890 2440
rect 5629 2363 5687 2369
rect 5629 2360 5641 2363
rect 2976 2332 5641 2360
rect 5629 2329 5641 2332
rect 5675 2360 5687 2363
rect 15194 2360 15200 2372
rect 5675 2332 15200 2360
rect 5675 2329 5687 2332
rect 5629 2323 5687 2329
rect 15194 2320 15200 2332
rect 15252 2320 15258 2372
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2292 2835 2295
rect 2866 2292 2872 2304
rect 2823 2264 2872 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 35802 2292 35808 2304
rect 35763 2264 35808 2292
rect 35802 2252 35808 2264
rect 35860 2252 35866 2304
rect 38010 2292 38016 2304
rect 37971 2264 38016 2292
rect 38010 2252 38016 2264
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 3142 1300 3148 1352
rect 3200 1340 3206 1352
rect 14458 1340 14464 1352
rect 3200 1312 14464 1340
rect 3200 1300 3206 1312
rect 14458 1300 14464 1312
rect 14516 1300 14522 1352
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2596 37408 2648 37460
rect 3884 37340 3936 37392
rect 2044 37315 2096 37324
rect 2044 37281 2053 37315
rect 2053 37281 2087 37315
rect 2087 37281 2096 37315
rect 2044 37272 2096 37281
rect 3700 37272 3752 37324
rect 1860 37247 1912 37256
rect 1860 37213 1869 37247
rect 1869 37213 1903 37247
rect 1903 37213 1912 37247
rect 1860 37204 1912 37213
rect 3884 37247 3936 37256
rect 3884 37213 3893 37247
rect 3893 37213 3927 37247
rect 3927 37213 3936 37247
rect 3884 37204 3936 37213
rect 4620 37204 4672 37256
rect 33876 37247 33928 37256
rect 33876 37213 33885 37247
rect 33885 37213 33919 37247
rect 33919 37213 33928 37247
rect 33876 37204 33928 37213
rect 2596 37179 2648 37188
rect 2596 37145 2605 37179
rect 2605 37145 2639 37179
rect 2639 37145 2648 37179
rect 2596 37136 2648 37145
rect 4068 37179 4120 37188
rect 4068 37145 4077 37179
rect 4077 37145 4111 37179
rect 4111 37145 4120 37179
rect 4068 37136 4120 37145
rect 26792 37136 26844 37188
rect 35072 37204 35124 37256
rect 35716 37247 35768 37256
rect 35716 37213 35725 37247
rect 35725 37213 35759 37247
rect 35759 37213 35768 37247
rect 35716 37204 35768 37213
rect 37188 37272 37240 37324
rect 35440 37136 35492 37188
rect 1768 37068 1820 37120
rect 3884 37068 3936 37120
rect 3976 37068 4028 37120
rect 34520 37068 34572 37120
rect 35348 37068 35400 37120
rect 35808 37068 35860 37120
rect 36636 37111 36688 37120
rect 36636 37077 36645 37111
rect 36645 37077 36679 37111
rect 36679 37077 36688 37111
rect 36636 37068 36688 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 3332 36907 3384 36916
rect 3332 36873 3341 36907
rect 3341 36873 3375 36907
rect 3375 36873 3384 36907
rect 3332 36864 3384 36873
rect 3884 36864 3936 36916
rect 29736 36907 29788 36916
rect 29736 36873 29745 36907
rect 29745 36873 29779 36907
rect 29779 36873 29788 36907
rect 29736 36864 29788 36873
rect 35532 36864 35584 36916
rect 1768 36796 1820 36848
rect 2872 36796 2924 36848
rect 22468 36796 22520 36848
rect 3332 36728 3384 36780
rect 3516 36771 3568 36780
rect 3516 36737 3525 36771
rect 3525 36737 3559 36771
rect 3559 36737 3568 36771
rect 3516 36728 3568 36737
rect 3976 36771 4028 36780
rect 3976 36737 3985 36771
rect 3985 36737 4019 36771
rect 4019 36737 4028 36771
rect 3976 36728 4028 36737
rect 24308 36660 24360 36712
rect 4068 36592 4120 36644
rect 2780 36524 2832 36576
rect 3792 36524 3844 36576
rect 24768 36567 24820 36576
rect 24768 36533 24777 36567
rect 24777 36533 24811 36567
rect 24811 36533 24820 36567
rect 24768 36524 24820 36533
rect 34704 36728 34756 36780
rect 34796 36728 34848 36780
rect 35992 36771 36044 36780
rect 35992 36737 36001 36771
rect 36001 36737 36035 36771
rect 36035 36737 36044 36771
rect 35992 36728 36044 36737
rect 37280 36771 37332 36780
rect 37280 36737 37289 36771
rect 37289 36737 37323 36771
rect 37323 36737 37332 36771
rect 37280 36728 37332 36737
rect 25504 36524 25556 36576
rect 30748 36524 30800 36576
rect 35900 36524 35952 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3332 36320 3384 36372
rect 5172 36363 5224 36372
rect 5172 36329 5181 36363
rect 5181 36329 5215 36363
rect 5215 36329 5224 36363
rect 5172 36320 5224 36329
rect 2136 36252 2188 36304
rect 30288 36320 30340 36372
rect 35716 36320 35768 36372
rect 36176 36363 36228 36372
rect 36176 36329 36185 36363
rect 36185 36329 36219 36363
rect 36219 36329 36228 36363
rect 36176 36320 36228 36329
rect 37188 36320 37240 36372
rect 24308 36252 24360 36304
rect 34796 36252 34848 36304
rect 2780 36159 2832 36168
rect 2780 36125 2789 36159
rect 2789 36125 2823 36159
rect 2823 36125 2832 36159
rect 2780 36116 2832 36125
rect 1860 36091 1912 36100
rect 1860 36057 1869 36091
rect 1869 36057 1903 36091
rect 1903 36057 1912 36091
rect 1860 36048 1912 36057
rect 2872 36048 2924 36100
rect 21456 36159 21508 36168
rect 21456 36125 21465 36159
rect 21465 36125 21499 36159
rect 21499 36125 21508 36159
rect 21456 36116 21508 36125
rect 22468 36159 22520 36168
rect 2596 36023 2648 36032
rect 2596 35989 2605 36023
rect 2605 35989 2639 36023
rect 2639 35989 2648 36023
rect 2596 35980 2648 35989
rect 4160 35980 4212 36032
rect 20444 36023 20496 36032
rect 20444 35989 20453 36023
rect 20453 35989 20487 36023
rect 20487 35989 20496 36023
rect 20444 35980 20496 35989
rect 20536 35980 20588 36032
rect 21916 36048 21968 36100
rect 22468 36125 22477 36159
rect 22477 36125 22511 36159
rect 22511 36125 22520 36159
rect 22468 36116 22520 36125
rect 25504 36116 25556 36168
rect 25964 36159 26016 36168
rect 25964 36125 25973 36159
rect 25973 36125 26007 36159
rect 26007 36125 26016 36159
rect 25964 36116 26016 36125
rect 29736 36184 29788 36236
rect 30012 36116 30064 36168
rect 30748 36159 30800 36168
rect 29828 36048 29880 36100
rect 30748 36125 30757 36159
rect 30757 36125 30791 36159
rect 30791 36125 30800 36159
rect 30748 36116 30800 36125
rect 37372 36184 37424 36236
rect 35532 36116 35584 36168
rect 35992 36159 36044 36168
rect 35992 36125 36001 36159
rect 36001 36125 36035 36159
rect 36035 36125 36044 36159
rect 35992 36116 36044 36125
rect 36360 36116 36412 36168
rect 34520 36048 34572 36100
rect 26792 36023 26844 36032
rect 26792 35989 26801 36023
rect 26801 35989 26835 36023
rect 26835 35989 26844 36023
rect 26792 35980 26844 35989
rect 35440 35980 35492 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 2964 35819 3016 35828
rect 2964 35785 2973 35819
rect 2973 35785 3007 35819
rect 3007 35785 3016 35819
rect 2964 35776 3016 35785
rect 3516 35776 3568 35828
rect 4160 35776 4212 35828
rect 4620 35776 4672 35828
rect 21456 35776 21508 35828
rect 21916 35776 21968 35828
rect 25964 35776 26016 35828
rect 33876 35776 33928 35828
rect 35532 35819 35584 35828
rect 35532 35785 35541 35819
rect 35541 35785 35575 35819
rect 35575 35785 35584 35819
rect 35532 35776 35584 35785
rect 3056 35640 3108 35692
rect 35900 35708 35952 35760
rect 20536 35640 20588 35692
rect 3700 35572 3752 35624
rect 24768 35640 24820 35692
rect 30012 35640 30064 35692
rect 36360 35683 36412 35692
rect 36360 35649 36369 35683
rect 36369 35649 36403 35683
rect 36403 35649 36412 35683
rect 36360 35640 36412 35649
rect 25504 35572 25556 35624
rect 36544 35615 36596 35624
rect 36544 35581 36553 35615
rect 36553 35581 36587 35615
rect 36587 35581 36596 35615
rect 36544 35572 36596 35581
rect 25504 35479 25556 35488
rect 25504 35445 25513 35479
rect 25513 35445 25547 35479
rect 25547 35445 25556 35479
rect 25504 35436 25556 35445
rect 36176 35479 36228 35488
rect 36176 35445 36185 35479
rect 36185 35445 36219 35479
rect 36219 35445 36228 35479
rect 36176 35436 36228 35445
rect 37188 35436 37240 35488
rect 38016 35479 38068 35488
rect 38016 35445 38025 35479
rect 38025 35445 38059 35479
rect 38059 35445 38068 35479
rect 38016 35436 38068 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2780 35232 2832 35284
rect 3976 35275 4028 35284
rect 3976 35241 3985 35275
rect 3985 35241 4019 35275
rect 4019 35241 4028 35275
rect 3976 35232 4028 35241
rect 36544 35275 36596 35284
rect 36544 35241 36553 35275
rect 36553 35241 36587 35275
rect 36587 35241 36596 35275
rect 36544 35232 36596 35241
rect 37372 35164 37424 35216
rect 1492 34935 1544 34944
rect 1492 34901 1501 34935
rect 1501 34901 1535 34935
rect 1535 34901 1544 34935
rect 1492 34892 1544 34901
rect 2228 34935 2280 34944
rect 2228 34901 2237 34935
rect 2237 34901 2271 34935
rect 2271 34901 2280 34935
rect 2228 34892 2280 34901
rect 2688 35028 2740 35080
rect 20444 35028 20496 35080
rect 36728 35071 36780 35080
rect 36728 35037 36737 35071
rect 36737 35037 36771 35071
rect 36771 35037 36780 35071
rect 36728 35028 36780 35037
rect 37188 35028 37240 35080
rect 3976 34960 4028 35012
rect 36176 34960 36228 35012
rect 36820 34960 36872 35012
rect 4620 34892 4672 34944
rect 25504 34892 25556 34944
rect 37280 34892 37332 34944
rect 38016 34935 38068 34944
rect 38016 34901 38025 34935
rect 38025 34901 38059 34935
rect 38059 34901 38068 34935
rect 38016 34892 38068 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2688 34731 2740 34740
rect 2688 34697 2697 34731
rect 2697 34697 2731 34731
rect 2731 34697 2740 34731
rect 2688 34688 2740 34697
rect 3976 34731 4028 34740
rect 3976 34697 3985 34731
rect 3985 34697 4019 34731
rect 4019 34697 4028 34731
rect 3976 34688 4028 34697
rect 1860 34595 1912 34604
rect 1860 34561 1869 34595
rect 1869 34561 1903 34595
rect 1903 34561 1912 34595
rect 1860 34552 1912 34561
rect 37372 34620 37424 34672
rect 30012 34595 30064 34604
rect 30012 34561 30021 34595
rect 30021 34561 30055 34595
rect 30055 34561 30064 34595
rect 30012 34552 30064 34561
rect 37280 34595 37332 34604
rect 37280 34561 37289 34595
rect 37289 34561 37323 34595
rect 37323 34561 37332 34595
rect 37280 34552 37332 34561
rect 36820 34484 36872 34536
rect 36360 34416 36412 34468
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3056 34187 3108 34196
rect 3056 34153 3065 34187
rect 3065 34153 3099 34187
rect 3099 34153 3108 34187
rect 3056 34144 3108 34153
rect 29276 33940 29328 33992
rect 35348 33940 35400 33992
rect 36360 33940 36412 33992
rect 37372 33983 37424 33992
rect 37372 33949 37381 33983
rect 37381 33949 37415 33983
rect 37415 33949 37424 33983
rect 37372 33940 37424 33949
rect 37832 33983 37884 33992
rect 37832 33949 37841 33983
rect 37841 33949 37875 33983
rect 37875 33949 37884 33983
rect 37832 33940 37884 33949
rect 1860 33915 1912 33924
rect 1860 33881 1869 33915
rect 1869 33881 1903 33915
rect 1903 33881 1912 33915
rect 1860 33872 1912 33881
rect 4620 33804 4672 33856
rect 38016 33847 38068 33856
rect 38016 33813 38025 33847
rect 38025 33813 38059 33847
rect 38059 33813 38068 33847
rect 38016 33804 38068 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1952 33600 2004 33652
rect 29276 33643 29328 33652
rect 29276 33609 29285 33643
rect 29285 33609 29319 33643
rect 29319 33609 29328 33643
rect 29276 33600 29328 33609
rect 37832 33600 37884 33652
rect 2688 33464 2740 33516
rect 30012 33507 30064 33516
rect 30012 33473 30021 33507
rect 30021 33473 30055 33507
rect 30055 33473 30064 33507
rect 30012 33464 30064 33473
rect 37832 33507 37884 33516
rect 37832 33473 37841 33507
rect 37841 33473 37875 33507
rect 37875 33473 37884 33507
rect 37832 33464 37884 33473
rect 38108 33328 38160 33380
rect 1492 33303 1544 33312
rect 1492 33269 1501 33303
rect 1501 33269 1535 33303
rect 1535 33269 1544 33303
rect 1492 33260 1544 33269
rect 38016 33303 38068 33312
rect 38016 33269 38025 33303
rect 38025 33269 38059 33303
rect 38059 33269 38068 33303
rect 38016 33260 38068 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 35348 33056 35400 33108
rect 36268 32988 36320 33040
rect 2780 32852 2832 32904
rect 26056 32852 26108 32904
rect 35808 32852 35860 32904
rect 37464 32895 37516 32904
rect 37464 32861 37473 32895
rect 37473 32861 37507 32895
rect 37507 32861 37516 32895
rect 37464 32852 37516 32861
rect 38108 32895 38160 32904
rect 38108 32861 38117 32895
rect 38117 32861 38151 32895
rect 38151 32861 38160 32895
rect 38108 32852 38160 32861
rect 1860 32827 1912 32836
rect 1860 32793 1869 32827
rect 1869 32793 1903 32827
rect 1903 32793 1912 32827
rect 1860 32784 1912 32793
rect 1952 32759 2004 32768
rect 1952 32725 1961 32759
rect 1961 32725 1995 32759
rect 1995 32725 2004 32759
rect 1952 32716 2004 32725
rect 6184 32716 6236 32768
rect 37832 32784 37884 32836
rect 35808 32716 35860 32768
rect 37280 32759 37332 32768
rect 37280 32725 37289 32759
rect 37289 32725 37323 32759
rect 37323 32725 37332 32759
rect 37280 32716 37332 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1952 32512 2004 32564
rect 26056 32555 26108 32564
rect 1860 32444 1912 32496
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 26056 32521 26065 32555
rect 26065 32521 26099 32555
rect 26099 32521 26108 32555
rect 26056 32512 26108 32521
rect 30012 32512 30064 32564
rect 2688 32283 2740 32292
rect 2688 32249 2697 32283
rect 2697 32249 2731 32283
rect 2731 32249 2740 32283
rect 2688 32240 2740 32249
rect 26240 32376 26292 32428
rect 28724 32376 28776 32428
rect 37280 32419 37332 32428
rect 37280 32385 37289 32419
rect 37289 32385 37323 32419
rect 37323 32385 37332 32419
rect 37280 32376 37332 32385
rect 37648 32376 37700 32428
rect 3516 32308 3568 32360
rect 25412 32308 25464 32360
rect 1492 32215 1544 32224
rect 1492 32181 1501 32215
rect 1501 32181 1535 32215
rect 1535 32181 1544 32215
rect 1492 32172 1544 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3516 31968 3568 32020
rect 1676 31900 1728 31952
rect 38016 32011 38068 32020
rect 25412 31943 25464 31952
rect 25412 31909 25421 31943
rect 25421 31909 25455 31943
rect 25455 31909 25464 31943
rect 25412 31900 25464 31909
rect 37280 31943 37332 31952
rect 37280 31909 37289 31943
rect 37289 31909 37323 31943
rect 37323 31909 37332 31943
rect 37280 31900 37332 31909
rect 1860 31807 1912 31816
rect 1860 31773 1869 31807
rect 1869 31773 1903 31807
rect 1903 31773 1912 31807
rect 1860 31764 1912 31773
rect 7656 31807 7708 31816
rect 7656 31773 7665 31807
rect 7665 31773 7699 31807
rect 7699 31773 7708 31807
rect 7656 31764 7708 31773
rect 11980 31807 12032 31816
rect 11980 31773 11989 31807
rect 11989 31773 12023 31807
rect 12023 31773 12032 31807
rect 11980 31764 12032 31773
rect 17408 31764 17460 31816
rect 19064 31764 19116 31816
rect 16856 31739 16908 31748
rect 16856 31705 16890 31739
rect 16890 31705 16908 31739
rect 25412 31764 25464 31816
rect 26240 31764 26292 31816
rect 16856 31696 16908 31705
rect 7288 31628 7340 31680
rect 11888 31628 11940 31680
rect 17960 31671 18012 31680
rect 17960 31637 17969 31671
rect 17969 31637 18003 31671
rect 18003 31637 18012 31671
rect 17960 31628 18012 31637
rect 20996 31671 21048 31680
rect 20996 31637 21005 31671
rect 21005 31637 21039 31671
rect 21039 31637 21048 31671
rect 20996 31628 21048 31637
rect 35900 31764 35952 31816
rect 38016 31977 38025 32011
rect 38025 31977 38059 32011
rect 38059 31977 38068 32011
rect 38016 31968 38068 31977
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 7656 31424 7708 31476
rect 16856 31467 16908 31476
rect 16856 31433 16865 31467
rect 16865 31433 16899 31467
rect 16899 31433 16908 31467
rect 16856 31424 16908 31433
rect 26240 31424 26292 31476
rect 27160 31424 27212 31476
rect 35900 31467 35952 31476
rect 35900 31433 35909 31467
rect 35909 31433 35943 31467
rect 35943 31433 35952 31467
rect 35900 31424 35952 31433
rect 12348 31356 12400 31408
rect 2136 31331 2188 31340
rect 2136 31297 2145 31331
rect 2145 31297 2179 31331
rect 2179 31297 2188 31331
rect 2136 31288 2188 31297
rect 7748 31331 7800 31340
rect 7748 31297 7757 31331
rect 7757 31297 7791 31331
rect 7791 31297 7800 31331
rect 7748 31288 7800 31297
rect 11888 31331 11940 31340
rect 11888 31297 11922 31331
rect 11922 31297 11940 31331
rect 11888 31288 11940 31297
rect 16488 31288 16540 31340
rect 20996 31288 21048 31340
rect 27712 31288 27764 31340
rect 36084 31331 36136 31340
rect 36084 31297 36093 31331
rect 36093 31297 36127 31331
rect 36127 31297 36136 31331
rect 36084 31288 36136 31297
rect 1492 31127 1544 31136
rect 1492 31093 1501 31127
rect 1501 31093 1535 31127
rect 1535 31093 1544 31127
rect 1492 31084 1544 31093
rect 6184 31220 6236 31272
rect 8024 31263 8076 31272
rect 8024 31229 8033 31263
rect 8033 31229 8067 31263
rect 8067 31229 8076 31263
rect 8024 31220 8076 31229
rect 9036 31220 9088 31272
rect 36268 31263 36320 31272
rect 36268 31229 36277 31263
rect 36277 31229 36311 31263
rect 36311 31229 36320 31263
rect 36268 31220 36320 31229
rect 12992 31195 13044 31204
rect 12992 31161 13001 31195
rect 13001 31161 13035 31195
rect 13035 31161 13044 31195
rect 12992 31152 13044 31161
rect 8484 31084 8536 31136
rect 20996 31084 21048 31136
rect 27712 31127 27764 31136
rect 27712 31093 27721 31127
rect 27721 31093 27755 31127
rect 27755 31093 27764 31127
rect 27712 31084 27764 31093
rect 28724 31084 28776 31136
rect 38016 31127 38068 31136
rect 38016 31093 38025 31127
rect 38025 31093 38059 31127
rect 38059 31093 38068 31127
rect 38016 31084 38068 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 9036 30923 9088 30932
rect 9036 30889 9045 30923
rect 9045 30889 9079 30923
rect 9079 30889 9088 30923
rect 9036 30880 9088 30889
rect 11980 30880 12032 30932
rect 8484 30812 8536 30864
rect 36084 30880 36136 30932
rect 37648 30880 37700 30932
rect 16488 30855 16540 30864
rect 16488 30821 16497 30855
rect 16497 30821 16531 30855
rect 16531 30821 16540 30855
rect 16488 30812 16540 30821
rect 12348 30787 12400 30796
rect 12348 30753 12357 30787
rect 12357 30753 12391 30787
rect 12391 30753 12400 30787
rect 12348 30744 12400 30753
rect 16120 30744 16172 30796
rect 7288 30719 7340 30728
rect 7288 30685 7322 30719
rect 7322 30685 7340 30719
rect 7288 30676 7340 30685
rect 12992 30676 13044 30728
rect 19064 30812 19116 30864
rect 17960 30744 18012 30796
rect 1860 30651 1912 30660
rect 1860 30617 1869 30651
rect 1869 30617 1903 30651
rect 1903 30617 1912 30651
rect 1860 30608 1912 30617
rect 1952 30583 2004 30592
rect 1952 30549 1961 30583
rect 1961 30549 1995 30583
rect 1995 30549 2004 30583
rect 1952 30540 2004 30549
rect 7748 30540 7800 30592
rect 35348 30676 35400 30728
rect 35808 30676 35860 30728
rect 37372 30719 37424 30728
rect 37372 30685 37381 30719
rect 37381 30685 37415 30719
rect 37415 30685 37424 30719
rect 37372 30676 37424 30685
rect 37832 30719 37884 30728
rect 37832 30685 37841 30719
rect 37841 30685 37875 30719
rect 37875 30685 37884 30719
rect 37832 30676 37884 30685
rect 36176 30608 36228 30660
rect 16028 30583 16080 30592
rect 16028 30549 16037 30583
rect 16037 30549 16071 30583
rect 16071 30549 16080 30583
rect 16028 30540 16080 30549
rect 20996 30583 21048 30592
rect 20996 30549 21005 30583
rect 21005 30549 21039 30583
rect 21039 30549 21048 30583
rect 20996 30540 21048 30549
rect 21824 30583 21876 30592
rect 21824 30549 21833 30583
rect 21833 30549 21867 30583
rect 21867 30549 21876 30583
rect 21824 30540 21876 30549
rect 37188 30583 37240 30592
rect 37188 30549 37197 30583
rect 37197 30549 37231 30583
rect 37231 30549 37240 30583
rect 37188 30540 37240 30549
rect 38016 30583 38068 30592
rect 38016 30549 38025 30583
rect 38025 30549 38059 30583
rect 38059 30549 38068 30583
rect 38016 30540 38068 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 36176 30311 36228 30320
rect 36176 30277 36185 30311
rect 36185 30277 36219 30311
rect 36219 30277 36228 30311
rect 36176 30268 36228 30277
rect 16028 30200 16080 30252
rect 21824 30200 21876 30252
rect 2228 30175 2280 30184
rect 2228 30141 2237 30175
rect 2237 30141 2271 30175
rect 2271 30141 2280 30175
rect 2228 30132 2280 30141
rect 1952 30064 2004 30116
rect 27160 30243 27212 30252
rect 27160 30209 27169 30243
rect 27169 30209 27203 30243
rect 27203 30209 27212 30243
rect 37648 30268 37700 30320
rect 27160 30200 27212 30209
rect 37188 30200 37240 30252
rect 37464 30200 37516 30252
rect 37280 30132 37332 30184
rect 37832 30064 37884 30116
rect 3332 30039 3384 30048
rect 3332 30005 3341 30039
rect 3341 30005 3375 30039
rect 3375 30005 3384 30039
rect 3332 29996 3384 30005
rect 37372 30039 37424 30048
rect 37372 30005 37381 30039
rect 37381 30005 37415 30039
rect 37415 30005 37424 30039
rect 37372 29996 37424 30005
rect 38108 29996 38160 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3332 29792 3384 29844
rect 35440 29792 35492 29844
rect 3332 29588 3384 29640
rect 26332 29588 26384 29640
rect 37188 29631 37240 29640
rect 37188 29597 37197 29631
rect 37197 29597 37231 29631
rect 37231 29597 37240 29631
rect 37188 29588 37240 29597
rect 37280 29588 37332 29640
rect 1860 29563 1912 29572
rect 1860 29529 1869 29563
rect 1869 29529 1903 29563
rect 1903 29529 1912 29563
rect 1860 29520 1912 29529
rect 2780 29452 2832 29504
rect 37556 29452 37608 29504
rect 38016 29495 38068 29504
rect 38016 29461 38025 29495
rect 38025 29461 38059 29495
rect 38059 29461 38068 29495
rect 38016 29452 38068 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 26332 29291 26384 29300
rect 26332 29257 26341 29291
rect 26341 29257 26375 29291
rect 26375 29257 26384 29291
rect 26332 29248 26384 29257
rect 35440 29291 35492 29300
rect 35440 29257 35449 29291
rect 35449 29257 35483 29291
rect 35483 29257 35492 29291
rect 35440 29248 35492 29257
rect 1860 29180 1912 29232
rect 16304 29112 16356 29164
rect 27160 29155 27212 29164
rect 27160 29121 27169 29155
rect 27169 29121 27203 29155
rect 27203 29121 27212 29155
rect 27160 29112 27212 29121
rect 37372 29112 37424 29164
rect 37648 29180 37700 29232
rect 37556 29155 37608 29164
rect 37556 29121 37565 29155
rect 37565 29121 37599 29155
rect 37599 29121 37608 29155
rect 37556 29112 37608 29121
rect 2228 29087 2280 29096
rect 2228 29053 2237 29087
rect 2237 29053 2271 29087
rect 2271 29053 2280 29087
rect 2228 29044 2280 29053
rect 37464 28976 37516 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 16120 28611 16172 28620
rect 16120 28577 16129 28611
rect 16129 28577 16163 28611
rect 16163 28577 16172 28611
rect 16120 28568 16172 28577
rect 16304 28611 16356 28620
rect 16304 28577 16313 28611
rect 16313 28577 16347 28611
rect 16347 28577 16356 28611
rect 16304 28568 16356 28577
rect 17224 28636 17276 28688
rect 20996 28611 21048 28620
rect 20996 28577 21005 28611
rect 21005 28577 21039 28611
rect 21039 28577 21048 28611
rect 20996 28568 21048 28577
rect 21456 28543 21508 28552
rect 21456 28509 21465 28543
rect 21465 28509 21499 28543
rect 21499 28509 21508 28543
rect 21456 28500 21508 28509
rect 21548 28500 21600 28552
rect 27160 28500 27212 28552
rect 37188 28543 37240 28552
rect 37188 28509 37197 28543
rect 37197 28509 37231 28543
rect 37231 28509 37240 28543
rect 37188 28500 37240 28509
rect 35808 28432 35860 28484
rect 1492 28407 1544 28416
rect 1492 28373 1501 28407
rect 1501 28373 1535 28407
rect 1535 28373 1544 28407
rect 1492 28364 1544 28373
rect 1860 28364 1912 28416
rect 17316 28364 17368 28416
rect 18236 28364 18288 28416
rect 27896 28364 27948 28416
rect 37556 28364 37608 28416
rect 38016 28407 38068 28416
rect 38016 28373 38025 28407
rect 38025 28373 38059 28407
rect 38059 28373 38068 28407
rect 38016 28364 38068 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 17408 28203 17460 28212
rect 17408 28169 17417 28203
rect 17417 28169 17451 28203
rect 17451 28169 17460 28203
rect 17408 28160 17460 28169
rect 35808 28203 35860 28212
rect 35808 28169 35817 28203
rect 35817 28169 35851 28203
rect 35851 28169 35860 28203
rect 35808 28160 35860 28169
rect 17224 28092 17276 28144
rect 1860 28067 1912 28076
rect 1860 28033 1869 28067
rect 1869 28033 1903 28067
rect 1903 28033 1912 28067
rect 1860 28024 1912 28033
rect 2780 28024 2832 28076
rect 18236 28135 18288 28144
rect 18236 28101 18270 28135
rect 18270 28101 18288 28135
rect 18236 28092 18288 28101
rect 27896 28067 27948 28076
rect 27896 28033 27905 28067
rect 27905 28033 27939 28067
rect 27939 28033 27948 28067
rect 27896 28024 27948 28033
rect 37372 28024 37424 28076
rect 37556 28067 37608 28076
rect 37556 28033 37565 28067
rect 37565 28033 37599 28067
rect 37599 28033 37608 28067
rect 37556 28024 37608 28033
rect 37096 27888 37148 27940
rect 2688 27863 2740 27872
rect 2688 27829 2697 27863
rect 2697 27829 2731 27863
rect 2731 27829 2740 27863
rect 2688 27820 2740 27829
rect 17316 27820 17368 27872
rect 21456 27820 21508 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2688 27616 2740 27668
rect 12256 27616 12308 27668
rect 9036 27591 9088 27600
rect 9036 27557 9045 27591
rect 9045 27557 9079 27591
rect 9079 27557 9088 27591
rect 9036 27548 9088 27557
rect 37280 27591 37332 27600
rect 37280 27557 37289 27591
rect 37289 27557 37323 27591
rect 37323 27557 37332 27591
rect 37280 27548 37332 27557
rect 1492 27319 1544 27328
rect 1492 27285 1501 27319
rect 1501 27285 1535 27319
rect 1535 27285 1544 27319
rect 1492 27276 1544 27285
rect 1952 27276 2004 27328
rect 8300 27412 8352 27464
rect 11980 27412 12032 27464
rect 37096 27455 37148 27464
rect 37096 27421 37105 27455
rect 37105 27421 37139 27455
rect 37139 27421 37148 27455
rect 37096 27412 37148 27421
rect 37832 27455 37884 27464
rect 37832 27421 37841 27455
rect 37841 27421 37875 27455
rect 37875 27421 37884 27455
rect 37832 27412 37884 27421
rect 7104 27344 7156 27396
rect 34796 27344 34848 27396
rect 8392 27319 8444 27328
rect 8392 27285 8401 27319
rect 8401 27285 8435 27319
rect 8435 27285 8444 27319
rect 8392 27276 8444 27285
rect 12072 27319 12124 27328
rect 12072 27285 12081 27319
rect 12081 27285 12115 27319
rect 12115 27285 12124 27319
rect 12072 27276 12124 27285
rect 38016 27319 38068 27328
rect 38016 27285 38025 27319
rect 38025 27285 38059 27319
rect 38059 27285 38068 27319
rect 38016 27276 38068 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 12072 27047 12124 27056
rect 12072 27013 12106 27047
rect 12106 27013 12124 27047
rect 12072 27004 12124 27013
rect 16488 26936 16540 26988
rect 23848 26936 23900 26988
rect 31300 26936 31352 26988
rect 2228 26911 2280 26920
rect 2228 26877 2237 26911
rect 2237 26877 2271 26911
rect 2271 26877 2280 26911
rect 2228 26868 2280 26877
rect 10968 26911 11020 26920
rect 10968 26877 10977 26911
rect 10977 26877 11011 26911
rect 11011 26877 11020 26911
rect 10968 26868 11020 26877
rect 1860 26732 1912 26784
rect 13176 26775 13228 26784
rect 13176 26741 13185 26775
rect 13185 26741 13219 26775
rect 13219 26741 13228 26775
rect 13176 26732 13228 26741
rect 23480 26732 23532 26784
rect 37832 26732 37884 26784
rect 38016 26775 38068 26784
rect 38016 26741 38025 26775
rect 38025 26741 38059 26775
rect 38059 26741 38068 26775
rect 38016 26732 38068 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 7104 26571 7156 26580
rect 7104 26537 7113 26571
rect 7113 26537 7147 26571
rect 7147 26537 7156 26571
rect 7104 26528 7156 26537
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 11980 26528 12032 26537
rect 2780 26460 2832 26512
rect 31300 26571 31352 26580
rect 23848 26503 23900 26512
rect 23848 26469 23857 26503
rect 23857 26469 23891 26503
rect 23891 26469 23900 26503
rect 23848 26460 23900 26469
rect 12256 26392 12308 26444
rect 16120 26392 16172 26444
rect 23480 26435 23532 26444
rect 23480 26401 23489 26435
rect 23489 26401 23523 26435
rect 23523 26401 23532 26435
rect 23480 26392 23532 26401
rect 31300 26537 31309 26571
rect 31309 26537 31343 26571
rect 31343 26537 31352 26571
rect 31300 26528 31352 26537
rect 34796 26528 34848 26580
rect 1860 26367 1912 26376
rect 1860 26333 1869 26367
rect 1869 26333 1903 26367
rect 1903 26333 1912 26367
rect 1860 26324 1912 26333
rect 3884 26324 3936 26376
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 6920 26324 6972 26333
rect 13176 26324 13228 26376
rect 23388 26256 23440 26308
rect 29644 26324 29696 26376
rect 35256 26367 35308 26376
rect 35256 26333 35265 26367
rect 35265 26333 35299 26367
rect 35299 26333 35308 26367
rect 35256 26324 35308 26333
rect 38108 26367 38160 26376
rect 38108 26333 38117 26367
rect 38117 26333 38151 26367
rect 38151 26333 38160 26367
rect 38108 26324 38160 26333
rect 8300 26188 8352 26240
rect 10968 26188 11020 26240
rect 37740 26188 37792 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 16488 25984 16540 26036
rect 1952 25916 2004 25968
rect 3792 25916 3844 25968
rect 3884 25916 3936 25968
rect 35256 25984 35308 26036
rect 2964 25891 3016 25900
rect 2964 25857 2998 25891
rect 2998 25857 3016 25891
rect 2964 25848 3016 25857
rect 29644 25891 29696 25900
rect 15844 25780 15896 25832
rect 16120 25780 16172 25832
rect 19340 25780 19392 25832
rect 29644 25857 29653 25891
rect 29653 25857 29687 25891
rect 29687 25857 29696 25891
rect 29644 25848 29696 25857
rect 30012 25848 30064 25900
rect 23388 25780 23440 25832
rect 29000 25780 29052 25832
rect 4068 25687 4120 25696
rect 4068 25653 4077 25687
rect 4077 25653 4111 25687
rect 4111 25653 4120 25687
rect 4068 25644 4120 25653
rect 8300 25644 8352 25696
rect 17040 25644 17092 25696
rect 29000 25687 29052 25696
rect 29000 25653 29009 25687
rect 29009 25653 29043 25687
rect 29043 25653 29052 25687
rect 29000 25644 29052 25653
rect 31484 25644 31536 25696
rect 35440 25891 35492 25900
rect 35440 25857 35449 25891
rect 35449 25857 35483 25891
rect 35483 25857 35492 25891
rect 35440 25848 35492 25857
rect 36452 25848 36504 25900
rect 37740 25848 37792 25900
rect 38016 25755 38068 25764
rect 38016 25721 38025 25755
rect 38025 25721 38059 25755
rect 38059 25721 38068 25755
rect 38016 25712 38068 25721
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2964 25440 3016 25492
rect 3792 25440 3844 25492
rect 6920 25440 6972 25492
rect 29000 25440 29052 25492
rect 35440 25440 35492 25492
rect 7380 25304 7432 25356
rect 38016 25415 38068 25424
rect 38016 25381 38025 25415
rect 38025 25381 38059 25415
rect 38059 25381 38068 25415
rect 38016 25372 38068 25381
rect 2136 25279 2188 25288
rect 2136 25245 2145 25279
rect 2145 25245 2179 25279
rect 2179 25245 2188 25279
rect 2136 25236 2188 25245
rect 2688 25168 2740 25220
rect 1492 25143 1544 25152
rect 1492 25109 1501 25143
rect 1501 25109 1535 25143
rect 1535 25109 1544 25143
rect 1492 25100 1544 25109
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 23388 25279 23440 25288
rect 4068 25100 4120 25152
rect 5540 25100 5592 25152
rect 5632 25100 5684 25152
rect 8392 25168 8444 25220
rect 23388 25245 23397 25279
rect 23397 25245 23431 25279
rect 23431 25245 23440 25279
rect 23388 25236 23440 25245
rect 24860 25236 24912 25288
rect 28724 25279 28776 25288
rect 17224 25143 17276 25152
rect 17224 25109 17233 25143
rect 17233 25109 17267 25143
rect 17267 25109 17276 25143
rect 17224 25100 17276 25109
rect 26240 25100 26292 25152
rect 26516 25143 26568 25152
rect 26516 25109 26525 25143
rect 26525 25109 26559 25143
rect 26559 25109 26568 25143
rect 26516 25100 26568 25109
rect 27620 25100 27672 25152
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 31484 25279 31536 25288
rect 31484 25245 31493 25279
rect 31493 25245 31527 25279
rect 31527 25245 31536 25279
rect 31484 25236 31536 25245
rect 36544 25279 36596 25288
rect 36544 25245 36553 25279
rect 36553 25245 36587 25279
rect 36587 25245 36596 25279
rect 36544 25236 36596 25245
rect 37372 25279 37424 25288
rect 37372 25245 37381 25279
rect 37381 25245 37415 25279
rect 37415 25245 37424 25279
rect 37372 25236 37424 25245
rect 30012 25100 30064 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 2136 24896 2188 24948
rect 19340 24939 19392 24948
rect 19340 24905 19349 24939
rect 19349 24905 19383 24939
rect 19383 24905 19392 24939
rect 19340 24896 19392 24905
rect 37372 24939 37424 24948
rect 37372 24905 37381 24939
rect 37381 24905 37415 24939
rect 37415 24905 37424 24939
rect 37372 24896 37424 24905
rect 26516 24828 26568 24880
rect 1860 24803 1912 24812
rect 1860 24769 1869 24803
rect 1869 24769 1903 24803
rect 1903 24769 1912 24803
rect 1860 24760 1912 24769
rect 8024 24760 8076 24812
rect 15384 24760 15436 24812
rect 17224 24760 17276 24812
rect 23388 24803 23440 24812
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 24860 24760 24912 24812
rect 17408 24692 17460 24744
rect 15844 24624 15896 24676
rect 1952 24599 2004 24608
rect 1952 24565 1961 24599
rect 1961 24565 1995 24599
rect 1995 24565 2004 24599
rect 1952 24556 2004 24565
rect 7380 24556 7432 24608
rect 17132 24556 17184 24608
rect 22652 24599 22704 24608
rect 22652 24565 22661 24599
rect 22661 24565 22695 24599
rect 22695 24565 22704 24599
rect 22652 24556 22704 24565
rect 38016 24599 38068 24608
rect 38016 24565 38025 24599
rect 38025 24565 38059 24599
rect 38059 24565 38068 24599
rect 38016 24556 38068 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1952 24352 2004 24404
rect 5540 24284 5592 24336
rect 22652 24284 22704 24336
rect 5632 24216 5684 24268
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 2688 24191 2740 24200
rect 2688 24157 2697 24191
rect 2697 24157 2731 24191
rect 2731 24157 2740 24191
rect 2688 24148 2740 24157
rect 15384 24148 15436 24200
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 26240 24148 26292 24157
rect 30012 24216 30064 24268
rect 35348 24148 35400 24200
rect 36544 24191 36596 24200
rect 36544 24157 36553 24191
rect 36553 24157 36587 24191
rect 36587 24157 36596 24191
rect 36544 24148 36596 24157
rect 37372 24191 37424 24200
rect 37372 24157 37381 24191
rect 37381 24157 37415 24191
rect 37415 24157 37424 24191
rect 37372 24148 37424 24157
rect 8024 24012 8076 24064
rect 26424 24055 26476 24064
rect 26424 24021 26433 24055
rect 26433 24021 26467 24055
rect 26467 24021 26476 24055
rect 26424 24012 26476 24021
rect 35900 24012 35952 24064
rect 38016 24055 38068 24064
rect 38016 24021 38025 24055
rect 38025 24021 38059 24055
rect 38059 24021 38068 24055
rect 38016 24012 38068 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 8300 23851 8352 23860
rect 8300 23817 8309 23851
rect 8309 23817 8343 23851
rect 8343 23817 8352 23851
rect 8300 23808 8352 23817
rect 37372 23783 37424 23792
rect 37372 23749 37381 23783
rect 37381 23749 37415 23783
rect 37415 23749 37424 23783
rect 37372 23740 37424 23749
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 15660 23672 15712 23724
rect 26424 23672 26476 23724
rect 29828 23536 29880 23588
rect 3148 23511 3200 23520
rect 3148 23477 3157 23511
rect 3157 23477 3191 23511
rect 3191 23477 3200 23511
rect 3148 23468 3200 23477
rect 35348 23511 35400 23520
rect 35348 23477 35357 23511
rect 35357 23477 35391 23511
rect 35391 23477 35400 23511
rect 35348 23468 35400 23477
rect 38016 23511 38068 23520
rect 38016 23477 38025 23511
rect 38025 23477 38059 23511
rect 38059 23477 38068 23511
rect 38016 23468 38068 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1492 23307 1544 23316
rect 1492 23273 1501 23307
rect 1501 23273 1535 23307
rect 1535 23273 1544 23307
rect 1492 23264 1544 23273
rect 3148 23264 3200 23316
rect 7380 23128 7432 23180
rect 2136 23103 2188 23112
rect 2136 23069 2145 23103
rect 2145 23069 2179 23103
rect 2179 23069 2188 23103
rect 2136 23060 2188 23069
rect 8300 23128 8352 23180
rect 9496 23128 9548 23180
rect 29828 23171 29880 23180
rect 29828 23137 29837 23171
rect 29837 23137 29871 23171
rect 29871 23137 29880 23171
rect 29828 23128 29880 23137
rect 35900 23128 35952 23180
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 30012 23103 30064 23112
rect 30012 23069 30021 23103
rect 30021 23069 30055 23103
rect 30055 23069 30064 23103
rect 30012 23060 30064 23069
rect 37372 23103 37424 23112
rect 37372 23069 37381 23103
rect 37381 23069 37415 23103
rect 37415 23069 37424 23103
rect 37372 23060 37424 23069
rect 21456 23035 21508 23044
rect 21088 22924 21140 22976
rect 21456 23001 21465 23035
rect 21465 23001 21499 23035
rect 21499 23001 21508 23035
rect 21456 22992 21508 23001
rect 22008 22967 22060 22976
rect 22008 22933 22017 22967
rect 22017 22933 22051 22967
rect 22051 22933 22060 22967
rect 22008 22924 22060 22933
rect 24952 22924 25004 22976
rect 38016 22967 38068 22976
rect 38016 22933 38025 22967
rect 38025 22933 38059 22967
rect 38059 22933 38068 22967
rect 38016 22924 38068 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9496 22763 9548 22772
rect 9496 22729 9505 22763
rect 9505 22729 9539 22763
rect 9539 22729 9548 22763
rect 9496 22720 9548 22729
rect 23388 22720 23440 22772
rect 22008 22584 22060 22636
rect 24952 22627 25004 22636
rect 24952 22593 24961 22627
rect 24961 22593 24995 22627
rect 24995 22593 25004 22627
rect 24952 22584 25004 22593
rect 30012 22584 30064 22636
rect 34520 22627 34572 22636
rect 34520 22593 34529 22627
rect 34529 22593 34563 22627
rect 34563 22593 34572 22627
rect 34520 22584 34572 22593
rect 37280 22584 37332 22636
rect 26332 22516 26384 22568
rect 29552 22516 29604 22568
rect 37372 22559 37424 22568
rect 37372 22525 37381 22559
rect 37381 22525 37415 22559
rect 37415 22525 37424 22559
rect 37372 22516 37424 22525
rect 1492 22423 1544 22432
rect 1492 22389 1501 22423
rect 1501 22389 1535 22423
rect 1535 22389 1544 22423
rect 1492 22380 1544 22389
rect 1860 22380 1912 22432
rect 3884 22380 3936 22432
rect 25136 22423 25188 22432
rect 25136 22389 25145 22423
rect 25145 22389 25179 22423
rect 25179 22389 25188 22423
rect 25136 22380 25188 22389
rect 29552 22423 29604 22432
rect 29552 22389 29561 22423
rect 29561 22389 29595 22423
rect 29595 22389 29604 22423
rect 29552 22380 29604 22389
rect 30472 22423 30524 22432
rect 30472 22389 30481 22423
rect 30481 22389 30515 22423
rect 30515 22389 30524 22423
rect 30472 22380 30524 22389
rect 38108 22380 38160 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 21088 22219 21140 22228
rect 21088 22185 21097 22219
rect 21097 22185 21131 22219
rect 21131 22185 21140 22219
rect 21088 22176 21140 22185
rect 25136 22176 25188 22228
rect 34520 22176 34572 22228
rect 1860 22015 1912 22024
rect 1860 21981 1869 22015
rect 1869 21981 1903 22015
rect 1903 21981 1912 22015
rect 1860 21972 1912 21981
rect 2780 21972 2832 22024
rect 29552 22040 29604 22092
rect 15108 21904 15160 21956
rect 3976 21836 4028 21888
rect 15200 21836 15252 21888
rect 21088 21972 21140 22024
rect 30472 21972 30524 22024
rect 35900 22015 35952 22024
rect 35900 21981 35909 22015
rect 35909 21981 35943 22015
rect 35943 21981 35952 22015
rect 35900 21972 35952 21981
rect 36084 22015 36136 22024
rect 36084 21981 36093 22015
rect 36093 21981 36127 22015
rect 36127 21981 36136 22015
rect 36084 21972 36136 21981
rect 37280 22040 37332 22092
rect 37372 22015 37424 22024
rect 17132 21836 17184 21888
rect 20720 21836 20772 21888
rect 37372 21981 37381 22015
rect 37381 21981 37415 22015
rect 37415 21981 37424 22015
rect 37372 21972 37424 21981
rect 36084 21836 36136 21888
rect 38016 21879 38068 21888
rect 38016 21845 38025 21879
rect 38025 21845 38059 21879
rect 38059 21845 38068 21879
rect 38016 21836 38068 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3884 21632 3936 21684
rect 8300 21632 8352 21684
rect 15108 21632 15160 21684
rect 15200 21632 15252 21684
rect 20536 21632 20588 21684
rect 21916 21632 21968 21684
rect 24952 21632 25004 21684
rect 25504 21632 25556 21684
rect 25964 21632 26016 21684
rect 2964 21539 3016 21548
rect 2964 21505 2998 21539
rect 2998 21505 3016 21539
rect 2964 21496 3016 21505
rect 15200 21496 15252 21548
rect 20628 21496 20680 21548
rect 25412 21539 25464 21548
rect 25412 21505 25421 21539
rect 25421 21505 25455 21539
rect 25455 21505 25464 21539
rect 25412 21496 25464 21505
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 28448 21539 28500 21548
rect 28448 21505 28457 21539
rect 28457 21505 28491 21539
rect 28491 21505 28500 21539
rect 28448 21496 28500 21505
rect 37832 21539 37884 21548
rect 37832 21505 37841 21539
rect 37841 21505 37875 21539
rect 37875 21505 37884 21539
rect 37832 21496 37884 21505
rect 20352 21471 20404 21480
rect 20352 21437 20361 21471
rect 20361 21437 20395 21471
rect 20395 21437 20404 21471
rect 20352 21428 20404 21437
rect 37464 21428 37516 21480
rect 1492 21335 1544 21344
rect 1492 21301 1501 21335
rect 1501 21301 1535 21335
rect 1535 21301 1544 21335
rect 1492 21292 1544 21301
rect 1860 21292 1912 21344
rect 4620 21292 4672 21344
rect 27620 21292 27672 21344
rect 30104 21292 30156 21344
rect 38108 21292 38160 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2964 21131 3016 21140
rect 2964 21097 2973 21131
rect 2973 21097 3007 21131
rect 3007 21097 3016 21131
rect 2964 21088 3016 21097
rect 4620 21088 4672 21140
rect 20352 21088 20404 21140
rect 25412 21088 25464 21140
rect 28448 21088 28500 21140
rect 3884 21020 3936 21072
rect 15200 21063 15252 21072
rect 3976 20952 4028 21004
rect 7380 20952 7432 21004
rect 12900 20952 12952 21004
rect 15200 21029 15209 21063
rect 15209 21029 15243 21063
rect 15243 21029 15252 21063
rect 15200 21020 15252 21029
rect 25596 21020 25648 21072
rect 4620 20884 4672 20936
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 15292 20884 15344 20936
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 36912 20884 36964 20936
rect 37096 20884 37148 20936
rect 37464 20884 37516 20936
rect 1860 20859 1912 20868
rect 1860 20825 1869 20859
rect 1869 20825 1903 20859
rect 1903 20825 1912 20859
rect 1860 20816 1912 20825
rect 2044 20859 2096 20868
rect 2044 20825 2053 20859
rect 2053 20825 2087 20859
rect 2087 20825 2096 20859
rect 2044 20816 2096 20825
rect 26148 20816 26200 20868
rect 7196 20791 7248 20800
rect 7196 20757 7205 20791
rect 7205 20757 7239 20791
rect 7239 20757 7248 20791
rect 7196 20748 7248 20757
rect 12532 20748 12584 20800
rect 17132 20791 17184 20800
rect 17132 20757 17141 20791
rect 17141 20757 17175 20791
rect 17175 20757 17184 20791
rect 17132 20748 17184 20757
rect 22008 20748 22060 20800
rect 25596 20791 25648 20800
rect 25596 20757 25605 20791
rect 25605 20757 25639 20791
rect 25639 20757 25648 20791
rect 25596 20748 25648 20757
rect 37280 20748 37332 20800
rect 38016 20791 38068 20800
rect 38016 20757 38025 20791
rect 38025 20757 38059 20791
rect 38059 20757 38068 20791
rect 38016 20748 38068 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 7012 20544 7064 20596
rect 15660 20544 15712 20596
rect 26424 20587 26476 20596
rect 26424 20553 26433 20587
rect 26433 20553 26467 20587
rect 26467 20553 26476 20587
rect 26424 20544 26476 20553
rect 37832 20544 37884 20596
rect 2044 20476 2096 20528
rect 2136 20451 2188 20460
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 2136 20417 2145 20451
rect 2145 20417 2179 20451
rect 2179 20417 2188 20451
rect 2136 20408 2188 20417
rect 7472 20408 7524 20460
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 21088 20408 21140 20460
rect 30288 20408 30340 20460
rect 32588 20408 32640 20460
rect 20536 20383 20588 20392
rect 20536 20349 20545 20383
rect 20545 20349 20579 20383
rect 20579 20349 20588 20383
rect 20536 20340 20588 20349
rect 25596 20340 25648 20392
rect 26148 20272 26200 20324
rect 11704 20204 11756 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 25596 20204 25648 20256
rect 37188 20204 37240 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 8300 20000 8352 20052
rect 11704 20000 11756 20052
rect 36912 20043 36964 20052
rect 36912 20009 36921 20043
rect 36921 20009 36955 20043
rect 36955 20009 36964 20043
rect 36912 20000 36964 20009
rect 22008 19864 22060 19916
rect 37280 19907 37332 19916
rect 37280 19873 37289 19907
rect 37289 19873 37323 19907
rect 37323 19873 37332 19907
rect 37280 19864 37332 19873
rect 7196 19839 7248 19848
rect 7196 19805 7230 19839
rect 7230 19805 7248 19839
rect 7196 19796 7248 19805
rect 7472 19796 7524 19848
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 20536 19796 20588 19848
rect 34520 19796 34572 19848
rect 36268 19796 36320 19848
rect 11520 19728 11572 19780
rect 36544 19728 36596 19780
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 12440 19660 12492 19669
rect 30196 19660 30248 19712
rect 38016 19703 38068 19712
rect 38016 19669 38025 19703
rect 38025 19669 38059 19703
rect 38059 19669 38068 19703
rect 38016 19660 38068 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 32588 19499 32640 19508
rect 32588 19465 32597 19499
rect 32597 19465 32631 19499
rect 32631 19465 32640 19499
rect 32588 19456 32640 19465
rect 36268 19456 36320 19508
rect 36544 19456 36596 19508
rect 12532 19388 12584 19440
rect 30104 19388 30156 19440
rect 35348 19388 35400 19440
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 30196 19320 30248 19372
rect 30288 19363 30340 19372
rect 30288 19329 30297 19363
rect 30297 19329 30331 19363
rect 30331 19329 30340 19363
rect 30288 19320 30340 19329
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 20904 19252 20956 19304
rect 1952 19184 2004 19236
rect 36268 19320 36320 19372
rect 37372 19252 37424 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 11704 18912 11756 18964
rect 26332 18912 26384 18964
rect 26884 18912 26936 18964
rect 37372 18955 37424 18964
rect 37372 18921 37381 18955
rect 37381 18921 37415 18955
rect 37415 18921 37424 18955
rect 37372 18912 37424 18921
rect 12900 18776 12952 18828
rect 34520 18776 34572 18828
rect 17132 18708 17184 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 12440 18640 12492 18692
rect 16856 18683 16908 18692
rect 16856 18649 16890 18683
rect 16890 18649 16908 18683
rect 16856 18640 16908 18649
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 17960 18615 18012 18624
rect 11888 18572 11940 18581
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 37188 18751 37240 18760
rect 37188 18717 37197 18751
rect 37197 18717 37231 18751
rect 37231 18717 37240 18751
rect 37188 18708 37240 18717
rect 25780 18640 25832 18692
rect 26148 18683 26200 18692
rect 26148 18649 26157 18683
rect 26157 18649 26191 18683
rect 26191 18649 26200 18683
rect 26148 18640 26200 18649
rect 24308 18572 24360 18624
rect 25596 18615 25648 18624
rect 25596 18581 25605 18615
rect 25605 18581 25639 18615
rect 25639 18581 25648 18615
rect 25596 18572 25648 18581
rect 38016 18615 38068 18624
rect 38016 18581 38025 18615
rect 38025 18581 38059 18615
rect 38059 18581 38068 18615
rect 38016 18572 38068 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1492 18411 1544 18420
rect 1492 18377 1501 18411
rect 1501 18377 1535 18411
rect 1535 18377 1544 18411
rect 1492 18368 1544 18377
rect 1952 18368 2004 18420
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 16672 18275 16724 18284
rect 16672 18241 16681 18275
rect 16681 18241 16715 18275
rect 16715 18241 16724 18275
rect 16672 18232 16724 18241
rect 21088 18232 21140 18284
rect 12440 18164 12492 18216
rect 27620 18232 27672 18284
rect 28908 18275 28960 18284
rect 28908 18241 28917 18275
rect 28917 18241 28951 18275
rect 28951 18241 28960 18275
rect 28908 18232 28960 18241
rect 29736 18232 29788 18284
rect 30288 18300 30340 18352
rect 36268 18232 36320 18284
rect 37924 18164 37976 18216
rect 11888 18096 11940 18148
rect 16856 18139 16908 18148
rect 16856 18105 16865 18139
rect 16865 18105 16899 18139
rect 16899 18105 16908 18139
rect 16856 18096 16908 18105
rect 29460 18096 29512 18148
rect 30288 18096 30340 18148
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 38016 18071 38068 18080
rect 38016 18037 38025 18071
rect 38025 18037 38059 18071
rect 38059 18037 38068 18071
rect 38016 18028 38068 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 15660 17824 15712 17876
rect 16672 17867 16724 17876
rect 16672 17833 16681 17867
rect 16681 17833 16715 17867
rect 16715 17833 16724 17867
rect 16672 17824 16724 17833
rect 25780 17867 25832 17876
rect 25780 17833 25789 17867
rect 25789 17833 25823 17867
rect 25823 17833 25832 17867
rect 25780 17824 25832 17833
rect 29736 17867 29788 17876
rect 29736 17833 29745 17867
rect 29745 17833 29779 17867
rect 29779 17833 29788 17867
rect 29736 17824 29788 17833
rect 37924 17867 37976 17876
rect 37924 17833 37933 17867
rect 37933 17833 37967 17867
rect 37967 17833 37976 17867
rect 37924 17824 37976 17833
rect 16212 17688 16264 17740
rect 17960 17688 18012 17740
rect 22192 17688 22244 17740
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2228 17527 2280 17536
rect 2228 17493 2237 17527
rect 2237 17493 2271 17527
rect 2271 17493 2280 17527
rect 2228 17484 2280 17493
rect 2872 17484 2924 17536
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 24308 17620 24360 17672
rect 36820 17620 36872 17672
rect 38108 17663 38160 17672
rect 38108 17629 38117 17663
rect 38117 17629 38151 17663
rect 38151 17629 38160 17663
rect 38108 17620 38160 17629
rect 14464 17595 14516 17604
rect 14464 17561 14473 17595
rect 14473 17561 14507 17595
rect 14507 17561 14516 17595
rect 14464 17552 14516 17561
rect 24124 17552 24176 17604
rect 11704 17484 11756 17536
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 22560 17484 22612 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8024 17323 8076 17332
rect 4068 17212 4120 17264
rect 6920 17212 6972 17264
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 11704 17280 11756 17332
rect 24308 17323 24360 17332
rect 17132 17212 17184 17264
rect 24308 17289 24317 17323
rect 24317 17289 24351 17323
rect 24351 17289 24360 17323
rect 24308 17280 24360 17289
rect 3056 17187 3108 17196
rect 3056 17153 3090 17187
rect 3090 17153 3108 17187
rect 3056 17144 3108 17153
rect 8024 17144 8076 17196
rect 29184 17144 29236 17196
rect 29460 17187 29512 17196
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 36084 17144 36136 17196
rect 36820 17144 36872 17196
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 5080 16940 5132 16992
rect 12900 16940 12952 16992
rect 14464 16940 14516 16992
rect 21364 16940 21416 16992
rect 29644 16983 29696 16992
rect 29644 16949 29653 16983
rect 29653 16949 29687 16983
rect 29687 16949 29696 16983
rect 29644 16940 29696 16949
rect 37372 16983 37424 16992
rect 37372 16949 37381 16983
rect 37381 16949 37415 16983
rect 37415 16949 37424 16983
rect 37372 16940 37424 16949
rect 38016 16983 38068 16992
rect 38016 16949 38025 16983
rect 38025 16949 38059 16983
rect 38059 16949 38068 16983
rect 38016 16940 38068 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 21364 16736 21416 16788
rect 36084 16779 36136 16788
rect 36084 16745 36093 16779
rect 36093 16745 36127 16779
rect 36127 16745 36136 16779
rect 36084 16736 36136 16745
rect 4620 16668 4672 16720
rect 37832 16736 37884 16788
rect 7472 16600 7524 16652
rect 12900 16600 12952 16652
rect 16212 16600 16264 16652
rect 22560 16643 22612 16652
rect 22560 16609 22569 16643
rect 22569 16609 22603 16643
rect 22603 16609 22612 16643
rect 22560 16600 22612 16609
rect 4528 16532 4580 16584
rect 8024 16532 8076 16584
rect 29644 16532 29696 16584
rect 36268 16575 36320 16584
rect 36268 16541 36277 16575
rect 36277 16541 36311 16575
rect 36311 16541 36320 16575
rect 36268 16532 36320 16541
rect 37372 16575 37424 16584
rect 37372 16541 37381 16575
rect 37381 16541 37415 16575
rect 37415 16541 37424 16575
rect 37372 16532 37424 16541
rect 2872 16464 2924 16516
rect 2780 16396 2832 16448
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 5080 16439 5132 16448
rect 5080 16405 5089 16439
rect 5089 16405 5123 16439
rect 5123 16405 5132 16439
rect 5080 16396 5132 16405
rect 7472 16396 7524 16448
rect 38016 16439 38068 16448
rect 38016 16405 38025 16439
rect 38025 16405 38059 16439
rect 38059 16405 38068 16439
rect 38016 16396 38068 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3056 16192 3108 16244
rect 8024 16124 8076 16176
rect 36268 16124 36320 16176
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 3792 16056 3844 16108
rect 29184 16099 29236 16108
rect 29184 16065 29193 16099
rect 29193 16065 29227 16099
rect 29227 16065 29236 16099
rect 29184 16056 29236 16065
rect 36084 15988 36136 16040
rect 4620 15852 4672 15904
rect 7932 15895 7984 15904
rect 7932 15861 7941 15895
rect 7941 15861 7975 15895
rect 7975 15861 7984 15895
rect 7932 15852 7984 15861
rect 30564 15895 30616 15904
rect 30564 15861 30573 15895
rect 30573 15861 30607 15895
rect 30607 15861 30616 15895
rect 30564 15852 30616 15861
rect 36176 15895 36228 15904
rect 36176 15861 36185 15895
rect 36185 15861 36219 15895
rect 36219 15861 36228 15895
rect 36176 15852 36228 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4620 15648 4672 15700
rect 36176 15648 36228 15700
rect 38016 15691 38068 15700
rect 38016 15657 38025 15691
rect 38025 15657 38059 15691
rect 38059 15657 38068 15691
rect 38016 15648 38068 15657
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 16212 15555 16264 15564
rect 6920 15512 6972 15521
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 3884 15444 3936 15496
rect 8944 15487 8996 15496
rect 8944 15453 8953 15487
rect 8953 15453 8987 15487
rect 8987 15453 8996 15487
rect 8944 15444 8996 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 30564 15444 30616 15496
rect 37832 15487 37884 15496
rect 37832 15453 37841 15487
rect 37841 15453 37875 15487
rect 37875 15453 37884 15487
rect 37832 15444 37884 15453
rect 2780 15351 2832 15360
rect 2780 15317 2789 15351
rect 2789 15317 2823 15351
rect 2823 15317 2832 15351
rect 2780 15308 2832 15317
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 7288 15376 7340 15428
rect 19248 15376 19300 15428
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 11980 15308 12032 15360
rect 17316 15308 17368 15360
rect 36268 15351 36320 15360
rect 36268 15317 36277 15351
rect 36277 15317 36311 15351
rect 36311 15317 36320 15351
rect 36268 15308 36320 15317
rect 37280 15351 37332 15360
rect 37280 15317 37289 15351
rect 37289 15317 37323 15351
rect 37323 15317 37332 15351
rect 37280 15308 37332 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2228 15104 2280 15156
rect 7288 15147 7340 15156
rect 7288 15113 7297 15147
rect 7297 15113 7331 15147
rect 7331 15113 7340 15147
rect 7288 15104 7340 15113
rect 8944 15104 8996 15156
rect 3884 15036 3936 15088
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 6920 14968 6972 15020
rect 11980 15011 12032 15020
rect 11980 14977 12014 15011
rect 12014 14977 12032 15011
rect 11980 14968 12032 14977
rect 17316 15011 17368 15020
rect 17316 14977 17325 15011
rect 17325 14977 17359 15011
rect 17359 14977 17368 15011
rect 17316 14968 17368 14977
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 36084 15147 36136 15156
rect 36084 15113 36093 15147
rect 36093 15113 36127 15147
rect 36127 15113 36136 15147
rect 36084 15104 36136 15113
rect 23664 15011 23716 15020
rect 23664 14977 23673 15011
rect 23673 14977 23707 15011
rect 23707 14977 23716 15011
rect 23664 14968 23716 14977
rect 33232 14968 33284 15020
rect 36268 14968 36320 15020
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 19432 14900 19484 14952
rect 24768 14832 24820 14884
rect 36636 14832 36688 14884
rect 19340 14764 19392 14816
rect 24308 14764 24360 14816
rect 38016 14807 38068 14816
rect 38016 14773 38025 14807
rect 38025 14773 38059 14807
rect 38059 14773 38068 14807
rect 38016 14764 38068 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1952 14560 2004 14612
rect 21364 14560 21416 14612
rect 23664 14560 23716 14612
rect 26148 14560 26200 14612
rect 36636 14560 36688 14612
rect 5080 14492 5132 14544
rect 12900 14424 12952 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 13084 14424 13136 14476
rect 32496 14424 32548 14476
rect 24308 14356 24360 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 24860 14356 24912 14408
rect 26148 14356 26200 14408
rect 21364 14288 21416 14340
rect 27988 14288 28040 14340
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 19340 14220 19392 14272
rect 33232 14356 33284 14408
rect 37188 14356 37240 14408
rect 28448 14220 28500 14272
rect 36268 14220 36320 14272
rect 38016 14263 38068 14272
rect 38016 14229 38025 14263
rect 38025 14229 38059 14263
rect 38059 14229 38068 14263
rect 38016 14220 38068 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 2688 13948 2740 14000
rect 27988 14059 28040 14068
rect 27988 14025 27997 14059
rect 27997 14025 28031 14059
rect 28031 14025 28040 14059
rect 27988 14016 28040 14025
rect 32496 14059 32548 14068
rect 32496 14025 32505 14059
rect 32505 14025 32539 14059
rect 32539 14025 32548 14059
rect 32496 14016 32548 14025
rect 34520 14016 34572 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 24952 13948 25004 14000
rect 24400 13923 24452 13932
rect 2044 13787 2096 13796
rect 2044 13753 2053 13787
rect 2053 13753 2087 13787
rect 2087 13753 2096 13787
rect 2044 13744 2096 13753
rect 7472 13744 7524 13796
rect 8300 13812 8352 13864
rect 21364 13812 21416 13864
rect 21824 13855 21876 13864
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 33140 13880 33192 13932
rect 38108 13923 38160 13932
rect 38108 13889 38117 13923
rect 38117 13889 38151 13923
rect 38151 13889 38160 13923
rect 38108 13880 38160 13889
rect 24860 13812 24912 13864
rect 1952 13676 2004 13728
rect 37832 13676 37884 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1492 13515 1544 13524
rect 1492 13481 1501 13515
rect 1501 13481 1535 13515
rect 1535 13481 1544 13515
rect 1492 13472 1544 13481
rect 4712 13472 4764 13524
rect 24400 13472 24452 13524
rect 2688 13336 2740 13388
rect 34520 13336 34572 13388
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 24308 13268 24360 13320
rect 28448 13311 28500 13320
rect 2044 13200 2096 13252
rect 28448 13277 28457 13311
rect 28457 13277 28491 13311
rect 28491 13277 28500 13311
rect 28448 13268 28500 13277
rect 36084 13311 36136 13320
rect 36084 13277 36093 13311
rect 36093 13277 36127 13311
rect 36127 13277 36136 13311
rect 36084 13268 36136 13277
rect 36268 13268 36320 13320
rect 37832 13311 37884 13320
rect 37832 13277 37841 13311
rect 37841 13277 37875 13311
rect 37875 13277 37884 13311
rect 37832 13268 37884 13277
rect 28632 13175 28684 13184
rect 28632 13141 28641 13175
rect 28641 13141 28675 13175
rect 28675 13141 28684 13175
rect 28632 13132 28684 13141
rect 36268 13175 36320 13184
rect 36268 13141 36277 13175
rect 36277 13141 36311 13175
rect 36311 13141 36320 13175
rect 36268 13132 36320 13141
rect 37832 13132 37884 13184
rect 38016 13175 38068 13184
rect 38016 13141 38025 13175
rect 38025 13141 38059 13175
rect 38059 13141 38068 13175
rect 38016 13132 38068 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4068 12928 4120 12980
rect 15384 12928 15436 12980
rect 28632 12928 28684 12980
rect 36084 12928 36136 12980
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 3148 12835 3200 12844
rect 3148 12801 3182 12835
rect 3182 12801 3200 12835
rect 3148 12792 3200 12801
rect 14556 12792 14608 12844
rect 26884 12792 26936 12844
rect 33140 12835 33192 12844
rect 33140 12801 33149 12835
rect 33149 12801 33183 12835
rect 33183 12801 33192 12835
rect 33140 12792 33192 12801
rect 36268 12792 36320 12844
rect 21364 12724 21416 12776
rect 2044 12699 2096 12708
rect 2044 12665 2053 12699
rect 2053 12665 2087 12699
rect 2087 12665 2096 12699
rect 2044 12656 2096 12665
rect 8300 12656 8352 12708
rect 38016 12699 38068 12708
rect 38016 12665 38025 12699
rect 38025 12665 38059 12699
rect 38059 12665 38068 12699
rect 38016 12656 38068 12665
rect 4620 12588 4672 12640
rect 36636 12588 36688 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1492 12427 1544 12436
rect 1492 12393 1501 12427
rect 1501 12393 1535 12427
rect 1535 12393 1544 12427
rect 1492 12384 1544 12393
rect 3148 12384 3200 12436
rect 26884 12384 26936 12436
rect 30380 12384 30432 12436
rect 7380 12316 7432 12368
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 4620 12248 4672 12300
rect 32588 12248 32640 12300
rect 2688 12112 2740 12164
rect 24216 12112 24268 12164
rect 27804 12155 27856 12164
rect 27804 12121 27813 12155
rect 27813 12121 27847 12155
rect 27847 12121 27856 12155
rect 28448 12180 28500 12232
rect 30380 12223 30432 12232
rect 30380 12189 30389 12223
rect 30389 12189 30423 12223
rect 30423 12189 30432 12223
rect 30380 12180 30432 12189
rect 32312 12180 32364 12232
rect 33140 12316 33192 12368
rect 36636 12223 36688 12232
rect 36636 12189 36645 12223
rect 36645 12189 36679 12223
rect 36679 12189 36688 12223
rect 36636 12180 36688 12189
rect 37832 12223 37884 12232
rect 37832 12189 37841 12223
rect 37841 12189 37875 12223
rect 37875 12189 37884 12223
rect 37832 12180 37884 12189
rect 27804 12112 27856 12121
rect 14556 12087 14608 12096
rect 14556 12053 14565 12087
rect 14565 12053 14599 12087
rect 14599 12053 14608 12087
rect 14556 12044 14608 12053
rect 23112 12087 23164 12096
rect 23112 12053 23121 12087
rect 23121 12053 23155 12087
rect 23155 12053 23164 12087
rect 23112 12044 23164 12053
rect 28724 12087 28776 12096
rect 28724 12053 28733 12087
rect 28733 12053 28767 12087
rect 28767 12053 28776 12087
rect 28724 12044 28776 12053
rect 34704 12044 34756 12096
rect 37832 12044 37884 12096
rect 38016 12087 38068 12096
rect 38016 12053 38025 12087
rect 38025 12053 38059 12087
rect 38059 12053 38068 12087
rect 38016 12044 38068 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2136 11883 2188 11892
rect 2136 11849 2145 11883
rect 2145 11849 2179 11883
rect 2179 11849 2188 11883
rect 2136 11840 2188 11849
rect 24216 11883 24268 11892
rect 24216 11849 24225 11883
rect 24225 11849 24259 11883
rect 24259 11849 24268 11883
rect 24216 11840 24268 11849
rect 32588 11883 32640 11892
rect 32588 11849 32597 11883
rect 32597 11849 32631 11883
rect 32631 11849 32640 11883
rect 32588 11840 32640 11849
rect 15384 11704 15436 11756
rect 24308 11704 24360 11756
rect 28724 11704 28776 11756
rect 23388 11636 23440 11688
rect 36636 11636 36688 11688
rect 1676 11568 1728 11620
rect 23112 11568 23164 11620
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 17960 11500 18012 11552
rect 38016 11543 38068 11552
rect 38016 11509 38025 11543
rect 38025 11509 38059 11543
rect 38059 11509 38068 11543
rect 38016 11500 38068 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 36636 11296 36688 11348
rect 23388 11271 23440 11280
rect 23388 11237 23397 11271
rect 23397 11237 23431 11271
rect 23431 11237 23440 11271
rect 23388 11228 23440 11237
rect 35348 11228 35400 11280
rect 38016 11271 38068 11280
rect 38016 11237 38025 11271
rect 38025 11237 38059 11271
rect 38059 11237 38068 11271
rect 38016 11228 38068 11237
rect 2780 11092 2832 11144
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 8300 11092 8352 11144
rect 8760 11092 8812 11144
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 19432 11092 19484 11144
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 28448 11135 28500 11144
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 2044 11067 2096 11076
rect 2044 11033 2053 11067
rect 2053 11033 2087 11067
rect 2087 11033 2096 11067
rect 2044 11024 2096 11033
rect 23572 11067 23624 11076
rect 23572 11033 23581 11067
rect 23581 11033 23615 11067
rect 23615 11033 23624 11067
rect 23572 11024 23624 11033
rect 27712 11067 27764 11076
rect 27712 11033 27721 11067
rect 27721 11033 27755 11067
rect 27755 11033 27764 11067
rect 28448 11101 28457 11135
rect 28457 11101 28491 11135
rect 28491 11101 28500 11135
rect 28448 11092 28500 11101
rect 37004 11160 37056 11212
rect 34520 11092 34572 11144
rect 34704 11135 34756 11144
rect 34704 11101 34713 11135
rect 34713 11101 34747 11135
rect 34747 11101 34756 11135
rect 34704 11092 34756 11101
rect 37372 11135 37424 11144
rect 37372 11101 37381 11135
rect 37381 11101 37415 11135
rect 37415 11101 37424 11135
rect 37372 11092 37424 11101
rect 37832 11135 37884 11144
rect 37832 11101 37841 11135
rect 37841 11101 37875 11135
rect 37875 11101 37884 11135
rect 37832 11092 37884 11101
rect 27712 11024 27764 11033
rect 10324 10999 10376 11008
rect 10324 10965 10333 10999
rect 10333 10965 10367 10999
rect 10367 10965 10376 10999
rect 10324 10956 10376 10965
rect 18328 10956 18380 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1860 10752 1912 10804
rect 15660 10752 15712 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 23572 10752 23624 10804
rect 12256 10616 12308 10668
rect 14832 10616 14884 10668
rect 19340 10684 19392 10736
rect 18328 10659 18380 10668
rect 18328 10625 18362 10659
rect 18362 10625 18380 10659
rect 18328 10616 18380 10625
rect 24308 10616 24360 10668
rect 34520 10616 34572 10668
rect 37188 10616 37240 10668
rect 36360 10548 36412 10600
rect 12348 10480 12400 10532
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 37740 10412 37792 10464
rect 38016 10455 38068 10464
rect 38016 10421 38025 10455
rect 38025 10421 38059 10455
rect 38059 10421 38068 10455
rect 38016 10412 38068 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 8024 10208 8076 10260
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 12348 10208 12400 10260
rect 4068 10072 4120 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 10324 10072 10376 10124
rect 11704 10140 11756 10192
rect 18052 10208 18104 10260
rect 36360 10251 36412 10260
rect 36360 10217 36369 10251
rect 36369 10217 36403 10251
rect 36403 10217 36412 10251
rect 36360 10208 36412 10217
rect 37188 10251 37240 10260
rect 37188 10217 37197 10251
rect 37197 10217 37231 10251
rect 37231 10217 37240 10251
rect 37188 10208 37240 10217
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 14832 10115 14884 10124
rect 14832 10081 14841 10115
rect 14841 10081 14875 10115
rect 14875 10081 14884 10115
rect 14832 10072 14884 10081
rect 17960 10072 18012 10124
rect 36176 10072 36228 10124
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 36544 10047 36596 10056
rect 36544 10013 36553 10047
rect 36553 10013 36587 10047
rect 36587 10013 36596 10047
rect 36544 10004 36596 10013
rect 37004 10047 37056 10056
rect 37004 10013 37013 10047
rect 37013 10013 37047 10047
rect 37047 10013 37056 10047
rect 37004 10004 37056 10013
rect 37096 10004 37148 10056
rect 1860 9936 1912 9945
rect 12532 9936 12584 9988
rect 15200 9936 15252 9988
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 5540 9868 5592 9920
rect 7932 9868 7984 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 16212 9911 16264 9920
rect 16212 9877 16221 9911
rect 16221 9877 16255 9911
rect 16255 9877 16264 9911
rect 16212 9868 16264 9877
rect 19432 9936 19484 9988
rect 23204 9979 23256 9988
rect 23204 9945 23213 9979
rect 23213 9945 23247 9979
rect 23247 9945 23256 9979
rect 23204 9936 23256 9945
rect 29828 9936 29880 9988
rect 38108 9868 38160 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 16212 9664 16264 9716
rect 5540 9596 5592 9648
rect 23204 9596 23256 9648
rect 27620 9596 27672 9648
rect 28908 9596 28960 9648
rect 30104 9664 30156 9716
rect 37096 9664 37148 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 3056 9528 3108 9580
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 24308 9571 24360 9580
rect 24308 9537 24317 9571
rect 24317 9537 24351 9571
rect 24351 9537 24360 9571
rect 24308 9528 24360 9537
rect 31024 9528 31076 9580
rect 35348 9596 35400 9648
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 34796 9528 34848 9580
rect 36176 9528 36228 9580
rect 10324 9460 10376 9512
rect 12716 9392 12768 9444
rect 27620 9460 27672 9512
rect 27896 9460 27948 9512
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 34060 9392 34112 9444
rect 38016 9435 38068 9444
rect 38016 9401 38025 9435
rect 38025 9401 38059 9435
rect 38059 9401 38068 9435
rect 38016 9392 38068 9401
rect 36636 9324 36688 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 4068 9120 4120 9172
rect 5172 9095 5224 9104
rect 5172 9061 5181 9095
rect 5181 9061 5215 9095
rect 5215 9061 5224 9095
rect 5172 9052 5224 9061
rect 2688 8916 2740 8968
rect 2872 8891 2924 8900
rect 2872 8857 2881 8891
rect 2881 8857 2915 8891
rect 2915 8857 2924 8891
rect 2872 8848 2924 8857
rect 3424 8848 3476 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 31024 9052 31076 9104
rect 32312 8984 32364 9036
rect 34796 8916 34848 8968
rect 36636 8959 36688 8968
rect 36636 8925 36645 8959
rect 36645 8925 36679 8959
rect 36679 8925 36688 8959
rect 36636 8916 36688 8925
rect 37372 8916 37424 8968
rect 33784 8848 33836 8900
rect 2780 8780 2832 8789
rect 8300 8780 8352 8832
rect 37832 8780 37884 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 2872 8576 2924 8628
rect 5172 8576 5224 8628
rect 33784 8619 33836 8628
rect 33784 8585 33793 8619
rect 33793 8585 33827 8619
rect 33827 8585 33836 8619
rect 33784 8576 33836 8585
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 27896 8440 27948 8492
rect 34060 8508 34112 8560
rect 37372 8551 37424 8560
rect 37372 8517 37381 8551
rect 37381 8517 37415 8551
rect 37415 8517 37424 8551
rect 37372 8508 37424 8517
rect 37832 8483 37884 8492
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 34796 8372 34848 8424
rect 37004 8372 37056 8424
rect 37832 8304 37884 8356
rect 38016 8347 38068 8356
rect 38016 8313 38025 8347
rect 38025 8313 38059 8347
rect 38059 8313 38068 8347
rect 38016 8304 38068 8313
rect 34704 8279 34756 8288
rect 34704 8245 34713 8279
rect 34713 8245 34747 8279
rect 34747 8245 34756 8279
rect 34704 8236 34756 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2780 8032 2832 8084
rect 19340 7896 19392 7948
rect 19984 7896 20036 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 18604 7828 18656 7880
rect 3424 7760 3476 7812
rect 29828 7871 29880 7880
rect 29828 7837 29837 7871
rect 29837 7837 29871 7871
rect 29871 7837 29880 7871
rect 29828 7828 29880 7837
rect 36820 7828 36872 7880
rect 37004 7871 37056 7880
rect 37004 7837 37013 7871
rect 37013 7837 37047 7871
rect 37047 7837 37056 7871
rect 37004 7828 37056 7837
rect 2228 7735 2280 7744
rect 2228 7701 2237 7735
rect 2237 7701 2271 7735
rect 2271 7701 2280 7735
rect 2228 7692 2280 7701
rect 7380 7692 7432 7744
rect 9680 7692 9732 7744
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 32128 7760 32180 7812
rect 21456 7692 21508 7701
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1860 7488 1912 7540
rect 2228 7488 2280 7540
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 18604 7531 18656 7540
rect 7380 7488 7432 7497
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 19984 7531 20036 7540
rect 19984 7497 19993 7531
rect 19993 7497 20027 7531
rect 20027 7497 20036 7531
rect 19984 7488 20036 7497
rect 2044 7420 2096 7472
rect 2688 7352 2740 7404
rect 8300 7420 8352 7472
rect 8484 7395 8536 7404
rect 8484 7361 8518 7395
rect 8518 7361 8536 7395
rect 8484 7352 8536 7361
rect 21456 7420 21508 7472
rect 15292 7352 15344 7404
rect 32128 7395 32180 7404
rect 32128 7361 32137 7395
rect 32137 7361 32171 7395
rect 32171 7361 32180 7395
rect 32128 7352 32180 7361
rect 32312 7395 32364 7404
rect 32312 7361 32321 7395
rect 32321 7361 32355 7395
rect 32355 7361 32364 7395
rect 32312 7352 32364 7361
rect 34704 7352 34756 7404
rect 37832 7395 37884 7404
rect 37832 7361 37841 7395
rect 37841 7361 37875 7395
rect 37875 7361 37884 7395
rect 37832 7352 37884 7361
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 7932 7284 7984 7336
rect 9588 7284 9640 7336
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 8116 7148 8168 7200
rect 9680 7148 9732 7200
rect 30656 7191 30708 7200
rect 30656 7157 30665 7191
rect 30665 7157 30699 7191
rect 30699 7157 30708 7191
rect 33324 7216 33376 7268
rect 30656 7148 30708 7157
rect 32864 7148 32916 7200
rect 37832 7148 37884 7200
rect 38016 7191 38068 7200
rect 38016 7157 38025 7191
rect 38025 7157 38059 7191
rect 38059 7157 38068 7191
rect 38016 7148 38068 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 7932 6944 7984 6996
rect 8484 6944 8536 6996
rect 9680 6944 9732 6996
rect 30656 6944 30708 6996
rect 36820 6944 36872 6996
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 13268 6740 13320 6792
rect 15108 6740 15160 6792
rect 19340 6808 19392 6860
rect 1860 6715 1912 6724
rect 1860 6681 1869 6715
rect 1869 6681 1903 6715
rect 1903 6681 1912 6715
rect 1860 6672 1912 6681
rect 12072 6672 12124 6724
rect 34060 6808 34112 6860
rect 27896 6783 27948 6792
rect 13820 6604 13872 6656
rect 17224 6604 17276 6656
rect 27896 6749 27905 6783
rect 27905 6749 27939 6783
rect 27939 6749 27948 6783
rect 27896 6740 27948 6749
rect 36544 6740 36596 6792
rect 37372 6783 37424 6792
rect 37372 6749 37381 6783
rect 37381 6749 37415 6783
rect 37415 6749 37424 6783
rect 37372 6740 37424 6749
rect 37832 6783 37884 6792
rect 37832 6749 37841 6783
rect 37841 6749 37875 6783
rect 37875 6749 37884 6783
rect 37832 6740 37884 6749
rect 38016 6647 38068 6656
rect 38016 6613 38025 6647
rect 38025 6613 38059 6647
rect 38059 6613 38068 6647
rect 38016 6604 38068 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2688 6443 2740 6452
rect 2688 6409 2697 6443
rect 2697 6409 2731 6443
rect 2731 6409 2740 6443
rect 2688 6400 2740 6409
rect 7932 6400 7984 6452
rect 13268 6443 13320 6452
rect 3424 6264 3476 6316
rect 2228 6239 2280 6248
rect 2228 6205 2237 6239
rect 2237 6205 2271 6239
rect 2271 6205 2280 6239
rect 2228 6196 2280 6205
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 12072 6332 12124 6384
rect 17224 6332 17276 6384
rect 13820 6264 13872 6316
rect 24584 6307 24636 6316
rect 24584 6273 24618 6307
rect 24618 6273 24636 6307
rect 33324 6307 33376 6316
rect 24584 6264 24636 6273
rect 33324 6273 33333 6307
rect 33333 6273 33367 6307
rect 33367 6273 33376 6307
rect 33324 6264 33376 6273
rect 36544 6307 36596 6316
rect 36544 6273 36553 6307
rect 36553 6273 36587 6307
rect 36587 6273 36596 6307
rect 36544 6264 36596 6273
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 19340 6196 19392 6248
rect 15292 6128 15344 6180
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 25688 6103 25740 6112
rect 25688 6069 25697 6103
rect 25697 6069 25731 6103
rect 25731 6069 25740 6103
rect 25688 6060 25740 6069
rect 37832 6060 37884 6112
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3424 5856 3476 5908
rect 34060 5899 34112 5908
rect 34060 5865 34069 5899
rect 34069 5865 34103 5899
rect 34103 5865 34112 5899
rect 34060 5856 34112 5865
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 29736 5652 29788 5704
rect 34060 5652 34112 5704
rect 34796 5652 34848 5704
rect 37372 5695 37424 5704
rect 37372 5661 37381 5695
rect 37381 5661 37415 5695
rect 37415 5661 37424 5695
rect 37372 5652 37424 5661
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 12808 5584 12860 5636
rect 35072 5559 35124 5568
rect 35072 5525 35081 5559
rect 35081 5525 35115 5559
rect 35115 5525 35124 5559
rect 35072 5516 35124 5525
rect 38016 5559 38068 5568
rect 38016 5525 38025 5559
rect 38025 5525 38059 5559
rect 38059 5525 38068 5559
rect 38016 5516 38068 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2780 5176 2832 5228
rect 35072 5176 35124 5228
rect 27252 5040 27304 5092
rect 5816 4972 5868 5024
rect 38016 5015 38068 5024
rect 38016 4981 38025 5015
rect 38025 4981 38059 5015
rect 38059 4981 38068 5015
rect 38016 4972 38068 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1676 4768 1728 4820
rect 24124 4768 24176 4820
rect 27252 4811 27304 4820
rect 27252 4777 27261 4811
rect 27261 4777 27295 4811
rect 27295 4777 27304 4811
rect 27252 4768 27304 4777
rect 3884 4564 3936 4616
rect 7196 4632 7248 4684
rect 15016 4564 15068 4616
rect 24492 4564 24544 4616
rect 27896 4564 27948 4616
rect 32864 4607 32916 4616
rect 32864 4573 32873 4607
rect 32873 4573 32907 4607
rect 32907 4573 32916 4607
rect 32864 4564 32916 4573
rect 37188 4607 37240 4616
rect 37188 4573 37197 4607
rect 37197 4573 37231 4607
rect 37231 4573 37240 4607
rect 37188 4564 37240 4573
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 1860 4539 1912 4548
rect 1860 4505 1869 4539
rect 1869 4505 1903 4539
rect 1903 4505 1912 4539
rect 1860 4496 1912 4505
rect 5816 4539 5868 4548
rect 5816 4505 5825 4539
rect 5825 4505 5859 4539
rect 5859 4505 5868 4539
rect 5816 4496 5868 4505
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 5080 4428 5132 4480
rect 5724 4471 5776 4480
rect 5724 4437 5733 4471
rect 5733 4437 5767 4471
rect 5767 4437 5776 4471
rect 6644 4471 6696 4480
rect 5724 4428 5776 4437
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 24768 4539 24820 4548
rect 24768 4505 24777 4539
rect 24777 4505 24811 4539
rect 24811 4505 24820 4539
rect 24768 4496 24820 4505
rect 28172 4471 28224 4480
rect 23756 4428 23808 4437
rect 28172 4437 28181 4471
rect 28181 4437 28215 4471
rect 28215 4437 28224 4471
rect 28172 4428 28224 4437
rect 34520 4428 34572 4480
rect 36084 4428 36136 4480
rect 36360 4428 36412 4480
rect 38016 4471 38068 4480
rect 38016 4437 38025 4471
rect 38025 4437 38059 4471
rect 38059 4437 38068 4471
rect 38016 4428 38068 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 7196 4224 7248 4276
rect 28172 4224 28224 4276
rect 4896 4088 4948 4140
rect 11428 4088 11480 4140
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 1860 3884 1912 3936
rect 15568 4020 15620 4072
rect 17960 4088 18012 4140
rect 19340 4088 19392 4140
rect 20536 4131 20588 4140
rect 20536 4097 20554 4131
rect 20554 4097 20588 4131
rect 20536 4088 20588 4097
rect 7564 3952 7616 4004
rect 14556 3952 14608 4004
rect 15200 3952 15252 4004
rect 19616 3952 19668 4004
rect 4620 3884 4672 3936
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 20812 3884 20864 3936
rect 21364 3884 21416 3936
rect 22008 3884 22060 3936
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 24768 4156 24820 4208
rect 24124 4088 24176 4140
rect 24492 4088 24544 4140
rect 25688 4088 25740 4140
rect 29736 4088 29788 4140
rect 24584 3995 24636 4004
rect 24584 3961 24593 3995
rect 24593 3961 24627 3995
rect 24627 3961 24636 3995
rect 24584 3952 24636 3961
rect 29736 3952 29788 4004
rect 29920 3995 29972 4004
rect 29920 3961 29929 3995
rect 29929 3961 29963 3995
rect 29963 3961 29972 3995
rect 29920 3952 29972 3961
rect 32864 4020 32916 4072
rect 33600 4131 33652 4140
rect 33600 4097 33609 4131
rect 33609 4097 33643 4131
rect 33643 4097 33652 4131
rect 34796 4156 34848 4208
rect 33600 4088 33652 4097
rect 35808 4088 35860 4140
rect 36084 4131 36136 4140
rect 36084 4097 36093 4131
rect 36093 4097 36127 4131
rect 36127 4097 36136 4131
rect 36084 4088 36136 4097
rect 34520 4020 34572 4072
rect 37832 3952 37884 4004
rect 23204 3884 23256 3936
rect 31024 3884 31076 3936
rect 32864 3927 32916 3936
rect 32864 3893 32873 3927
rect 32873 3893 32907 3927
rect 32907 3893 32916 3927
rect 32864 3884 32916 3893
rect 35532 3884 35584 3936
rect 38016 3927 38068 3936
rect 38016 3893 38025 3927
rect 38025 3893 38059 3927
rect 38059 3893 38068 3927
rect 38016 3884 38068 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4896 3723 4948 3732
rect 4896 3689 4905 3723
rect 4905 3689 4939 3723
rect 4939 3689 4948 3723
rect 4896 3680 4948 3689
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 19616 3723 19668 3732
rect 15108 3680 15160 3689
rect 4620 3612 4672 3664
rect 15568 3655 15620 3664
rect 15568 3621 15577 3655
rect 15577 3621 15611 3655
rect 15611 3621 15620 3655
rect 15568 3612 15620 3621
rect 7564 3544 7616 3596
rect 2964 3519 3016 3528
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 3884 3476 3936 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 7196 3476 7248 3528
rect 8208 3476 8260 3528
rect 9588 3544 9640 3596
rect 19616 3689 19625 3723
rect 19625 3689 19659 3723
rect 19659 3689 19668 3723
rect 19616 3680 19668 3689
rect 20536 3680 20588 3732
rect 24124 3680 24176 3732
rect 37832 3680 37884 3732
rect 23204 3612 23256 3664
rect 3424 3408 3476 3460
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 16672 3519 16724 3528
rect 16672 3485 16690 3519
rect 16690 3485 16724 3519
rect 16672 3476 16724 3485
rect 11428 3408 11480 3460
rect 35808 3612 35860 3664
rect 36544 3612 36596 3664
rect 37188 3612 37240 3664
rect 19616 3476 19668 3528
rect 20812 3476 20864 3528
rect 21824 3476 21876 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 27160 3476 27212 3528
rect 27896 3519 27948 3528
rect 27896 3485 27905 3519
rect 27905 3485 27939 3519
rect 27939 3485 27948 3519
rect 27896 3476 27948 3485
rect 29736 3476 29788 3528
rect 33048 3476 33100 3528
rect 10508 3340 10560 3392
rect 33600 3476 33652 3528
rect 35532 3519 35584 3528
rect 35532 3485 35541 3519
rect 35541 3485 35575 3519
rect 35575 3485 35584 3519
rect 35532 3476 35584 3485
rect 36452 3519 36504 3528
rect 36452 3485 36461 3519
rect 36461 3485 36495 3519
rect 36495 3485 36504 3519
rect 36452 3476 36504 3485
rect 27160 3383 27212 3392
rect 27160 3349 27169 3383
rect 27169 3349 27203 3383
rect 27203 3349 27212 3383
rect 27160 3340 27212 3349
rect 28080 3383 28132 3392
rect 28080 3349 28089 3383
rect 28089 3349 28123 3383
rect 28123 3349 28132 3383
rect 28080 3340 28132 3349
rect 37280 3383 37332 3392
rect 37280 3349 37289 3383
rect 37289 3349 37323 3383
rect 37323 3349 37332 3383
rect 37280 3340 37332 3349
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3792 3136 3844 3188
rect 6644 3136 6696 3188
rect 1860 3111 1912 3120
rect 1860 3077 1869 3111
rect 1869 3077 1903 3111
rect 1903 3077 1912 3111
rect 1860 3068 1912 3077
rect 8944 3068 8996 3120
rect 9404 3136 9456 3188
rect 10508 3136 10560 3188
rect 11060 3136 11112 3188
rect 28080 3136 28132 3188
rect 36452 3136 36504 3188
rect 32864 3068 32916 3120
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 8208 3000 8260 3052
rect 17960 3000 18012 3052
rect 24492 3000 24544 3052
rect 31024 3000 31076 3052
rect 35624 3000 35676 3052
rect 1952 2932 2004 2984
rect 27160 2932 27212 2984
rect 23756 2864 23808 2916
rect 24584 2864 24636 2916
rect 37740 3000 37792 3052
rect 2780 2796 2832 2848
rect 3424 2839 3476 2848
rect 3424 2805 3433 2839
rect 3433 2805 3467 2839
rect 3467 2805 3476 2839
rect 3424 2796 3476 2805
rect 3976 2796 4028 2848
rect 4988 2839 5040 2848
rect 4988 2805 4997 2839
rect 4997 2805 5031 2839
rect 5031 2805 5040 2839
rect 4988 2796 5040 2805
rect 8944 2796 8996 2848
rect 15568 2796 15620 2848
rect 34796 2839 34848 2848
rect 34796 2805 34805 2839
rect 34805 2805 34839 2839
rect 34839 2805 34848 2839
rect 34796 2796 34848 2805
rect 38108 2796 38160 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2964 2592 3016 2644
rect 3884 2592 3936 2644
rect 33048 2592 33100 2644
rect 3056 2456 3108 2508
rect 35716 2524 35768 2576
rect 22008 2456 22060 2508
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4068 2388 4120 2440
rect 4988 2388 5040 2440
rect 34796 2388 34848 2440
rect 35256 2431 35308 2440
rect 35256 2397 35265 2431
rect 35265 2397 35299 2431
rect 35299 2397 35308 2431
rect 35256 2388 35308 2397
rect 36360 2388 36412 2440
rect 36544 2388 36596 2440
rect 37832 2431 37884 2440
rect 37832 2397 37841 2431
rect 37841 2397 37875 2431
rect 37875 2397 37884 2431
rect 37832 2388 37884 2397
rect 15200 2320 15252 2372
rect 2872 2252 2924 2304
rect 35808 2295 35860 2304
rect 35808 2261 35817 2295
rect 35817 2261 35851 2295
rect 35851 2261 35860 2295
rect 35808 2252 35860 2261
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3148 1300 3200 1352
rect 14464 1300 14516 1352
<< metal2 >>
rect 3790 39808 3846 39817
rect 3790 39743 3846 39752
rect 2962 38992 3018 39001
rect 2962 38927 3018 38936
rect 2594 38584 2650 38593
rect 2594 38519 2650 38528
rect 1766 37768 1822 37777
rect 1766 37703 1822 37712
rect 1780 37126 1808 37703
rect 2608 37466 2636 38519
rect 2596 37460 2648 37466
rect 2596 37402 2648 37408
rect 2044 37324 2096 37330
rect 2044 37266 2096 37272
rect 1860 37256 1912 37262
rect 1860 37198 1912 37204
rect 1768 37120 1820 37126
rect 1768 37062 1820 37068
rect 1780 36854 1808 37062
rect 1872 36961 1900 37198
rect 1858 36952 1914 36961
rect 1858 36887 1914 36896
rect 1768 36848 1820 36854
rect 1768 36790 1820 36796
rect 2056 36281 2084 37266
rect 2134 37224 2190 37233
rect 2608 37194 2636 37402
rect 2134 37159 2190 37168
rect 2596 37188 2648 37194
rect 2148 36310 2176 37159
rect 2596 37130 2648 37136
rect 2872 36848 2924 36854
rect 2872 36790 2924 36796
rect 2780 36576 2832 36582
rect 2778 36544 2780 36553
rect 2832 36544 2834 36553
rect 2778 36479 2834 36488
rect 2136 36304 2188 36310
rect 2042 36272 2098 36281
rect 2136 36246 2188 36252
rect 2042 36207 2098 36216
rect 2780 36168 2832 36174
rect 1858 36136 1914 36145
rect 2780 36110 2832 36116
rect 1858 36071 1860 36080
rect 1912 36071 1914 36080
rect 1860 36042 1912 36048
rect 2596 36032 2648 36038
rect 2596 35974 2648 35980
rect 2608 35737 2636 35974
rect 2594 35728 2650 35737
rect 2594 35663 2650 35672
rect 2792 35290 2820 36110
rect 2884 36106 2912 36790
rect 2872 36100 2924 36106
rect 2872 36042 2924 36048
rect 2976 35834 3004 38927
rect 3330 37360 3386 37369
rect 3330 37295 3386 37304
rect 3700 37324 3752 37330
rect 3344 36922 3372 37295
rect 3700 37266 3752 37272
rect 3332 36916 3384 36922
rect 3332 36858 3384 36864
rect 3332 36780 3384 36786
rect 3332 36722 3384 36728
rect 3516 36780 3568 36786
rect 3516 36722 3568 36728
rect 3344 36378 3372 36722
rect 3332 36372 3384 36378
rect 3332 36314 3384 36320
rect 3528 35834 3556 36722
rect 2964 35828 3016 35834
rect 2964 35770 3016 35776
rect 3516 35828 3568 35834
rect 3516 35770 3568 35776
rect 3056 35692 3108 35698
rect 3056 35634 3108 35640
rect 3068 35329 3096 35634
rect 3712 35630 3740 37266
rect 3804 36582 3832 39743
rect 34518 39672 34574 39681
rect 34518 39607 34574 39616
rect 3882 39400 3938 39409
rect 3882 39335 3938 39344
rect 3896 37398 3924 39335
rect 3974 38176 4030 38185
rect 3974 38111 4030 38120
rect 3884 37392 3936 37398
rect 3884 37334 3936 37340
rect 3896 37262 3924 37334
rect 3884 37256 3936 37262
rect 3884 37198 3936 37204
rect 3988 37126 4016 38111
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4620 37256 4672 37262
rect 33876 37256 33928 37262
rect 4620 37198 4672 37204
rect 29734 37224 29790 37233
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 3896 36922 3924 37062
rect 3884 36916 3936 36922
rect 3884 36858 3936 36864
rect 3976 36780 4028 36786
rect 3976 36722 4028 36728
rect 3792 36576 3844 36582
rect 3792 36518 3844 36524
rect 3700 35624 3752 35630
rect 3700 35566 3752 35572
rect 3054 35320 3110 35329
rect 2780 35284 2832 35290
rect 3988 35290 4016 36722
rect 4080 36650 4108 37130
rect 4068 36644 4120 36650
rect 4068 36586 4120 36592
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4160 36032 4212 36038
rect 4160 35974 4212 35980
rect 4172 35834 4200 35974
rect 4632 35834 4660 37198
rect 26792 37188 26844 37194
rect 33876 37198 33928 37204
rect 29734 37159 29790 37168
rect 26792 37130 26844 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 22468 36848 22520 36854
rect 22468 36790 22520 36796
rect 5170 36544 5226 36553
rect 5170 36479 5226 36488
rect 5184 36378 5212 36479
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 22480 36174 22508 36790
rect 24308 36712 24360 36718
rect 24308 36654 24360 36660
rect 24320 36310 24348 36654
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 25504 36576 25556 36582
rect 25504 36518 25556 36524
rect 24308 36304 24360 36310
rect 24308 36246 24360 36252
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20536 36032 20588 36038
rect 20536 35974 20588 35980
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 4160 35828 4212 35834
rect 4160 35770 4212 35776
rect 4620 35828 4672 35834
rect 4620 35770 4672 35776
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 3054 35255 3110 35264
rect 3976 35284 4028 35290
rect 2780 35226 2832 35232
rect 2688 35080 2740 35086
rect 2688 35022 2740 35028
rect 1492 34944 1544 34950
rect 2228 34944 2280 34950
rect 1492 34886 1544 34892
rect 2226 34912 2228 34921
rect 2280 34912 2282 34921
rect 1504 34105 1532 34886
rect 2226 34847 2282 34856
rect 2700 34746 2728 35022
rect 2688 34740 2740 34746
rect 2688 34682 2740 34688
rect 1860 34604 1912 34610
rect 1860 34546 1912 34552
rect 1872 34513 1900 34546
rect 1858 34504 1914 34513
rect 1914 34462 1992 34490
rect 1858 34439 1914 34448
rect 1490 34096 1546 34105
rect 1490 34031 1546 34040
rect 1860 33924 1912 33930
rect 1860 33866 1912 33872
rect 1872 33697 1900 33866
rect 1858 33688 1914 33697
rect 1964 33658 1992 34462
rect 3068 34202 3096 35255
rect 3976 35226 4028 35232
rect 20456 35086 20484 35974
rect 20548 35698 20576 35974
rect 21468 35834 21496 36110
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21928 35834 21956 36042
rect 21456 35828 21508 35834
rect 21456 35770 21508 35776
rect 21916 35828 21968 35834
rect 21916 35770 21968 35776
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 3976 35012 4028 35018
rect 3976 34954 4028 34960
rect 3988 34746 4016 34954
rect 4620 34944 4672 34950
rect 4620 34886 4672 34892
rect 3976 34740 4028 34746
rect 3976 34682 4028 34688
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 3056 34196 3108 34202
rect 3056 34138 3108 34144
rect 4632 33862 4660 34886
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 4620 33856 4672 33862
rect 4620 33798 4672 33804
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 1858 33623 1914 33632
rect 1952 33652 2004 33658
rect 1952 33594 2004 33600
rect 2688 33516 2740 33522
rect 2688 33458 2740 33464
rect 1492 33312 1544 33318
rect 1490 33280 1492 33289
rect 1544 33280 1546 33289
rect 1490 33215 1546 33224
rect 1858 32872 1914 32881
rect 1858 32807 1860 32816
rect 1912 32807 1914 32816
rect 1860 32778 1912 32784
rect 1872 32502 1900 32778
rect 1952 32768 2004 32774
rect 1952 32710 2004 32716
rect 1964 32570 1992 32710
rect 1952 32564 2004 32570
rect 1952 32506 2004 32512
rect 1860 32496 1912 32502
rect 1860 32438 1912 32444
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1492 32224 1544 32230
rect 1492 32166 1544 32172
rect 1504 32065 1532 32166
rect 1490 32056 1546 32065
rect 1490 31991 1546 32000
rect 1688 31958 1716 32370
rect 2700 32298 2728 33458
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 2792 32473 2820 32846
rect 6184 32768 6236 32774
rect 6184 32710 6236 32716
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 3516 32360 3568 32366
rect 3516 32302 3568 32308
rect 2688 32292 2740 32298
rect 2688 32234 2740 32240
rect 3528 32026 3556 32302
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 1676 31952 1728 31958
rect 1676 31894 1728 31900
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1872 31657 1900 31758
rect 1858 31648 1914 31657
rect 1858 31583 1914 31592
rect 2136 31340 2188 31346
rect 2136 31282 2188 31288
rect 2148 31249 2176 31282
rect 6196 31278 6224 32710
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 7656 31816 7708 31822
rect 7656 31758 7708 31764
rect 11980 31816 12032 31822
rect 11980 31758 12032 31764
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 7288 31680 7340 31686
rect 7288 31622 7340 31628
rect 6184 31272 6236 31278
rect 2134 31240 2190 31249
rect 6184 31214 6236 31220
rect 2134 31175 2190 31184
rect 1492 31136 1544 31142
rect 1492 31078 1544 31084
rect 1504 30841 1532 31078
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 1490 30832 1546 30841
rect 1490 30767 1546 30776
rect 7300 30734 7328 31622
rect 7668 31482 7696 31758
rect 11888 31680 11940 31686
rect 11888 31622 11940 31628
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 11900 31346 11928 31622
rect 7748 31340 7800 31346
rect 7748 31282 7800 31288
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 1860 30660 1912 30666
rect 1860 30602 1912 30608
rect 1872 30433 1900 30602
rect 7760 30598 7788 31282
rect 8024 31272 8076 31278
rect 8024 31214 8076 31220
rect 9036 31272 9088 31278
rect 9036 31214 9088 31220
rect 1952 30592 2004 30598
rect 1952 30534 2004 30540
rect 7748 30592 7800 30598
rect 7748 30534 7800 30540
rect 1858 30424 1914 30433
rect 1858 30359 1914 30368
rect 1964 30122 1992 30534
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 1952 30116 2004 30122
rect 1952 30058 2004 30064
rect 2240 30025 2268 30126
rect 3332 30048 3384 30054
rect 2226 30016 2282 30025
rect 3332 29990 3384 29996
rect 2226 29951 2282 29960
rect 3344 29850 3372 29990
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 3332 29844 3384 29850
rect 3332 29786 3384 29792
rect 3344 29646 3372 29786
rect 3332 29640 3384 29646
rect 2778 29608 2834 29617
rect 1860 29572 1912 29578
rect 3332 29582 3384 29588
rect 2778 29543 2834 29552
rect 1860 29514 1912 29520
rect 1872 29238 1900 29514
rect 2792 29510 2820 29543
rect 2780 29504 2832 29510
rect 2780 29446 2832 29452
rect 1860 29232 1912 29238
rect 1858 29200 1860 29209
rect 1912 29200 1914 29209
rect 1858 29135 1914 29144
rect 1872 29109 1900 29135
rect 2228 29096 2280 29102
rect 2228 29038 2280 29044
rect 2240 28801 2268 29038
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 2226 28792 2282 28801
rect 4214 28784 4522 28804
rect 2226 28727 2282 28736
rect 1492 28416 1544 28422
rect 1490 28384 1492 28393
rect 1860 28416 1912 28422
rect 1544 28384 1546 28393
rect 1860 28358 1912 28364
rect 1490 28319 1546 28328
rect 1872 28082 1900 28358
rect 1860 28076 1912 28082
rect 1860 28018 1912 28024
rect 2780 28076 2832 28082
rect 2780 28018 2832 28024
rect 1872 27985 1900 28018
rect 1858 27976 1914 27985
rect 1858 27911 1914 27920
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2700 27674 2728 27814
rect 2688 27668 2740 27674
rect 2688 27610 2740 27616
rect 2792 27577 2820 28018
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 2778 27568 2834 27577
rect 2778 27503 2834 27512
rect 7104 27396 7156 27402
rect 7104 27338 7156 27344
rect 1492 27328 1544 27334
rect 1492 27270 1544 27276
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 1504 27169 1532 27270
rect 1490 27160 1546 27169
rect 1490 27095 1546 27104
rect 1858 26888 1914 26897
rect 1858 26823 1914 26832
rect 1872 26790 1900 26823
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1872 26382 1900 26726
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1964 25974 1992 27270
rect 2228 26920 2280 26926
rect 2228 26862 2280 26868
rect 2240 26489 2268 26862
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 7116 26586 7144 27338
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 2780 26512 2832 26518
rect 2226 26480 2282 26489
rect 2780 26454 2832 26460
rect 2226 26415 2282 26424
rect 2792 26081 2820 26454
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 3896 25974 3924 26318
rect 1952 25968 2004 25974
rect 1952 25910 2004 25916
rect 3792 25968 3844 25974
rect 3792 25910 3844 25916
rect 3884 25968 3936 25974
rect 3884 25910 3936 25916
rect 1964 25673 1992 25910
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 1950 25664 2006 25673
rect 1950 25599 2006 25608
rect 2976 25498 3004 25842
rect 3804 25498 3832 25910
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 3792 25492 3844 25498
rect 3792 25434 3844 25440
rect 2136 25288 2188 25294
rect 2134 25256 2136 25265
rect 2188 25256 2190 25265
rect 2134 25191 2190 25200
rect 2688 25220 2740 25226
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1504 24857 1532 25094
rect 2148 24954 2176 25191
rect 2688 25162 2740 25168
rect 2136 24948 2188 24954
rect 2136 24890 2188 24896
rect 1490 24848 1546 24857
rect 1490 24783 1546 24792
rect 1860 24812 1912 24818
rect 1860 24754 1912 24760
rect 1872 24449 1900 24754
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1858 24440 1914 24449
rect 1964 24410 1992 24550
rect 1858 24375 1914 24384
rect 1952 24404 2004 24410
rect 1952 24346 2004 24352
rect 2700 24206 2728 25162
rect 4080 25158 4108 25638
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 6932 25498 6960 26318
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 5552 24342 5580 25094
rect 5540 24336 5592 24342
rect 5540 24278 5592 24284
rect 5644 24274 5672 25094
rect 7392 24614 7420 25298
rect 8036 24818 8064 31214
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8496 30870 8524 31078
rect 9048 30938 9076 31214
rect 11992 30938 12020 31758
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16868 31482 16896 31690
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 9036 30932 9088 30938
rect 9036 30874 9088 30880
rect 11980 30932 12032 30938
rect 11980 30874 12032 30880
rect 8484 30864 8536 30870
rect 8484 30806 8536 30812
rect 9048 27606 9076 30874
rect 12360 30802 12388 31350
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 12992 31204 13044 31210
rect 12992 31146 13044 31152
rect 12348 30796 12400 30802
rect 12348 30738 12400 30744
rect 13004 30734 13032 31146
rect 16500 30870 16528 31282
rect 16488 30864 16540 30870
rect 16488 30806 16540 30812
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 16028 30592 16080 30598
rect 16028 30534 16080 30540
rect 16040 30258 16068 30534
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 16132 28626 16160 30738
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 16316 28626 16344 29106
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 16120 28620 16172 28626
rect 16120 28562 16172 28568
rect 16304 28620 16356 28626
rect 16304 28562 16356 28568
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 8300 27464 8352 27470
rect 8300 27406 8352 27412
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 8312 26246 8340 27406
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8312 25702 8340 26182
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 1412 24041 1440 24142
rect 1398 24032 1454 24041
rect 1398 23967 1454 23976
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1490 23624 1546 23633
rect 1490 23559 1546 23568
rect 1504 23322 1532 23559
rect 1492 23316 1544 23322
rect 1492 23258 1544 23264
rect 1872 23225 1900 23666
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 3160 23322 3188 23462
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 3148 23316 3200 23322
rect 3148 23258 3200 23264
rect 1858 23216 1914 23225
rect 7392 23186 7420 24550
rect 8036 24070 8064 24754
rect 8024 24064 8076 24070
rect 8024 24006 8076 24012
rect 1858 23151 1914 23160
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 2136 23112 2188 23118
rect 2136 23054 2188 23060
rect 2148 22817 2176 23054
rect 2134 22808 2190 22817
rect 2134 22743 2190 22752
rect 1492 22432 1544 22438
rect 1490 22400 1492 22409
rect 1860 22432 1912 22438
rect 1544 22400 1546 22409
rect 1860 22374 1912 22380
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 1490 22335 1546 22344
rect 1872 22030 1900 22374
rect 1860 22024 1912 22030
rect 1858 21992 1860 22001
rect 2780 22024 2832 22030
rect 1912 21992 1914 22001
rect 2780 21966 2832 21972
rect 1858 21927 1914 21936
rect 2792 21593 2820 21966
rect 3896 21690 3924 22374
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 2778 21584 2834 21593
rect 2778 21519 2834 21528
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 1492 21344 1544 21350
rect 1492 21286 1544 21292
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1504 21185 1532 21286
rect 1490 21176 1546 21185
rect 1490 21111 1546 21120
rect 1872 20874 1900 21286
rect 2976 21146 3004 21490
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 3896 21078 3924 21626
rect 3884 21072 3936 21078
rect 3884 21014 3936 21020
rect 3988 21010 4016 21830
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4632 21146 4660 21286
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4632 20942 4660 21082
rect 7392 21010 7420 23122
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 2044 20868 2096 20874
rect 2044 20810 2096 20816
rect 1872 20777 1900 20810
rect 1858 20768 1914 20777
rect 1858 20703 1914 20712
rect 2056 20534 2084 20810
rect 7024 20602 7052 20878
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 2044 20528 2096 20534
rect 2044 20470 2096 20476
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2148 20369 2176 20402
rect 2134 20360 2190 20369
rect 2134 20295 2190 20304
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1504 19961 1532 20198
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 1490 19952 1546 19961
rect 1490 19887 1546 19896
rect 7208 19854 7236 20742
rect 7392 20398 7420 20946
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7484 19854 7512 20402
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1872 19553 1900 19722
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1858 19544 1914 19553
rect 1858 19479 1914 19488
rect 1964 19242 1992 19654
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 1952 19236 2004 19242
rect 1952 19178 2004 19184
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 1490 18728 1546 18737
rect 1490 18663 1546 18672
rect 1860 18692 1912 18698
rect 1504 18426 1532 18663
rect 1860 18634 1912 18640
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1872 18329 1900 18634
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18426 1992 18566
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2148 17921 2176 18226
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 2134 17912 2190 17921
rect 4214 17904 4522 17924
rect 2134 17847 2190 17856
rect 1492 17536 1544 17542
rect 1490 17504 1492 17513
rect 2228 17536 2280 17542
rect 1544 17504 1546 17513
rect 2228 17478 2280 17484
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 1490 17439 1546 17448
rect 2240 17134 2268 17478
rect 2228 17128 2280 17134
rect 2884 17105 2912 17478
rect 8036 17338 8064 24006
rect 8312 23866 8340 25638
rect 8404 25226 8432 27270
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10980 26246 11008 26862
rect 11992 26586 12020 27406
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12084 27062 12112 27270
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 12268 26450 12296 27610
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 13188 26382 13216 26726
rect 16132 26450 16160 28562
rect 17236 28150 17264 28630
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17224 28144 17276 28150
rect 17224 28086 17276 28092
rect 17328 27878 17356 28358
rect 17420 28218 17448 31758
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 30802 18000 31622
rect 19076 30870 19104 31758
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 21008 31346 21036 31622
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21008 31142 21036 31282
rect 20996 31136 21048 31142
rect 20996 31078 21048 31084
rect 19064 30864 19116 30870
rect 19064 30806 19116 30812
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 21008 30598 21036 31078
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 21008 28626 21036 30534
rect 21836 30258 21864 30534
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 16132 25838 16160 26386
rect 16500 26042 16528 26930
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 15844 25832 15896 25838
rect 15844 25774 15896 25780
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 8392 25220 8444 25226
rect 8392 25162 8444 25168
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 24206 15424 24754
rect 15856 24682 15884 25774
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 17052 25294 17080 25638
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17236 24818 17264 25094
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17420 24750 17448 28154
rect 18248 28150 18276 28358
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 21468 27878 21496 28494
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 21560 26234 21588 28494
rect 21468 26206 21588 26234
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19352 24954 19380 25774
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 15844 24676 15896 24682
rect 15844 24618 15896 24624
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8312 23186 8340 23802
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 8312 21690 8340 23122
rect 9508 22778 9536 23122
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 15108 21956 15160 21962
rect 15108 21898 15160 21904
rect 15120 21690 15148 21898
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15212 21706 15240 21830
rect 15212 21690 15332 21706
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15200 21684 15332 21690
rect 15252 21678 15332 21684
rect 15200 21626 15252 21632
rect 8312 20058 8340 21626
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15212 21078 15240 21490
rect 15200 21072 15252 21078
rect 15200 21014 15252 21020
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11716 20058 11744 20198
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19514 11560 19722
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11716 18970 11744 19314
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 12452 18698 12480 19654
rect 12544 19446 12572 20742
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12912 18834 12940 20946
rect 15304 20942 15332 21678
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11900 18154 11928 18566
rect 12452 18222 12480 18634
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11716 17338 11744 17478
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2228 17070 2280 17076
rect 2870 17096 2926 17105
rect 2240 16697 2268 17070
rect 2870 17031 2926 17040
rect 2226 16688 2282 16697
rect 2226 16623 2282 16632
rect 2884 16522 2912 17031
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16289 2820 16390
rect 2778 16280 2834 16289
rect 3068 16250 3096 17138
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 2778 16215 2834 16224
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3804 16114 3832 16390
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 1872 15881 1900 16050
rect 1858 15872 1914 15881
rect 1858 15807 1914 15816
rect 2228 15496 2280 15502
rect 2226 15464 2228 15473
rect 3884 15496 3936 15502
rect 2280 15464 2282 15473
rect 3884 15438 3936 15444
rect 2226 15399 2282 15408
rect 2240 15162 2268 15399
rect 3896 15366 3924 15438
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2792 15065 2820 15302
rect 3896 15094 3924 15302
rect 3884 15088 3936 15094
rect 2778 15056 2834 15065
rect 1860 15020 1912 15026
rect 3884 15030 3936 15036
rect 2778 14991 2834 15000
rect 1860 14962 1912 14968
rect 1872 14657 1900 14962
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1858 14648 1914 14657
rect 1964 14618 1992 14758
rect 1858 14583 1914 14592
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 14249 1440 14350
rect 2688 14272 2740 14278
rect 1398 14240 1454 14249
rect 2688 14214 2740 14220
rect 1398 14175 1454 14184
rect 2700 14006 2728 14214
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1490 13832 1546 13841
rect 1490 13767 1546 13776
rect 1504 13530 1532 13767
rect 1872 13569 1900 13874
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1858 13560 1914 13569
rect 1492 13524 1544 13530
rect 1858 13495 1914 13504
rect 1492 13466 1544 13472
rect 1964 13410 1992 13670
rect 1872 13382 1992 13410
rect 1872 12850 1900 13382
rect 2056 13258 2084 13738
rect 2700 13394 2728 13942
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2148 13161 2176 13262
rect 2134 13152 2190 13161
rect 2134 13087 2190 13096
rect 4080 12986 4108 17206
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4528 16584 4580 16590
rect 4632 16574 4660 16662
rect 4632 16546 4752 16574
rect 4528 16526 4580 16532
rect 4540 15892 4568 16526
rect 4620 15904 4672 15910
rect 4540 15864 4620 15892
rect 4620 15846 4672 15852
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4632 15706 4660 15846
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4724 13530 4752 16546
rect 5092 16454 5120 16934
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5092 14550 5120 16390
rect 6932 15570 6960 17206
rect 8036 17202 8064 17274
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7484 16454 7512 16594
rect 8036 16590 8064 17138
rect 12912 16998 12940 18770
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14476 16998 14504 17546
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 12912 16658 12940 16934
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 15162 7328 15370
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 6932 14074 6960 14962
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 1490 12744 1546 12753
rect 1490 12679 1546 12688
rect 1504 12442 1532 12679
rect 1872 12481 1900 12786
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1858 12472 1914 12481
rect 1492 12436 1544 12442
rect 1858 12407 1914 12416
rect 1492 12378 1544 12384
rect 1676 12232 1728 12238
rect 2056 12209 2084 12650
rect 3160 12442 3188 12786
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 4632 12306 4660 12582
rect 7392 12374 7420 13806
rect 7484 13802 7512 16390
rect 8036 16182 8064 16526
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 2136 12232 2188 12238
rect 1676 12174 1728 12180
rect 2042 12200 2098 12209
rect 1688 11626 1716 12174
rect 4356 12186 4384 12242
rect 2136 12174 2188 12180
rect 2042 12135 2098 12144
rect 2148 11937 2176 12174
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 4080 12158 4384 12186
rect 2134 11928 2190 11937
rect 2134 11863 2136 11872
rect 2188 11863 2190 11872
rect 2136 11834 2188 11840
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1492 11552 1544 11558
rect 1490 11520 1492 11529
rect 1544 11520 1546 11529
rect 1490 11455 1546 11464
rect 2700 11354 2728 12106
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2780 11144 2832 11150
rect 1858 11112 1914 11121
rect 1858 11047 1860 11056
rect 1912 11047 1914 11056
rect 2042 11112 2098 11121
rect 2780 11086 2832 11092
rect 2042 11047 2044 11056
rect 1860 11018 1912 11024
rect 2096 11047 2098 11056
rect 2044 11018 2096 11024
rect 1872 10810 1900 11018
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 2792 10713 2820 11086
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10305 1532 10406
rect 1490 10296 1546 10305
rect 1490 10231 1546 10240
rect 4080 10130 4108 12158
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 7484 10130 7512 13738
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1872 9897 1900 9930
rect 3056 9920 3108 9926
rect 1858 9888 1914 9897
rect 3056 9862 3108 9868
rect 1858 9823 1914 9832
rect 3068 9586 3096 9862
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 1412 9489 1440 9522
rect 1398 9480 1454 9489
rect 1398 9415 1454 9424
rect 2056 9081 2084 9522
rect 3252 9178 3280 9522
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 2042 9072 2098 9081
rect 2042 9007 2098 9016
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8673 1532 8774
rect 1490 8664 1546 8673
rect 2700 8634 2728 8910
rect 3436 8906 3464 9318
rect 4080 9178 4108 10066
rect 7944 9926 7972 15846
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 13870 8340 15302
rect 8956 15162 8984 15438
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 12714 8340 13806
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8956 12434 8984 15098
rect 11716 14278 11744 15438
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 15026 12020 15302
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12912 14482 12940 16594
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14482 13124 14758
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 8772 12406 8984 12434
rect 8772 11558 8800 12406
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 11150 8800 11494
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8036 10266 8064 11086
rect 8312 10470 8340 11086
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 5552 9654 5580 9862
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 1490 8599 1546 8608
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8265 1900 8434
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1400 7880 1452 7886
rect 1398 7848 1400 7857
rect 1452 7848 1454 7857
rect 1398 7783 1454 7792
rect 1872 7546 1900 8191
rect 2792 8090 2820 8774
rect 2884 8634 2912 8842
rect 5184 8634 5212 9046
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 2056 7478 2084 7822
rect 3436 7818 3464 8366
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 2240 7546 2268 7686
rect 7392 7546 7420 7686
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 2044 7472 2096 7478
rect 2042 7440 2044 7449
rect 2096 7440 2098 7449
rect 2042 7375 2098 7384
rect 2688 7404 2740 7410
rect 2056 7349 2084 7375
rect 2688 7346 2740 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 7041 1532 7142
rect 1490 7032 1546 7041
rect 1490 6967 1546 6976
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6633 1900 6666
rect 1858 6624 1914 6633
rect 1858 6559 1914 6568
rect 2700 6458 2728 7346
rect 7944 7342 7972 9862
rect 8312 8838 8340 10406
rect 10336 10130 10364 10950
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10266 12296 10610
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 10266 12388 10474
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10336 9518 10364 10066
rect 11716 9926 11744 10134
rect 12544 9994 12572 10406
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 12728 9450 12756 10066
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 7478 8340 8774
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2228 6248 2280 6254
rect 2134 6216 2190 6225
rect 2228 6190 2280 6196
rect 2134 6151 2190 6160
rect 2148 5710 2176 6151
rect 2240 5817 2268 6190
rect 3436 6118 3464 6258
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5914 3464 6054
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 2226 5808 2282 5817
rect 2226 5743 2282 5752
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1504 5409 1532 5510
rect 1490 5400 1546 5409
rect 1490 5335 1546 5344
rect 1688 4826 1716 5646
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 1872 5001 1900 5170
rect 1858 4992 1914 5001
rect 1858 4927 1914 4936
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 2792 4593 2820 5170
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3884 4616 3936 4622
rect 2778 4584 2834 4593
rect 1860 4548 1912 4554
rect 3884 4558 3936 4564
rect 2778 4519 2834 4528
rect 1860 4490 1912 4496
rect 1872 4185 1900 4490
rect 3896 4486 3924 4558
rect 5828 4554 5856 4966
rect 7208 4690 7236 7278
rect 7944 7002 7972 7278
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7944 6458 7972 6938
rect 8128 6798 8156 7142
rect 8496 7002 8524 7346
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 1858 4176 1914 4185
rect 1858 4111 1914 4120
rect 3896 4049 3924 4422
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 1504 3777 1532 3878
rect 1490 3768 1546 3777
rect 1490 3703 1546 3712
rect 1872 3466 1900 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3670 4660 3878
rect 4908 3738 4936 4082
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 5092 3534 5120 4422
rect 5736 4282 5764 4422
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1872 3369 1900 3402
rect 1952 3392 2004 3398
rect 1858 3360 1914 3369
rect 1952 3334 2004 3340
rect 1858 3295 1914 3304
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1872 2553 1900 3062
rect 1964 2990 1992 3334
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1858 2544 1914 2553
rect 1858 2479 1914 2488
rect 2792 1737 2820 2790
rect 2976 2650 3004 3470
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3252 2961 3280 2994
rect 3238 2952 3294 2961
rect 3238 2887 3294 2896
rect 3436 2854 3464 3402
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3194 3832 3334
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3896 2650 3924 3470
rect 6656 3194 6684 4422
rect 7208 4282 7236 4626
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7208 3534 7236 4218
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7576 3602 7604 3946
rect 9600 3602 9628 7278
rect 9692 7206 9720 7686
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 7002 9720 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12084 6390 12112 6666
rect 13280 6458 13308 6734
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6458 13860 6598
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 13832 6322 13860 6394
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5642 12848 6190
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 8220 3058 8248 3470
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 9416 3194 9444 3334
rect 10520 3194 10548 3334
rect 11072 3194 11100 3470
rect 11440 3466 11468 4082
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8956 2854 8984 3062
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2778 1728 2834 1737
rect 2778 1663 2834 1672
rect 2884 241 2912 2246
rect 3068 1329 3096 2450
rect 3988 2446 4016 2790
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5000 2446 5028 2790
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 3148 1352 3200 1358
rect 3054 1320 3110 1329
rect 3148 1294 3200 1300
rect 3054 1255 3110 1264
rect 3160 513 3188 1294
rect 3988 921 4016 2382
rect 4080 2145 4108 2382
rect 4066 2136 4122 2145
rect 4066 2071 4122 2080
rect 14476 1358 14504 16934
rect 15396 12986 15424 24142
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15672 20942 15700 23666
rect 17144 21894 17172 24550
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 21468 23050 21496 26206
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 21100 22234 21128 22918
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 21100 22030 21128 22170
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20602 15700 20878
rect 17144 20806 17172 21830
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20364 21146 20392 21422
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20548 20942 20576 21626
rect 20628 21548 20680 21554
rect 20732 21536 20760 21830
rect 20680 21508 20760 21536
rect 20628 21490 20680 21496
rect 20732 20942 20760 21508
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15672 17882 15700 20538
rect 17144 18766 17172 20742
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 20732 20466 20760 20878
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20548 19854 20576 20334
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 20916 19310 20944 20198
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 17882 16712 18226
rect 16868 18154 16896 18634
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12102 14596 12786
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 4010 14596 12038
rect 15396 11762 15424 12922
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15672 10810 15700 17818
rect 17972 17746 18000 18566
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 21100 18290 21128 20402
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 16224 16658 16252 17682
rect 21100 17678 21128 18226
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17270 17172 17478
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 16794 21404 16934
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 15570 16252 16594
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17328 15026 17356 15302
rect 19260 15042 19288 15370
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 17316 15020 17368 15026
rect 19260 15014 19472 15042
rect 17316 14962 17368 14968
rect 19444 14958 19472 15014
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 14278 19380 14758
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21376 14346 21404 14554
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 10130 14872 10610
rect 17972 10130 18000 11494
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10266 18092 11086
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10674 18368 10950
rect 19352 10742 19380 14214
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 21376 12782 21404 13806
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10810 19472 11086
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15212 9874 15240 9930
rect 15028 9846 15240 9874
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 15028 4622 15056 9846
rect 16224 9722 16252 9862
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 15120 3738 15148 6734
rect 15304 6186 15332 7346
rect 17972 7342 18000 10066
rect 19352 7954 19380 10678
rect 19444 9994 19472 10746
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18616 7546 18644 7822
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6390 17264 6598
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 17972 4146 18000 7278
rect 19352 6866 19380 7890
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19996 7546 20024 7890
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6254 19380 6802
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19352 4146 19380 6190
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15212 2378 15240 3946
rect 15580 3670 15608 4014
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15580 2854 15608 3606
rect 16684 3534 16712 3878
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 17972 3058 18000 4082
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19628 3738 19656 3946
rect 20548 3738 20576 4082
rect 21376 3942 21404 12718
rect 21468 11150 21496 22986
rect 21928 21690 21956 35770
rect 24780 35698 24808 36518
rect 25516 36174 25544 36518
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 25516 35630 25544 36110
rect 25976 35834 26004 36110
rect 26804 36038 26832 37130
rect 29748 36922 29776 37159
rect 29826 36952 29882 36961
rect 29736 36916 29788 36922
rect 29826 36887 29882 36896
rect 29736 36858 29788 36864
rect 29748 36242 29776 36858
rect 29736 36236 29788 36242
rect 29736 36178 29788 36184
rect 29840 36106 29868 36887
rect 30748 36576 30800 36582
rect 30748 36518 30800 36524
rect 30288 36372 30340 36378
rect 30288 36314 30340 36320
rect 30012 36168 30064 36174
rect 30300 36145 30328 36314
rect 30760 36281 30788 36518
rect 30746 36272 30802 36281
rect 30746 36207 30802 36216
rect 30760 36174 30788 36207
rect 30748 36168 30800 36174
rect 30012 36110 30064 36116
rect 30286 36136 30342 36145
rect 29828 36100 29880 36106
rect 29828 36042 29880 36048
rect 26792 36032 26844 36038
rect 26792 35974 26844 35980
rect 25964 35828 26016 35834
rect 25964 35770 26016 35776
rect 30024 35698 30052 36110
rect 30748 36110 30800 36116
rect 30286 36071 30342 36080
rect 33888 35834 33916 37198
rect 34532 37126 34560 39607
rect 37370 39264 37426 39273
rect 37370 39199 37426 39208
rect 35530 38856 35586 38865
rect 35530 38791 35586 38800
rect 35346 38040 35402 38049
rect 35346 37975 35402 37984
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35072 37256 35124 37262
rect 35072 37198 35124 37204
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 35084 36961 35112 37198
rect 35360 37126 35388 37975
rect 35440 37188 35492 37194
rect 35440 37130 35492 37136
rect 35348 37120 35400 37126
rect 35348 37062 35400 37068
rect 35070 36952 35126 36961
rect 35070 36887 35126 36896
rect 34702 36816 34758 36825
rect 34702 36751 34704 36760
rect 34756 36751 34758 36760
rect 34796 36780 34848 36786
rect 34704 36722 34756 36728
rect 34796 36722 34848 36728
rect 34808 36310 34836 36722
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34796 36304 34848 36310
rect 34796 36246 34848 36252
rect 34518 36136 34574 36145
rect 34518 36071 34520 36080
rect 34572 36071 34574 36080
rect 34520 36042 34572 36048
rect 35452 36038 35480 37130
rect 35544 36922 35572 38791
rect 37278 38448 37334 38457
rect 37278 38383 37334 38392
rect 37186 37632 37242 37641
rect 37186 37567 37242 37576
rect 37200 37330 37228 37567
rect 37188 37324 37240 37330
rect 37188 37266 37240 37272
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35806 37224 35862 37233
rect 35532 36916 35584 36922
rect 35532 36858 35584 36864
rect 35728 36378 35756 37198
rect 35806 37159 35862 37168
rect 35820 37126 35848 37159
rect 35808 37120 35860 37126
rect 35808 37062 35860 37068
rect 36636 37120 36688 37126
rect 36636 37062 36688 37068
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35900 36576 35952 36582
rect 35900 36518 35952 36524
rect 35716 36372 35768 36378
rect 35716 36314 35768 36320
rect 35532 36168 35584 36174
rect 35532 36110 35584 36116
rect 35440 36032 35492 36038
rect 35544 36009 35572 36110
rect 35440 35974 35492 35980
rect 35530 36000 35586 36009
rect 35530 35935 35586 35944
rect 35544 35834 35572 35935
rect 33876 35828 33928 35834
rect 33876 35770 33928 35776
rect 35532 35828 35584 35834
rect 35532 35770 35584 35776
rect 35912 35766 35940 36518
rect 36004 36174 36032 36722
rect 36174 36680 36230 36689
rect 36174 36615 36230 36624
rect 36188 36378 36216 36615
rect 36648 36417 36676 37062
rect 36634 36408 36690 36417
rect 36176 36372 36228 36378
rect 37200 36378 37228 37266
rect 37292 36786 37320 38383
rect 37280 36780 37332 36786
rect 37280 36722 37332 36728
rect 36634 36343 36690 36352
rect 37188 36372 37240 36378
rect 36176 36314 36228 36320
rect 37188 36314 37240 36320
rect 35992 36168 36044 36174
rect 35992 36110 36044 36116
rect 36360 36168 36412 36174
rect 36360 36110 36412 36116
rect 35900 35760 35952 35766
rect 35900 35702 35952 35708
rect 36372 35698 36400 36110
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 36360 35692 36412 35698
rect 36360 35634 36412 35640
rect 25504 35624 25556 35630
rect 25504 35566 25556 35572
rect 25516 35494 25544 35566
rect 25504 35488 25556 35494
rect 25504 35430 25556 35436
rect 25516 34950 25544 35430
rect 25504 34944 25556 34950
rect 25504 34886 25556 34892
rect 25412 32360 25464 32366
rect 25412 32302 25464 32308
rect 25424 31958 25452 32302
rect 25412 31952 25464 31958
rect 25412 31894 25464 31900
rect 25424 31822 25452 31894
rect 25412 31816 25464 31822
rect 25412 31758 25464 31764
rect 23848 26988 23900 26994
rect 23848 26930 23900 26936
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23492 26450 23520 26726
rect 23860 26518 23888 26930
rect 23848 26512 23900 26518
rect 23848 26454 23900 26460
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23388 26308 23440 26314
rect 23388 26250 23440 26256
rect 23400 25838 23428 26250
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23400 25294 23428 25774
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 23400 24818 23428 25230
rect 24872 24818 24900 25230
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22664 24342 22692 24550
rect 22652 24336 22704 24342
rect 22652 24278 22704 24284
rect 23400 23118 23428 24754
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22020 22642 22048 22918
rect 23400 22778 23428 23054
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 24964 22642 24992 22918
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25148 22234 25176 22374
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25516 21690 25544 34886
rect 30024 34610 30052 35634
rect 36176 35488 36228 35494
rect 36176 35430 36228 35436
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 36188 35018 36216 35430
rect 36176 35012 36228 35018
rect 36176 34954 36228 34960
rect 30012 34604 30064 34610
rect 30012 34546 30064 34552
rect 29276 33992 29328 33998
rect 29276 33934 29328 33940
rect 29288 33658 29316 33934
rect 29276 33652 29328 33658
rect 29276 33594 29328 33600
rect 30024 33522 30052 34546
rect 36372 34474 36400 35634
rect 36544 35624 36596 35630
rect 36544 35566 36596 35572
rect 36556 35290 36584 35566
rect 37188 35488 37240 35494
rect 37188 35430 37240 35436
rect 36544 35284 36596 35290
rect 36544 35226 36596 35232
rect 37200 35086 37228 35430
rect 36728 35080 36780 35086
rect 36726 35048 36728 35057
rect 37188 35080 37240 35086
rect 36780 35048 36782 35057
rect 37188 35022 37240 35028
rect 37292 35034 37320 36722
rect 37384 36242 37412 39199
rect 37372 36236 37424 36242
rect 37372 36178 37424 36184
rect 37384 35222 37412 36178
rect 38016 35488 38068 35494
rect 38014 35456 38016 35465
rect 38068 35456 38070 35465
rect 38014 35391 38070 35400
rect 37372 35216 37424 35222
rect 37372 35158 37424 35164
rect 36726 34983 36782 34992
rect 36820 35012 36872 35018
rect 36820 34954 36872 34960
rect 36832 34542 36860 34954
rect 36820 34536 36872 34542
rect 36820 34478 36872 34484
rect 36360 34468 36412 34474
rect 36360 34410 36412 34416
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 36372 33998 36400 34410
rect 37200 34241 37228 35022
rect 37292 35006 37412 35034
rect 37280 34944 37332 34950
rect 37280 34886 37332 34892
rect 37292 34610 37320 34886
rect 37384 34678 37412 35006
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 37372 34672 37424 34678
rect 38028 34649 38056 34886
rect 37372 34614 37424 34620
rect 38014 34640 38070 34649
rect 37280 34604 37332 34610
rect 38014 34575 38070 34584
rect 37280 34546 37332 34552
rect 37186 34232 37242 34241
rect 37186 34167 37242 34176
rect 35348 33992 35400 33998
rect 35348 33934 35400 33940
rect 36360 33992 36412 33998
rect 36360 33934 36412 33940
rect 37372 33992 37424 33998
rect 37372 33934 37424 33940
rect 37832 33992 37884 33998
rect 37832 33934 37884 33940
rect 30012 33516 30064 33522
rect 30012 33458 30064 33464
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26068 32570 26096 32846
rect 30024 32570 30052 33458
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35360 33114 35388 33934
rect 37384 33425 37412 33934
rect 37844 33658 37872 33934
rect 38016 33856 38068 33862
rect 38014 33824 38016 33833
rect 38068 33824 38070 33833
rect 38014 33759 38070 33768
rect 37832 33652 37884 33658
rect 37832 33594 37884 33600
rect 37832 33516 37884 33522
rect 37832 33458 37884 33464
rect 37370 33416 37426 33425
rect 37370 33351 37426 33360
rect 35348 33108 35400 33114
rect 35348 33050 35400 33056
rect 36268 33040 36320 33046
rect 36268 32982 36320 32988
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35820 32774 35848 32846
rect 35808 32768 35860 32774
rect 35808 32710 35860 32716
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 30012 32564 30064 32570
rect 30012 32506 30064 32512
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 26252 31822 26280 32370
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 26252 31482 26280 31758
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 27160 31476 27212 31482
rect 27160 31418 27212 31424
rect 27172 30258 27200 31418
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 27724 31142 27752 31282
rect 28736 31142 28764 32370
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 27712 31136 27764 31142
rect 27712 31078 27764 31084
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 27160 30252 27212 30258
rect 27160 30194 27212 30200
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26344 29306 26372 29582
rect 26332 29300 26384 29306
rect 26332 29242 26384 29248
rect 27172 29170 27200 30194
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 27172 28558 27200 29106
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27908 28082 27936 28358
rect 27896 28076 27948 28082
rect 27896 28018 27948 28024
rect 28736 25294 28764 31078
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35820 30734 35848 32710
rect 35900 31816 35952 31822
rect 35900 31758 35952 31764
rect 35912 31482 35940 31758
rect 35900 31476 35952 31482
rect 35900 31418 35952 31424
rect 36084 31340 36136 31346
rect 36084 31282 36136 31288
rect 36096 30938 36124 31282
rect 36280 31278 36308 32982
rect 37464 32904 37516 32910
rect 37464 32846 37516 32852
rect 37280 32768 37332 32774
rect 37280 32710 37332 32716
rect 37292 32434 37320 32710
rect 37476 32609 37504 32846
rect 37844 32842 37872 33458
rect 38108 33380 38160 33386
rect 38108 33322 38160 33328
rect 38016 33312 38068 33318
rect 38016 33254 38068 33260
rect 38028 33017 38056 33254
rect 38014 33008 38070 33017
rect 38014 32943 38070 32952
rect 38120 32910 38148 33322
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 37832 32836 37884 32842
rect 37832 32778 37884 32784
rect 37462 32600 37518 32609
rect 37462 32535 37518 32544
rect 37280 32428 37332 32434
rect 37280 32370 37332 32376
rect 37648 32428 37700 32434
rect 37648 32370 37700 32376
rect 37280 31952 37332 31958
rect 37280 31894 37332 31900
rect 37292 31793 37320 31894
rect 37278 31784 37334 31793
rect 37278 31719 37334 31728
rect 36268 31272 36320 31278
rect 36268 31214 36320 31220
rect 37660 30938 37688 32370
rect 38014 32192 38070 32201
rect 38014 32127 38070 32136
rect 38028 32026 38056 32127
rect 38016 32020 38068 32026
rect 38016 31962 38068 31968
rect 38120 31385 38148 32846
rect 38106 31376 38162 31385
rect 38106 31311 38162 31320
rect 38016 31136 38068 31142
rect 38016 31078 38068 31084
rect 36084 30932 36136 30938
rect 36084 30874 36136 30880
rect 37648 30932 37700 30938
rect 37648 30874 37700 30880
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 35808 30728 35860 30734
rect 35808 30670 35860 30676
rect 37372 30728 37424 30734
rect 37372 30670 37424 30676
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34796 27396 34848 27402
rect 34796 27338 34848 27344
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31312 26586 31340 26930
rect 34808 26586 34836 27338
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 35256 26376 35308 26382
rect 35256 26318 35308 26324
rect 29656 25906 29684 26318
rect 35268 26042 35296 26318
rect 35256 26036 35308 26042
rect 35256 25978 35308 25984
rect 29644 25900 29696 25906
rect 29644 25842 29696 25848
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 29000 25832 29052 25838
rect 29000 25774 29052 25780
rect 29012 25702 29040 25774
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 29012 25498 29040 25638
rect 29000 25492 29052 25498
rect 29000 25434 29052 25440
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 30024 25158 30052 25842
rect 31484 25696 31536 25702
rect 31484 25638 31536 25644
rect 31496 25294 31524 25638
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 26252 24206 26280 25094
rect 26528 24886 26556 25094
rect 26516 24880 26568 24886
rect 26516 24822 26568 24828
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26436 23730 26464 24006
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26332 22568 26384 22574
rect 26332 22510 26384 22516
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22020 19922 22048 20742
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 17746 22232 18022
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 24320 17678 24348 18566
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 24124 17604 24176 17610
rect 24124 17546 24176 17552
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 16658 22600 17478
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23676 14618 23704 14962
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 7478 21496 7686
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 19628 3534 19656 3674
rect 20824 3534 20852 3878
rect 21836 3534 21864 13806
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11626 23152 12038
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23400 11286 23428 11630
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23584 10810 23612 11018
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23204 9988 23256 9994
rect 23204 9930 23256 9936
rect 23216 9654 23244 9930
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 24136 4826 24164 17546
rect 24320 17338 24348 17614
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24964 15162 24992 21626
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25424 21146 25452 21490
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25596 21072 25648 21078
rect 25596 21014 25648 21020
rect 25608 20806 25636 21014
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25608 20398 25636 20742
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25608 20262 25636 20334
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25608 18630 25636 20198
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 16574 25636 18566
rect 25792 17882 25820 18634
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25976 16574 26004 21626
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26160 20330 26188 20810
rect 26148 20324 26200 20330
rect 26148 20266 26200 20272
rect 26160 18698 26188 20266
rect 26344 18970 26372 22510
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26436 20602 26464 21490
rect 27632 21350 27660 25094
rect 30024 24274 30052 25094
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 29828 23588 29880 23594
rect 29828 23530 29880 23536
rect 29840 23186 29868 23530
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 30024 23118 30052 24210
rect 35360 24206 35388 30670
rect 36176 30660 36228 30666
rect 36176 30602 36228 30608
rect 36188 30326 36216 30602
rect 37188 30592 37240 30598
rect 37188 30534 37240 30540
rect 36176 30320 36228 30326
rect 36176 30262 36228 30268
rect 37200 30258 37228 30534
rect 37188 30252 37240 30258
rect 37188 30194 37240 30200
rect 37280 30184 37332 30190
rect 37280 30126 37332 30132
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 35452 29306 35480 29786
rect 37292 29646 37320 30126
rect 37384 30054 37412 30670
rect 37660 30326 37688 30874
rect 38028 30841 38056 31078
rect 38014 30832 38070 30841
rect 38014 30767 38070 30776
rect 37832 30728 37884 30734
rect 37832 30670 37884 30676
rect 37648 30320 37700 30326
rect 37648 30262 37700 30268
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 37372 30048 37424 30054
rect 37370 30016 37372 30025
rect 37424 30016 37426 30025
rect 37370 29951 37426 29960
rect 37188 29640 37240 29646
rect 37188 29582 37240 29588
rect 37280 29640 37332 29646
rect 37280 29582 37332 29588
rect 35440 29300 35492 29306
rect 35440 29242 35492 29248
rect 37200 28801 37228 29582
rect 37372 29164 37424 29170
rect 37372 29106 37424 29112
rect 37186 28792 37242 28801
rect 37186 28727 37242 28736
rect 37188 28552 37240 28558
rect 37188 28494 37240 28500
rect 35808 28484 35860 28490
rect 35808 28426 35860 28432
rect 35820 28218 35848 28426
rect 35808 28212 35860 28218
rect 35808 28154 35860 28160
rect 37096 27940 37148 27946
rect 37096 27882 37148 27888
rect 37108 27470 37136 27882
rect 37200 27577 37228 28494
rect 37384 28082 37412 29106
rect 37476 29034 37504 30194
rect 37556 29504 37608 29510
rect 37556 29446 37608 29452
rect 37568 29170 37596 29446
rect 37660 29238 37688 30262
rect 37844 30122 37872 30670
rect 38016 30592 38068 30598
rect 38016 30534 38068 30540
rect 38028 30433 38056 30534
rect 38014 30424 38070 30433
rect 38014 30359 38070 30368
rect 37832 30116 37884 30122
rect 37832 30058 37884 30064
rect 38108 30048 38160 30054
rect 38108 29990 38160 29996
rect 38014 29608 38070 29617
rect 38014 29543 38070 29552
rect 38028 29510 38056 29543
rect 38016 29504 38068 29510
rect 38016 29446 38068 29452
rect 37648 29232 37700 29238
rect 38120 29209 38148 29990
rect 37648 29174 37700 29180
rect 38106 29200 38162 29209
rect 37556 29164 37608 29170
rect 38106 29135 38162 29144
rect 37556 29106 37608 29112
rect 37464 29028 37516 29034
rect 37464 28970 37516 28976
rect 37556 28416 37608 28422
rect 38016 28416 38068 28422
rect 37556 28358 37608 28364
rect 38014 28384 38016 28393
rect 38068 28384 38070 28393
rect 37568 28082 37596 28358
rect 38014 28319 38070 28328
rect 37372 28076 37424 28082
rect 37372 28018 37424 28024
rect 37556 28076 37608 28082
rect 37556 28018 37608 28024
rect 37278 27976 37334 27985
rect 37278 27911 37334 27920
rect 37292 27606 37320 27911
rect 37280 27600 37332 27606
rect 37186 27568 37242 27577
rect 37280 27542 37332 27548
rect 37186 27503 37242 27512
rect 37096 27464 37148 27470
rect 37096 27406 37148 27412
rect 37832 27464 37884 27470
rect 37832 27406 37884 27412
rect 37844 26790 37872 27406
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 38028 27169 38056 27270
rect 38014 27160 38070 27169
rect 38014 27095 38070 27104
rect 37832 26784 37884 26790
rect 37832 26726 37884 26732
rect 38016 26784 38068 26790
rect 38016 26726 38068 26732
rect 38028 26625 38056 26726
rect 38014 26616 38070 26625
rect 38014 26551 38070 26560
rect 38108 26376 38160 26382
rect 38108 26318 38160 26324
rect 37740 26240 37792 26246
rect 38120 26217 38148 26318
rect 37740 26182 37792 26188
rect 38106 26208 38162 26217
rect 37752 25906 37780 26182
rect 38106 26143 38162 26152
rect 35440 25900 35492 25906
rect 35440 25842 35492 25848
rect 36452 25900 36504 25906
rect 37740 25900 37792 25906
rect 36504 25860 36584 25888
rect 36452 25842 36504 25848
rect 35452 25498 35480 25842
rect 35440 25492 35492 25498
rect 35440 25434 35492 25440
rect 36556 25294 36584 25860
rect 37740 25842 37792 25848
rect 38014 25800 38070 25809
rect 38014 25735 38016 25744
rect 38068 25735 38070 25744
rect 38016 25706 38068 25712
rect 38016 25424 38068 25430
rect 38014 25392 38016 25401
rect 38068 25392 38070 25401
rect 38014 25327 38070 25336
rect 36544 25288 36596 25294
rect 36544 25230 36596 25236
rect 37372 25288 37424 25294
rect 37372 25230 37424 25236
rect 36556 24206 36584 25230
rect 37384 24993 37412 25230
rect 37370 24984 37426 24993
rect 37370 24919 37372 24928
rect 37424 24919 37426 24928
rect 37372 24890 37424 24896
rect 38016 24608 38068 24614
rect 38014 24576 38016 24585
rect 38068 24576 38070 24585
rect 38014 24511 38070 24520
rect 35348 24200 35400 24206
rect 35348 24142 35400 24148
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 38014 24168 38070 24177
rect 35360 23526 35388 24142
rect 35900 24064 35952 24070
rect 35900 24006 35952 24012
rect 35348 23520 35400 23526
rect 35348 23462 35400 23468
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 30024 22642 30052 23054
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29564 22438 29592 22510
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 29564 22098 29592 22374
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 30484 22030 30512 22374
rect 34532 22234 34560 22578
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34520 22228 34572 22234
rect 34520 22170 34572 22176
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 25608 16546 25728 16574
rect 25976 16546 26188 16574
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24320 14414 24348 14758
rect 24780 14414 24808 14826
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24320 13326 24348 14350
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24412 13530 24440 13874
rect 24872 13870 24900 14350
rect 24964 14006 24992 15098
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24308 13320 24360 13326
rect 24308 13262 24360 13268
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 24228 11898 24256 12106
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24320 11762 24348 13262
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24320 10674 24348 11698
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24320 9586 24348 10610
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23216 3942 23244 4082
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 22020 2514 22048 3878
rect 23216 3670 23244 3878
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 23768 2922 23796 4422
rect 24504 4146 24532 4558
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24136 3738 24164 4082
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24504 3058 24532 4082
rect 24596 4010 24624 6258
rect 25700 6118 25728 16546
rect 26160 14618 26188 16546
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 26160 14414 26188 14554
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26896 12850 26924 18906
rect 27632 18290 27660 21286
rect 28460 21146 28488 21490
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 30116 19446 30144 21286
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30104 19440 30156 19446
rect 30104 19382 30156 19388
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 28908 18284 28960 18290
rect 28908 18226 28960 18232
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 28000 14074 28028 14282
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 28460 13326 28488 14214
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 26884 12844 26936 12850
rect 26884 12786 26936 12792
rect 26896 12442 26924 12786
rect 26884 12436 26936 12442
rect 26884 12378 26936 12384
rect 28460 12238 28488 13262
rect 28632 13184 28684 13190
rect 28632 13126 28684 13132
rect 28644 12986 28672 13126
rect 28632 12980 28684 12986
rect 28632 12922 28684 12928
rect 28448 12232 28500 12238
rect 27802 12200 27858 12209
rect 28448 12174 28500 12180
rect 27802 12135 27804 12144
rect 27856 12135 27858 12144
rect 27804 12106 27856 12112
rect 28460 11150 28488 12174
rect 28724 12096 28776 12102
rect 28724 12038 28776 12044
rect 28736 11762 28764 12038
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28448 11144 28500 11150
rect 27710 11112 27766 11121
rect 28448 11086 28500 11092
rect 27710 11047 27712 11056
rect 27764 11047 27766 11056
rect 27712 11018 27764 11024
rect 28460 10062 28488 11086
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28920 9654 28948 18226
rect 29460 18148 29512 18154
rect 29460 18090 29512 18096
rect 29472 17202 29500 18090
rect 29748 17882 29776 18226
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29196 16114 29224 17138
rect 29644 16992 29696 16998
rect 29644 16934 29696 16940
rect 29656 16590 29684 16934
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 29184 16108 29236 16114
rect 29184 16050 29236 16056
rect 30116 10062 30144 19382
rect 30208 19378 30236 19654
rect 30300 19378 30328 20402
rect 32600 19514 32628 20402
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30300 18358 30328 19314
rect 34532 18834 34560 19790
rect 35360 19446 35388 23462
rect 35912 23186 35940 24006
rect 37384 23798 37412 24142
rect 38014 24103 38070 24112
rect 38028 24070 38056 24103
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 37372 23792 37424 23798
rect 37370 23760 37372 23769
rect 37424 23760 37426 23769
rect 37370 23695 37426 23704
rect 38016 23520 38068 23526
rect 38016 23462 38068 23468
rect 38028 23361 38056 23462
rect 38014 23352 38070 23361
rect 38014 23287 38070 23296
rect 35900 23180 35952 23186
rect 35900 23122 35952 23128
rect 35912 22030 35940 23122
rect 37372 23112 37424 23118
rect 37372 23054 37424 23060
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 37292 22098 37320 22578
rect 37384 22574 37412 23054
rect 38016 22976 38068 22982
rect 38014 22944 38016 22953
rect 38068 22944 38070 22953
rect 38014 22879 38070 22888
rect 37372 22568 37424 22574
rect 37370 22536 37372 22545
rect 37424 22536 37426 22545
rect 37370 22471 37426 22480
rect 38108 22432 38160 22438
rect 38108 22374 38160 22380
rect 37280 22092 37332 22098
rect 37280 22034 37332 22040
rect 35900 22024 35952 22030
rect 35900 21966 35952 21972
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 38014 21992 38070 22001
rect 36096 21894 36124 21966
rect 36084 21888 36136 21894
rect 36084 21830 36136 21836
rect 37384 21185 37412 21966
rect 38014 21927 38070 21936
rect 38028 21894 38056 21927
rect 38016 21888 38068 21894
rect 38016 21830 38068 21836
rect 38120 21593 38148 22374
rect 38106 21584 38162 21593
rect 37832 21548 37884 21554
rect 38106 21519 38162 21528
rect 37832 21490 37884 21496
rect 37464 21480 37516 21486
rect 37464 21422 37516 21428
rect 37370 21176 37426 21185
rect 37370 21111 37426 21120
rect 37476 20942 37504 21422
rect 36912 20936 36964 20942
rect 36912 20878 36964 20884
rect 37096 20936 37148 20942
rect 37096 20878 37148 20884
rect 37464 20936 37516 20942
rect 37464 20878 37516 20884
rect 36924 20058 36952 20878
rect 36912 20052 36964 20058
rect 36912 19994 36964 20000
rect 37108 19961 37136 20878
rect 37280 20800 37332 20806
rect 37280 20742 37332 20748
rect 37188 20256 37240 20262
rect 37188 20198 37240 20204
rect 37094 19952 37150 19961
rect 37094 19887 37150 19896
rect 36268 19848 36320 19854
rect 36268 19790 36320 19796
rect 36280 19514 36308 19790
rect 36544 19780 36596 19786
rect 36544 19722 36596 19728
rect 36556 19514 36584 19722
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 36544 19508 36596 19514
rect 36544 19450 36596 19456
rect 35348 19440 35400 19446
rect 35348 19382 35400 19388
rect 36280 19378 36308 19450
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 30288 18352 30340 18358
rect 30288 18294 30340 18300
rect 30300 18154 30328 18294
rect 36280 18290 36308 19314
rect 37200 19145 37228 20198
rect 37292 19922 37320 20742
rect 37844 20602 37872 21490
rect 38108 21344 38160 21350
rect 38108 21286 38160 21292
rect 38016 20800 38068 20806
rect 38014 20768 38016 20777
rect 38068 20768 38070 20777
rect 38014 20703 38070 20712
rect 37832 20596 37884 20602
rect 37832 20538 37884 20544
rect 38120 20369 38148 21286
rect 38106 20360 38162 20369
rect 38106 20295 38162 20304
rect 37280 19916 37332 19922
rect 37280 19858 37332 19864
rect 38016 19712 38068 19718
rect 38016 19654 38068 19660
rect 38028 19553 38056 19654
rect 38014 19544 38070 19553
rect 38014 19479 38070 19488
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37186 19136 37242 19145
rect 37186 19071 37242 19080
rect 37384 18970 37412 19246
rect 37372 18964 37424 18970
rect 37372 18906 37424 18912
rect 37188 18760 37240 18766
rect 37186 18728 37188 18737
rect 37240 18728 37242 18737
rect 37186 18663 37242 18672
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 38028 18329 38056 18566
rect 38014 18320 38070 18329
rect 36268 18284 36320 18290
rect 38014 18255 38070 18264
rect 36268 18226 36320 18232
rect 30288 18148 30340 18154
rect 30288 18090 30340 18096
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 36096 16794 36124 17138
rect 36084 16788 36136 16794
rect 36084 16730 36136 16736
rect 36280 16590 36308 18226
rect 37924 18216 37976 18222
rect 37924 18158 37976 18164
rect 37936 17882 37964 18158
rect 38016 18080 38068 18086
rect 38016 18022 38068 18028
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 38028 17785 38056 18022
rect 38014 17776 38070 17785
rect 38014 17711 38070 17720
rect 36820 17672 36872 17678
rect 36820 17614 36872 17620
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 36832 17202 36860 17614
rect 38120 17377 38148 17614
rect 38106 17368 38162 17377
rect 38106 17303 38162 17312
rect 36820 17196 36872 17202
rect 36820 17138 36872 17144
rect 37372 16992 37424 16998
rect 38016 16992 38068 16998
rect 37372 16934 37424 16940
rect 38014 16960 38016 16969
rect 38068 16960 38070 16969
rect 37384 16590 37412 16934
rect 38014 16895 38070 16904
rect 37832 16788 37884 16794
rect 37832 16730 37884 16736
rect 36268 16584 36320 16590
rect 36268 16526 36320 16532
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 36280 16182 36308 16526
rect 36268 16176 36320 16182
rect 37384 16153 37412 16526
rect 36268 16118 36320 16124
rect 37370 16144 37426 16153
rect 37370 16079 37426 16088
rect 36084 16040 36136 16046
rect 36084 15982 36136 15988
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30576 15502 30604 15846
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 36096 15162 36124 15982
rect 36176 15904 36228 15910
rect 36176 15846 36228 15852
rect 36188 15706 36216 15846
rect 36176 15700 36228 15706
rect 36176 15642 36228 15648
rect 37844 15502 37872 16730
rect 38014 16552 38070 16561
rect 38014 16487 38070 16496
rect 38028 16454 38056 16487
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 38014 15736 38070 15745
rect 38014 15671 38016 15680
rect 38068 15671 38070 15680
rect 38016 15642 38068 15648
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 36268 15360 36320 15366
rect 37280 15360 37332 15366
rect 36268 15302 36320 15308
rect 37278 15328 37280 15337
rect 37332 15328 37334 15337
rect 36084 15156 36136 15162
rect 36084 15098 36136 15104
rect 36280 15026 36308 15302
rect 37278 15263 37334 15272
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 36268 15020 36320 15026
rect 36268 14962 36320 14968
rect 32496 14476 32548 14482
rect 32496 14418 32548 14424
rect 32508 14074 32536 14418
rect 33244 14414 33272 14962
rect 36280 14929 36308 14962
rect 36266 14920 36322 14929
rect 36266 14855 36322 14864
rect 36636 14884 36688 14890
rect 36636 14826 36688 14832
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 36648 14618 36676 14826
rect 38016 14816 38068 14822
rect 38016 14758 38068 14764
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 38028 14521 38056 14758
rect 38014 14512 38070 14521
rect 38014 14447 38070 14456
rect 33232 14408 33284 14414
rect 33152 14368 33232 14396
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 33152 13938 33180 14368
rect 33232 14350 33284 14356
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33152 12850 33180 13874
rect 34532 13394 34560 14010
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34520 13388 34572 13394
rect 34520 13330 34572 13336
rect 36280 13326 36308 14214
rect 37200 13705 37228 14350
rect 38016 14272 38068 14278
rect 38016 14214 38068 14220
rect 38028 14113 38056 14214
rect 38014 14104 38070 14113
rect 38014 14039 38070 14048
rect 38108 13932 38160 13938
rect 38108 13874 38160 13880
rect 37832 13728 37884 13734
rect 37186 13696 37242 13705
rect 37832 13670 37884 13676
rect 37186 13631 37242 13640
rect 37844 13326 37872 13670
rect 36084 13320 36136 13326
rect 36084 13262 36136 13268
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 36096 12986 36124 13262
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 37832 13184 37884 13190
rect 38016 13184 38068 13190
rect 37832 13126 37884 13132
rect 38014 13152 38016 13161
rect 38068 13152 38070 13161
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 36280 12850 36308 13126
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 30380 12436 30432 12442
rect 30380 12378 30432 12384
rect 30392 12238 30420 12378
rect 33152 12374 33180 12786
rect 36636 12640 36688 12646
rect 36636 12582 36688 12588
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 33140 12368 33192 12374
rect 33140 12310 33192 12316
rect 32588 12300 32640 12306
rect 32588 12242 32640 12248
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 32312 12232 32364 12238
rect 32312 12174 32364 12180
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 27632 9518 27660 9590
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27908 8498 27936 9454
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27908 6798 27936 8434
rect 29840 7886 29868 9930
rect 30116 9722 30144 9998
rect 30104 9716 30156 9722
rect 30104 9658 30156 9664
rect 32324 9586 32352 12174
rect 32600 11898 32628 12242
rect 36648 12238 36676 12582
rect 37844 12238 37872 13126
rect 38014 13087 38070 13096
rect 38014 12744 38070 12753
rect 38014 12679 38016 12688
rect 38068 12679 38070 12688
rect 38016 12650 38068 12656
rect 38120 12345 38148 13874
rect 38106 12336 38162 12345
rect 38106 12271 38162 12280
rect 36636 12232 36688 12238
rect 36636 12174 36688 12180
rect 37832 12232 37884 12238
rect 37832 12174 37884 12180
rect 34704 12096 34756 12102
rect 34704 12038 34756 12044
rect 37832 12096 37884 12102
rect 37832 12038 37884 12044
rect 38016 12096 38068 12102
rect 38016 12038 38068 12044
rect 32588 11892 32640 11898
rect 32588 11834 32640 11840
rect 34716 11150 34744 12038
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 36648 11354 36676 11630
rect 36636 11348 36688 11354
rect 36636 11290 36688 11296
rect 35348 11280 35400 11286
rect 35348 11222 35400 11228
rect 34520 11144 34572 11150
rect 34520 11086 34572 11092
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 34532 10674 34560 11086
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 35360 9654 35388 11222
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36372 10266 36400 10542
rect 36360 10260 36412 10266
rect 36360 10202 36412 10208
rect 36176 10124 36228 10130
rect 36176 10066 36228 10072
rect 35348 9648 35400 9654
rect 35348 9590 35400 9596
rect 36188 9586 36216 10066
rect 37016 10062 37044 11154
rect 37844 11150 37872 12038
rect 38028 11937 38056 12038
rect 38014 11928 38070 11937
rect 38014 11863 38070 11872
rect 38016 11552 38068 11558
rect 38014 11520 38016 11529
rect 38068 11520 38070 11529
rect 38014 11455 38070 11464
rect 38016 11280 38068 11286
rect 38016 11222 38068 11228
rect 37372 11144 37424 11150
rect 37370 11112 37372 11121
rect 37832 11144 37884 11150
rect 37424 11112 37426 11121
rect 37832 11086 37884 11092
rect 37370 11047 37426 11056
rect 38028 10713 38056 11222
rect 38014 10704 38070 10713
rect 37188 10668 37240 10674
rect 38014 10639 38070 10648
rect 37188 10610 37240 10616
rect 37200 10266 37228 10610
rect 37740 10464 37792 10470
rect 37740 10406 37792 10412
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 37188 10260 37240 10266
rect 37188 10202 37240 10208
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 37004 10056 37056 10062
rect 37004 9998 37056 10004
rect 37096 10056 37148 10062
rect 37096 9998 37148 10004
rect 36556 9897 36584 9998
rect 36542 9888 36598 9897
rect 36542 9823 36598 9832
rect 37108 9722 37136 9998
rect 37096 9716 37148 9722
rect 37096 9658 37148 9664
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 36176 9580 36228 9586
rect 36176 9522 36228 9528
rect 31036 9110 31064 9522
rect 31024 9104 31076 9110
rect 31024 9046 31076 9052
rect 32324 9042 32352 9522
rect 34060 9444 34112 9450
rect 34060 9386 34112 9392
rect 32312 9036 32364 9042
rect 32312 8978 32364 8984
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29840 6914 29868 7822
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 32140 7410 32168 7754
rect 32324 7410 32352 8978
rect 33784 8900 33836 8906
rect 33784 8842 33836 8848
rect 33796 8634 33824 8842
rect 33784 8628 33836 8634
rect 33784 8570 33836 8576
rect 34072 8566 34100 9386
rect 34808 8974 34836 9522
rect 36636 9376 36688 9382
rect 36636 9318 36688 9324
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 36648 8974 36676 9318
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 37372 8968 37424 8974
rect 37372 8910 37424 8916
rect 34060 8560 34112 8566
rect 34060 8502 34112 8508
rect 34808 8430 34836 8910
rect 37384 8566 37412 8910
rect 37372 8560 37424 8566
rect 37370 8528 37372 8537
rect 37424 8528 37426 8537
rect 37370 8463 37426 8472
rect 34796 8424 34848 8430
rect 34796 8366 34848 8372
rect 37004 8424 37056 8430
rect 37004 8366 37056 8372
rect 34704 8288 34756 8294
rect 34704 8230 34756 8236
rect 34716 7410 34744 8230
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 33324 7268 33376 7274
rect 33324 7210 33376 7216
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 32864 7200 32916 7206
rect 32864 7142 32916 7148
rect 30668 7002 30696 7142
rect 30656 6996 30708 7002
rect 30656 6938 30708 6944
rect 29748 6886 29868 6914
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 24768 4548 24820 4554
rect 24768 4490 24820 4496
rect 24780 4214 24808 4490
rect 24768 4208 24820 4214
rect 24768 4150 24820 4156
rect 25700 4146 25728 6054
rect 27252 5092 27304 5098
rect 27252 5034 27304 5040
rect 27264 4826 27292 5034
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 27908 4622 27936 6734
rect 29748 5710 29776 6886
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 24584 4004 24636 4010
rect 24584 3946 24636 3952
rect 27908 3534 27936 4558
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28184 4282 28212 4422
rect 28172 4276 28224 4282
rect 28172 4218 28224 4224
rect 29748 4146 29776 5646
rect 32876 4622 32904 7142
rect 33336 6322 33364 7210
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 34072 5914 34100 6802
rect 34060 5908 34112 5914
rect 34060 5850 34112 5856
rect 34072 5710 34100 5850
rect 34808 5710 34836 8366
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 37016 7886 37044 8366
rect 36820 7880 36872 7886
rect 36820 7822 36872 7828
rect 37004 7880 37056 7886
rect 37004 7822 37056 7828
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 36832 7002 36860 7822
rect 37370 7304 37426 7313
rect 37370 7239 37426 7248
rect 36820 6996 36872 7002
rect 36820 6938 36872 6944
rect 37384 6798 37412 7239
rect 36544 6792 36596 6798
rect 36544 6734 36596 6740
rect 37372 6792 37424 6798
rect 37372 6734 37424 6740
rect 36556 6322 36584 6734
rect 36544 6316 36596 6322
rect 36544 6258 36596 6264
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34796 5704 34848 5710
rect 37372 5704 37424 5710
rect 34796 5646 34848 5652
rect 37370 5672 37372 5681
rect 37424 5672 37426 5681
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 29748 4010 29776 4082
rect 32864 4072 32916 4078
rect 29918 4040 29974 4049
rect 29736 4004 29788 4010
rect 32864 4014 32916 4020
rect 29918 3975 29920 3984
rect 29736 3946 29788 3952
rect 29972 3975 29974 3984
rect 29920 3946 29972 3952
rect 29748 3534 29776 3946
rect 32876 3942 32904 4014
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24596 2922 24624 3470
rect 27172 3398 27200 3470
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 27172 2990 27200 3334
rect 28092 3194 28120 3334
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 31036 3058 31064 3878
rect 32876 3126 32904 3878
rect 33612 3534 33640 4082
rect 34532 4078 34560 4422
rect 34808 4214 34836 5646
rect 37370 5607 37426 5616
rect 35072 5568 35124 5574
rect 35072 5510 35124 5516
rect 35084 5234 35112 5510
rect 35072 5228 35124 5234
rect 35072 5170 35124 5176
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 36084 4480 36136 4486
rect 36084 4422 36136 4428
rect 36360 4480 36412 4486
rect 36360 4422 36412 4428
rect 34796 4208 34848 4214
rect 34796 4150 34848 4156
rect 36096 4146 36124 4422
rect 35808 4140 35860 4146
rect 35808 4082 35860 4088
rect 36084 4140 36136 4146
rect 36084 4082 36136 4088
rect 34520 4072 34572 4078
rect 34520 4014 34572 4020
rect 35532 3936 35584 3942
rect 35532 3878 35584 3884
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35544 3534 35572 3878
rect 35820 3670 35848 4082
rect 36096 3913 36124 4082
rect 36082 3904 36138 3913
rect 36082 3839 36138 3848
rect 35808 3664 35860 3670
rect 35808 3606 35860 3612
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 35532 3528 35584 3534
rect 35532 3470 35584 3476
rect 32864 3120 32916 3126
rect 32864 3062 32916 3068
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 33060 2650 33088 3470
rect 35624 3052 35676 3058
rect 35624 2994 35676 3000
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 33048 2644 33100 2650
rect 33048 2586 33100 2592
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 34808 2446 34836 2790
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 35268 2281 35296 2382
rect 35254 2272 35310 2281
rect 19574 2204 19882 2224
rect 35254 2207 35310 2216
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 3974 912 4030 921
rect 3974 847 4030 856
rect 3146 504 3202 513
rect 3146 439 3202 448
rect 35636 241 35664 2994
rect 35716 2576 35768 2582
rect 35716 2518 35768 2524
rect 35728 649 35756 2518
rect 36372 2446 36400 4422
rect 37200 3670 37228 4558
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 37188 3664 37240 3670
rect 37188 3606 37240 3612
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 36464 3194 36492 3470
rect 36452 3188 36504 3194
rect 36452 3130 36504 3136
rect 36556 2446 36584 3606
rect 37280 3392 37332 3398
rect 37280 3334 37332 3340
rect 37292 2689 37320 3334
rect 37752 3058 37780 10406
rect 38028 10305 38056 10406
rect 38014 10296 38070 10305
rect 38014 10231 38070 10240
rect 38108 9920 38160 9926
rect 38108 9862 38160 9868
rect 38014 9480 38070 9489
rect 38014 9415 38016 9424
rect 38068 9415 38070 9424
rect 38016 9386 38068 9392
rect 38120 8945 38148 9862
rect 38106 8936 38162 8945
rect 38106 8871 38162 8880
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37844 8498 37872 8774
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 37832 8356 37884 8362
rect 37832 8298 37884 8304
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 37844 7410 37872 8298
rect 38028 8129 38056 8298
rect 38014 8120 38070 8129
rect 38014 8055 38070 8064
rect 38016 7744 38068 7750
rect 38014 7712 38016 7721
rect 38068 7712 38070 7721
rect 38014 7647 38070 7656
rect 37832 7404 37884 7410
rect 37832 7346 37884 7352
rect 37832 7200 37884 7206
rect 37832 7142 37884 7148
rect 38016 7200 38068 7206
rect 38016 7142 38068 7148
rect 37844 6798 37872 7142
rect 38028 6905 38056 7142
rect 38014 6896 38070 6905
rect 38014 6831 38070 6840
rect 37832 6792 37884 6798
rect 37832 6734 37884 6740
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38028 6497 38056 6598
rect 38014 6488 38070 6497
rect 38014 6423 38070 6432
rect 37832 6112 37884 6118
rect 38016 6112 38068 6118
rect 37832 6054 37884 6060
rect 38014 6080 38016 6089
rect 38068 6080 38070 6089
rect 37844 5710 37872 6054
rect 38014 6015 38070 6024
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 38028 5273 38056 5510
rect 38014 5264 38070 5273
rect 38014 5199 38070 5208
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 38028 4865 38056 4966
rect 38014 4856 38070 4865
rect 38014 4791 38070 4800
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37844 4010 37872 4558
rect 38016 4480 38068 4486
rect 38016 4422 38068 4428
rect 38028 4321 38056 4422
rect 38014 4312 38070 4321
rect 38014 4247 38070 4256
rect 37832 4004 37884 4010
rect 37832 3946 37884 3952
rect 38016 3936 38068 3942
rect 38016 3878 38068 3884
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 37278 2680 37334 2689
rect 37278 2615 37334 2624
rect 37844 2446 37872 3674
rect 38028 3505 38056 3878
rect 38014 3496 38070 3505
rect 38014 3431 38070 3440
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 38028 3097 38056 3334
rect 38014 3088 38070 3097
rect 38014 3023 38070 3032
rect 38108 2848 38160 2854
rect 38108 2790 38160 2796
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 37832 2440 37884 2446
rect 37832 2382 37884 2388
rect 35808 2304 35860 2310
rect 35808 2246 35860 2252
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 35820 1057 35848 2246
rect 38028 1465 38056 2246
rect 38120 1873 38148 2790
rect 38106 1864 38162 1873
rect 38106 1799 38162 1808
rect 38014 1456 38070 1465
rect 38014 1391 38070 1400
rect 35806 1048 35862 1057
rect 35806 983 35862 992
rect 35714 640 35770 649
rect 35714 575 35770 584
rect 2870 232 2926 241
rect 2870 167 2926 176
rect 35622 232 35678 241
rect 35622 167 35678 176
<< via2 >>
rect 3790 39752 3846 39808
rect 2962 38936 3018 38992
rect 2594 38528 2650 38584
rect 1766 37712 1822 37768
rect 1858 36896 1914 36952
rect 2134 37168 2190 37224
rect 2778 36524 2780 36544
rect 2780 36524 2832 36544
rect 2832 36524 2834 36544
rect 2778 36488 2834 36524
rect 2042 36216 2098 36272
rect 1858 36100 1914 36136
rect 1858 36080 1860 36100
rect 1860 36080 1912 36100
rect 1912 36080 1914 36100
rect 2594 35672 2650 35728
rect 3330 37304 3386 37360
rect 34518 39616 34574 39672
rect 3882 39344 3938 39400
rect 3974 38120 4030 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3054 35264 3110 35320
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 29734 37168 29790 37224
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 5170 36488 5226 36544
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 2226 34892 2228 34912
rect 2228 34892 2280 34912
rect 2280 34892 2282 34912
rect 2226 34856 2282 34892
rect 1858 34448 1914 34504
rect 1490 34040 1546 34096
rect 1858 33632 1914 33688
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 1490 33260 1492 33280
rect 1492 33260 1544 33280
rect 1544 33260 1546 33280
rect 1490 33224 1546 33260
rect 1858 32836 1914 32872
rect 1858 32816 1860 32836
rect 1860 32816 1912 32836
rect 1912 32816 1914 32836
rect 1490 32000 1546 32056
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 2778 32408 2834 32464
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1858 31592 1914 31648
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 2134 31184 2190 31240
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 1490 30776 1546 30832
rect 1858 30368 1914 30424
rect 2226 29960 2282 30016
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 2778 29552 2834 29608
rect 1858 29180 1860 29200
rect 1860 29180 1912 29200
rect 1912 29180 1914 29200
rect 1858 29144 1914 29180
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 2226 28736 2282 28792
rect 1490 28364 1492 28384
rect 1492 28364 1544 28384
rect 1544 28364 1546 28384
rect 1490 28328 1546 28364
rect 1858 27920 1914 27976
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 2778 27512 2834 27568
rect 1490 27104 1546 27160
rect 1858 26832 1914 26888
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2226 26424 2282 26480
rect 2778 26016 2834 26072
rect 1950 25608 2006 25664
rect 2134 25236 2136 25256
rect 2136 25236 2188 25256
rect 2188 25236 2190 25256
rect 2134 25200 2190 25236
rect 1490 24792 1546 24848
rect 1858 24384 1914 24440
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1398 23976 1454 24032
rect 1490 23568 1546 23624
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 1858 23160 1914 23216
rect 2134 22752 2190 22808
rect 1490 22380 1492 22400
rect 1492 22380 1544 22400
rect 1544 22380 1546 22400
rect 1490 22344 1546 22380
rect 1858 21972 1860 21992
rect 1860 21972 1912 21992
rect 1912 21972 1914 21992
rect 1858 21936 1914 21972
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 2778 21528 2834 21584
rect 1490 21120 1546 21176
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1858 20712 1914 20768
rect 2134 20304 2190 20360
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1490 19896 1546 19952
rect 1858 19488 1914 19544
rect 2226 19080 2282 19136
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1490 18672 1546 18728
rect 1858 18264 1914 18320
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 2134 17856 2190 17912
rect 1490 17484 1492 17504
rect 1492 17484 1544 17504
rect 1544 17484 1546 17504
rect 1490 17448 1546 17484
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 2870 17040 2926 17096
rect 2226 16632 2282 16688
rect 2778 16224 2834 16280
rect 1858 15816 1914 15872
rect 2226 15444 2228 15464
rect 2228 15444 2280 15464
rect 2280 15444 2282 15464
rect 2226 15408 2282 15444
rect 2778 15000 2834 15056
rect 1858 14592 1914 14648
rect 1398 14184 1454 14240
rect 1490 13776 1546 13832
rect 1858 13504 1914 13560
rect 2134 13096 2190 13152
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1490 12688 1546 12744
rect 1858 12416 1914 12472
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 2042 12144 2098 12200
rect 2134 11892 2190 11928
rect 2134 11872 2136 11892
rect 2136 11872 2188 11892
rect 2188 11872 2190 11892
rect 1490 11500 1492 11520
rect 1492 11500 1544 11520
rect 1544 11500 1546 11520
rect 1490 11464 1546 11500
rect 1858 11076 1914 11112
rect 1858 11056 1860 11076
rect 1860 11056 1912 11076
rect 1912 11056 1914 11076
rect 2042 11076 2098 11112
rect 2042 11056 2044 11076
rect 2044 11056 2096 11076
rect 2096 11056 2098 11076
rect 2778 10648 2834 10704
rect 1490 10240 1546 10296
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1858 9832 1914 9888
rect 1398 9424 1454 9480
rect 2042 9016 2098 9072
rect 1490 8608 1546 8664
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1858 8200 1914 8256
rect 1398 7828 1400 7848
rect 1400 7828 1452 7848
rect 1452 7828 1454 7848
rect 1398 7792 1454 7828
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 2042 7420 2044 7440
rect 2044 7420 2096 7440
rect 2096 7420 2098 7440
rect 2042 7384 2098 7420
rect 1490 6976 1546 7032
rect 1858 6568 1914 6624
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2134 6160 2190 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 2226 5752 2282 5808
rect 1490 5344 1546 5400
rect 1858 4936 1914 4992
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2778 4528 2834 4584
rect 1858 4120 1914 4176
rect 3882 3984 3938 4040
rect 1490 3712 1546 3768
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1858 3304 1914 3360
rect 1858 2488 1914 2544
rect 3238 2896 3294 2952
rect 2778 1672 2834 1728
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3054 1264 3110 1320
rect 4066 2080 4122 2136
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 29826 36896 29882 36952
rect 30746 36216 30802 36272
rect 30286 36080 30342 36136
rect 37370 39208 37426 39264
rect 35530 38800 35586 38856
rect 35346 37984 35402 38040
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35070 36896 35126 36952
rect 34702 36780 34758 36816
rect 34702 36760 34704 36780
rect 34704 36760 34756 36780
rect 34756 36760 34758 36780
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34518 36100 34574 36136
rect 34518 36080 34520 36100
rect 34520 36080 34572 36100
rect 34572 36080 34574 36100
rect 37278 38392 37334 38448
rect 37186 37576 37242 37632
rect 35806 37168 35862 37224
rect 35530 35944 35586 36000
rect 36174 36624 36230 36680
rect 36634 36352 36690 36408
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 36726 35028 36728 35048
rect 36728 35028 36780 35048
rect 36780 35028 36782 35048
rect 36726 34992 36782 35028
rect 38014 35436 38016 35456
rect 38016 35436 38068 35456
rect 38068 35436 38070 35456
rect 38014 35400 38070 35436
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 38014 34584 38070 34640
rect 37186 34176 37242 34232
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 38014 33804 38016 33824
rect 38016 33804 38068 33824
rect 38068 33804 38070 33824
rect 38014 33768 38070 33804
rect 37370 33360 37426 33416
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 38014 32952 38070 33008
rect 37462 32544 37518 32600
rect 37278 31728 37334 31784
rect 38014 32136 38070 32192
rect 38106 31320 38162 31376
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 38014 30776 38070 30832
rect 37370 29996 37372 30016
rect 37372 29996 37424 30016
rect 37424 29996 37426 30016
rect 37370 29960 37426 29996
rect 37186 28736 37242 28792
rect 38014 30368 38070 30424
rect 38014 29552 38070 29608
rect 38106 29144 38162 29200
rect 38014 28364 38016 28384
rect 38016 28364 38068 28384
rect 38068 28364 38070 28384
rect 38014 28328 38070 28364
rect 37278 27920 37334 27976
rect 37186 27512 37242 27568
rect 38014 27104 38070 27160
rect 38014 26560 38070 26616
rect 38106 26152 38162 26208
rect 38014 25764 38070 25800
rect 38014 25744 38016 25764
rect 38016 25744 38068 25764
rect 38068 25744 38070 25764
rect 38014 25372 38016 25392
rect 38016 25372 38068 25392
rect 38068 25372 38070 25392
rect 38014 25336 38070 25372
rect 37370 24948 37426 24984
rect 37370 24928 37372 24948
rect 37372 24928 37424 24948
rect 37424 24928 37426 24948
rect 38014 24556 38016 24576
rect 38016 24556 38068 24576
rect 38068 24556 38070 24576
rect 38014 24520 38070 24556
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 27802 12164 27858 12200
rect 27802 12144 27804 12164
rect 27804 12144 27856 12164
rect 27856 12144 27858 12164
rect 27710 11076 27766 11112
rect 27710 11056 27712 11076
rect 27712 11056 27764 11076
rect 27764 11056 27766 11076
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 38014 24112 38070 24168
rect 37370 23740 37372 23760
rect 37372 23740 37424 23760
rect 37424 23740 37426 23760
rect 37370 23704 37426 23740
rect 38014 23296 38070 23352
rect 38014 22924 38016 22944
rect 38016 22924 38068 22944
rect 38068 22924 38070 22944
rect 38014 22888 38070 22924
rect 37370 22516 37372 22536
rect 37372 22516 37424 22536
rect 37424 22516 37426 22536
rect 37370 22480 37426 22516
rect 38014 21936 38070 21992
rect 38106 21528 38162 21584
rect 37370 21120 37426 21176
rect 37094 19896 37150 19952
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 38014 20748 38016 20768
rect 38016 20748 38068 20768
rect 38068 20748 38070 20768
rect 38014 20712 38070 20748
rect 38106 20304 38162 20360
rect 38014 19488 38070 19544
rect 37186 19080 37242 19136
rect 37186 18708 37188 18728
rect 37188 18708 37240 18728
rect 37240 18708 37242 18728
rect 37186 18672 37242 18708
rect 38014 18264 38070 18320
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 38014 17720 38070 17776
rect 38106 17312 38162 17368
rect 38014 16940 38016 16960
rect 38016 16940 38068 16960
rect 38068 16940 38070 16960
rect 38014 16904 38070 16940
rect 37370 16088 37426 16144
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38014 16496 38070 16552
rect 38014 15700 38070 15736
rect 38014 15680 38016 15700
rect 38016 15680 38068 15700
rect 38068 15680 38070 15700
rect 37278 15308 37280 15328
rect 37280 15308 37332 15328
rect 37332 15308 37334 15328
rect 37278 15272 37334 15308
rect 36266 14864 36322 14920
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38014 14456 38070 14512
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 38014 14048 38070 14104
rect 37186 13640 37242 13696
rect 38014 13132 38016 13152
rect 38016 13132 38068 13152
rect 38068 13132 38070 13152
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38014 13096 38070 13132
rect 38014 12708 38070 12744
rect 38014 12688 38016 12708
rect 38016 12688 38068 12708
rect 38068 12688 38070 12708
rect 38106 12280 38162 12336
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 38014 11872 38070 11928
rect 38014 11500 38016 11520
rect 38016 11500 38068 11520
rect 38068 11500 38070 11520
rect 38014 11464 38070 11500
rect 37370 11092 37372 11112
rect 37372 11092 37424 11112
rect 37424 11092 37426 11112
rect 37370 11056 37426 11092
rect 38014 10648 38070 10704
rect 36542 9832 36598 9888
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 37370 8508 37372 8528
rect 37372 8508 37424 8528
rect 37424 8508 37426 8528
rect 37370 8472 37426 8508
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37370 7248 37426 7304
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 37370 5652 37372 5672
rect 37372 5652 37424 5672
rect 37424 5652 37426 5672
rect 29918 4004 29974 4040
rect 29918 3984 29920 4004
rect 29920 3984 29972 4004
rect 29972 3984 29974 4004
rect 37370 5616 37426 5652
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36082 3848 36138 3904
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35254 2216 35310 2272
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 3974 856 4030 912
rect 3146 448 3202 504
rect 38014 10240 38070 10296
rect 38014 9444 38070 9480
rect 38014 9424 38016 9444
rect 38016 9424 38068 9444
rect 38068 9424 38070 9444
rect 38106 8880 38162 8936
rect 38014 8064 38070 8120
rect 38014 7692 38016 7712
rect 38016 7692 38068 7712
rect 38068 7692 38070 7712
rect 38014 7656 38070 7692
rect 38014 6840 38070 6896
rect 38014 6432 38070 6488
rect 38014 6060 38016 6080
rect 38016 6060 38068 6080
rect 38068 6060 38070 6080
rect 38014 6024 38070 6060
rect 38014 5208 38070 5264
rect 38014 4800 38070 4856
rect 38014 4256 38070 4312
rect 37278 2624 37334 2680
rect 38014 3440 38070 3496
rect 38014 3032 38070 3088
rect 38106 1808 38162 1864
rect 38014 1400 38070 1456
rect 35806 992 35862 1048
rect 35714 584 35770 640
rect 2870 176 2926 232
rect 35622 176 35678 232
<< metal3 >>
rect 0 39810 800 39840
rect 3785 39810 3851 39813
rect 0 39808 3851 39810
rect 0 39752 3790 39808
rect 3846 39752 3851 39808
rect 0 39750 3851 39752
rect 0 39720 800 39750
rect 3785 39747 3851 39750
rect 34513 39674 34579 39677
rect 39200 39674 40000 39704
rect 34513 39672 40000 39674
rect 34513 39616 34518 39672
rect 34574 39616 40000 39672
rect 34513 39614 40000 39616
rect 34513 39611 34579 39614
rect 39200 39584 40000 39614
rect 0 39402 800 39432
rect 3877 39402 3943 39405
rect 0 39400 3943 39402
rect 0 39344 3882 39400
rect 3938 39344 3943 39400
rect 0 39342 3943 39344
rect 0 39312 800 39342
rect 3877 39339 3943 39342
rect 37365 39266 37431 39269
rect 39200 39266 40000 39296
rect 37365 39264 40000 39266
rect 37365 39208 37370 39264
rect 37426 39208 40000 39264
rect 37365 39206 40000 39208
rect 37365 39203 37431 39206
rect 39200 39176 40000 39206
rect 0 38994 800 39024
rect 2957 38994 3023 38997
rect 0 38992 3023 38994
rect 0 38936 2962 38992
rect 3018 38936 3023 38992
rect 0 38934 3023 38936
rect 0 38904 800 38934
rect 2957 38931 3023 38934
rect 35525 38858 35591 38861
rect 39200 38858 40000 38888
rect 35525 38856 40000 38858
rect 35525 38800 35530 38856
rect 35586 38800 40000 38856
rect 35525 38798 40000 38800
rect 35525 38795 35591 38798
rect 39200 38768 40000 38798
rect 0 38586 800 38616
rect 2589 38586 2655 38589
rect 0 38584 2655 38586
rect 0 38528 2594 38584
rect 2650 38528 2655 38584
rect 0 38526 2655 38528
rect 0 38496 800 38526
rect 2589 38523 2655 38526
rect 37273 38450 37339 38453
rect 39200 38450 40000 38480
rect 37273 38448 40000 38450
rect 37273 38392 37278 38448
rect 37334 38392 40000 38448
rect 37273 38390 40000 38392
rect 37273 38387 37339 38390
rect 39200 38360 40000 38390
rect 0 38178 800 38208
rect 3969 38178 4035 38181
rect 0 38176 4035 38178
rect 0 38120 3974 38176
rect 4030 38120 4035 38176
rect 0 38118 4035 38120
rect 0 38088 800 38118
rect 3969 38115 4035 38118
rect 35341 38042 35407 38045
rect 39200 38042 40000 38072
rect 35341 38040 40000 38042
rect 35341 37984 35346 38040
rect 35402 37984 40000 38040
rect 35341 37982 40000 37984
rect 35341 37979 35407 37982
rect 39200 37952 40000 37982
rect 0 37770 800 37800
rect 1761 37770 1827 37773
rect 0 37768 1827 37770
rect 0 37712 1766 37768
rect 1822 37712 1827 37768
rect 0 37710 1827 37712
rect 0 37680 800 37710
rect 1761 37707 1827 37710
rect 37181 37634 37247 37637
rect 39200 37634 40000 37664
rect 37181 37632 40000 37634
rect 37181 37576 37186 37632
rect 37242 37576 40000 37632
rect 37181 37574 40000 37576
rect 37181 37571 37247 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 39200 37544 40000 37574
rect 34928 37503 35248 37504
rect 0 37362 800 37392
rect 3325 37362 3391 37365
rect 0 37360 3391 37362
rect 0 37304 3330 37360
rect 3386 37304 3391 37360
rect 0 37302 3391 37304
rect 0 37272 800 37302
rect 3325 37299 3391 37302
rect 2129 37226 2195 37229
rect 29729 37226 29795 37229
rect 2129 37224 29795 37226
rect 2129 37168 2134 37224
rect 2190 37168 29734 37224
rect 29790 37168 29795 37224
rect 2129 37166 29795 37168
rect 2129 37163 2195 37166
rect 29729 37163 29795 37166
rect 35801 37226 35867 37229
rect 39200 37226 40000 37256
rect 35801 37224 40000 37226
rect 35801 37168 35806 37224
rect 35862 37168 40000 37224
rect 35801 37166 40000 37168
rect 35801 37163 35867 37166
rect 39200 37136 40000 37166
rect 19568 37024 19888 37025
rect 0 36954 800 36984
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 1853 36954 1919 36957
rect 0 36952 1919 36954
rect 0 36896 1858 36952
rect 1914 36896 1919 36952
rect 0 36894 1919 36896
rect 0 36864 800 36894
rect 1853 36891 1919 36894
rect 29821 36954 29887 36957
rect 35065 36954 35131 36957
rect 29821 36952 35131 36954
rect 29821 36896 29826 36952
rect 29882 36896 35070 36952
rect 35126 36896 35131 36952
rect 29821 36894 35131 36896
rect 29821 36891 29887 36894
rect 35065 36891 35131 36894
rect 34697 36818 34763 36821
rect 39200 36818 40000 36848
rect 34697 36816 40000 36818
rect 34697 36760 34702 36816
rect 34758 36760 40000 36816
rect 34697 36758 40000 36760
rect 34697 36755 34763 36758
rect 39200 36728 40000 36758
rect 36169 36682 36235 36685
rect 26190 36680 36235 36682
rect 26190 36624 36174 36680
rect 36230 36624 36235 36680
rect 26190 36622 36235 36624
rect 0 36546 800 36576
rect 2773 36546 2839 36549
rect 0 36544 2839 36546
rect 0 36488 2778 36544
rect 2834 36488 2839 36544
rect 0 36486 2839 36488
rect 0 36456 800 36486
rect 2773 36483 2839 36486
rect 5165 36546 5231 36549
rect 26190 36546 26250 36622
rect 36169 36619 36235 36622
rect 5165 36544 26250 36546
rect 5165 36488 5170 36544
rect 5226 36488 26250 36544
rect 5165 36486 26250 36488
rect 5165 36483 5231 36486
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 36629 36410 36695 36413
rect 39200 36410 40000 36440
rect 36629 36408 40000 36410
rect 36629 36352 36634 36408
rect 36690 36352 40000 36408
rect 36629 36350 40000 36352
rect 36629 36347 36695 36350
rect 39200 36320 40000 36350
rect 2037 36274 2103 36277
rect 30741 36274 30807 36277
rect 2037 36272 30807 36274
rect 2037 36216 2042 36272
rect 2098 36216 30746 36272
rect 30802 36216 30807 36272
rect 2037 36214 30807 36216
rect 2037 36211 2103 36214
rect 30741 36211 30807 36214
rect 0 36138 800 36168
rect 1853 36138 1919 36141
rect 0 36136 1919 36138
rect 0 36080 1858 36136
rect 1914 36080 1919 36136
rect 0 36078 1919 36080
rect 0 36048 800 36078
rect 1853 36075 1919 36078
rect 30281 36138 30347 36141
rect 34513 36138 34579 36141
rect 30281 36136 34579 36138
rect 30281 36080 30286 36136
rect 30342 36080 34518 36136
rect 34574 36080 34579 36136
rect 30281 36078 34579 36080
rect 30281 36075 30347 36078
rect 34513 36075 34579 36078
rect 35525 36002 35591 36005
rect 39200 36002 40000 36032
rect 35525 36000 40000 36002
rect 35525 35944 35530 36000
rect 35586 35944 40000 36000
rect 35525 35942 40000 35944
rect 35525 35939 35591 35942
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 39200 35912 40000 35942
rect 19568 35871 19888 35872
rect 0 35730 800 35760
rect 2589 35730 2655 35733
rect 0 35728 2655 35730
rect 0 35672 2594 35728
rect 2650 35672 2655 35728
rect 0 35670 2655 35672
rect 0 35640 800 35670
rect 2589 35667 2655 35670
rect 38009 35458 38075 35461
rect 39200 35458 40000 35488
rect 38009 35456 40000 35458
rect 38009 35400 38014 35456
rect 38070 35400 40000 35456
rect 38009 35398 40000 35400
rect 38009 35395 38075 35398
rect 4208 35392 4528 35393
rect 0 35322 800 35352
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 39200 35368 40000 35398
rect 34928 35327 35248 35328
rect 3049 35322 3115 35325
rect 0 35320 3115 35322
rect 0 35264 3054 35320
rect 3110 35264 3115 35320
rect 0 35262 3115 35264
rect 0 35232 800 35262
rect 3049 35259 3115 35262
rect 36721 35050 36787 35053
rect 39200 35050 40000 35080
rect 36721 35048 40000 35050
rect 36721 34992 36726 35048
rect 36782 34992 40000 35048
rect 36721 34990 40000 34992
rect 36721 34987 36787 34990
rect 39200 34960 40000 34990
rect 0 34914 800 34944
rect 2221 34914 2287 34917
rect 0 34912 2287 34914
rect 0 34856 2226 34912
rect 2282 34856 2287 34912
rect 0 34854 2287 34856
rect 0 34824 800 34854
rect 2221 34851 2287 34854
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 38009 34642 38075 34645
rect 39200 34642 40000 34672
rect 38009 34640 40000 34642
rect 38009 34584 38014 34640
rect 38070 34584 40000 34640
rect 38009 34582 40000 34584
rect 38009 34579 38075 34582
rect 39200 34552 40000 34582
rect 0 34506 800 34536
rect 1853 34506 1919 34509
rect 0 34504 1919 34506
rect 0 34448 1858 34504
rect 1914 34448 1919 34504
rect 0 34446 1919 34448
rect 0 34416 800 34446
rect 1853 34443 1919 34446
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 37181 34234 37247 34237
rect 39200 34234 40000 34264
rect 37181 34232 40000 34234
rect 37181 34176 37186 34232
rect 37242 34176 40000 34232
rect 37181 34174 40000 34176
rect 37181 34171 37247 34174
rect 39200 34144 40000 34174
rect 0 34098 800 34128
rect 1485 34098 1551 34101
rect 0 34096 1551 34098
rect 0 34040 1490 34096
rect 1546 34040 1551 34096
rect 0 34038 1551 34040
rect 0 34008 800 34038
rect 1485 34035 1551 34038
rect 38009 33826 38075 33829
rect 39200 33826 40000 33856
rect 38009 33824 40000 33826
rect 38009 33768 38014 33824
rect 38070 33768 40000 33824
rect 38009 33766 40000 33768
rect 38009 33763 38075 33766
rect 19568 33760 19888 33761
rect 0 33690 800 33720
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 39200 33736 40000 33766
rect 19568 33695 19888 33696
rect 1853 33690 1919 33693
rect 0 33688 1919 33690
rect 0 33632 1858 33688
rect 1914 33632 1919 33688
rect 0 33630 1919 33632
rect 0 33600 800 33630
rect 1853 33627 1919 33630
rect 37365 33418 37431 33421
rect 39200 33418 40000 33448
rect 37365 33416 40000 33418
rect 37365 33360 37370 33416
rect 37426 33360 40000 33416
rect 37365 33358 40000 33360
rect 37365 33355 37431 33358
rect 39200 33328 40000 33358
rect 0 33282 800 33312
rect 1485 33282 1551 33285
rect 0 33280 1551 33282
rect 0 33224 1490 33280
rect 1546 33224 1551 33280
rect 0 33222 1551 33224
rect 0 33192 800 33222
rect 1485 33219 1551 33222
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 38009 33010 38075 33013
rect 39200 33010 40000 33040
rect 38009 33008 40000 33010
rect 38009 32952 38014 33008
rect 38070 32952 40000 33008
rect 38009 32950 40000 32952
rect 38009 32947 38075 32950
rect 39200 32920 40000 32950
rect 0 32874 800 32904
rect 1853 32874 1919 32877
rect 0 32872 1919 32874
rect 0 32816 1858 32872
rect 1914 32816 1919 32872
rect 0 32814 1919 32816
rect 0 32784 800 32814
rect 1853 32811 1919 32814
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 37457 32602 37523 32605
rect 39200 32602 40000 32632
rect 37457 32600 40000 32602
rect 37457 32544 37462 32600
rect 37518 32544 40000 32600
rect 37457 32542 40000 32544
rect 37457 32539 37523 32542
rect 39200 32512 40000 32542
rect 0 32466 800 32496
rect 2773 32466 2839 32469
rect 0 32464 2839 32466
rect 0 32408 2778 32464
rect 2834 32408 2839 32464
rect 0 32406 2839 32408
rect 0 32376 800 32406
rect 2773 32403 2839 32406
rect 38009 32194 38075 32197
rect 39200 32194 40000 32224
rect 38009 32192 40000 32194
rect 38009 32136 38014 32192
rect 38070 32136 40000 32192
rect 38009 32134 40000 32136
rect 38009 32131 38075 32134
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 39200 32104 40000 32134
rect 34928 32063 35248 32064
rect 1485 32058 1551 32061
rect 0 32056 1551 32058
rect 0 32000 1490 32056
rect 1546 32000 1551 32056
rect 0 31998 1551 32000
rect 0 31968 800 31998
rect 1485 31995 1551 31998
rect 37273 31786 37339 31789
rect 39200 31786 40000 31816
rect 37273 31784 40000 31786
rect 37273 31728 37278 31784
rect 37334 31728 40000 31784
rect 37273 31726 40000 31728
rect 37273 31723 37339 31726
rect 39200 31696 40000 31726
rect 0 31650 800 31680
rect 1853 31650 1919 31653
rect 0 31648 1919 31650
rect 0 31592 1858 31648
rect 1914 31592 1919 31648
rect 0 31590 1919 31592
rect 0 31560 800 31590
rect 1853 31587 1919 31590
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 38101 31378 38167 31381
rect 39200 31378 40000 31408
rect 38101 31376 40000 31378
rect 38101 31320 38106 31376
rect 38162 31320 40000 31376
rect 38101 31318 40000 31320
rect 38101 31315 38167 31318
rect 39200 31288 40000 31318
rect 0 31242 800 31272
rect 2129 31242 2195 31245
rect 0 31240 2195 31242
rect 0 31184 2134 31240
rect 2190 31184 2195 31240
rect 0 31182 2195 31184
rect 0 31152 800 31182
rect 2129 31179 2195 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30834 800 30864
rect 1485 30834 1551 30837
rect 0 30832 1551 30834
rect 0 30776 1490 30832
rect 1546 30776 1551 30832
rect 0 30774 1551 30776
rect 0 30744 800 30774
rect 1485 30771 1551 30774
rect 38009 30834 38075 30837
rect 39200 30834 40000 30864
rect 38009 30832 40000 30834
rect 38009 30776 38014 30832
rect 38070 30776 40000 30832
rect 38009 30774 40000 30776
rect 38009 30771 38075 30774
rect 39200 30744 40000 30774
rect 19568 30496 19888 30497
rect 0 30426 800 30456
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 1853 30426 1919 30429
rect 0 30424 1919 30426
rect 0 30368 1858 30424
rect 1914 30368 1919 30424
rect 0 30366 1919 30368
rect 0 30336 800 30366
rect 1853 30363 1919 30366
rect 38009 30426 38075 30429
rect 39200 30426 40000 30456
rect 38009 30424 40000 30426
rect 38009 30368 38014 30424
rect 38070 30368 40000 30424
rect 38009 30366 40000 30368
rect 38009 30363 38075 30366
rect 39200 30336 40000 30366
rect 0 30018 800 30048
rect 2221 30018 2287 30021
rect 0 30016 2287 30018
rect 0 29960 2226 30016
rect 2282 29960 2287 30016
rect 0 29958 2287 29960
rect 0 29928 800 29958
rect 2221 29955 2287 29958
rect 37365 30018 37431 30021
rect 39200 30018 40000 30048
rect 37365 30016 40000 30018
rect 37365 29960 37370 30016
rect 37426 29960 40000 30016
rect 37365 29958 40000 29960
rect 37365 29955 37431 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 39200 29928 40000 29958
rect 34928 29887 35248 29888
rect 0 29610 800 29640
rect 2773 29610 2839 29613
rect 0 29608 2839 29610
rect 0 29552 2778 29608
rect 2834 29552 2839 29608
rect 0 29550 2839 29552
rect 0 29520 800 29550
rect 2773 29547 2839 29550
rect 38009 29610 38075 29613
rect 39200 29610 40000 29640
rect 38009 29608 40000 29610
rect 38009 29552 38014 29608
rect 38070 29552 40000 29608
rect 38009 29550 40000 29552
rect 38009 29547 38075 29550
rect 39200 29520 40000 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 0 29202 800 29232
rect 1853 29202 1919 29205
rect 0 29200 1919 29202
rect 0 29144 1858 29200
rect 1914 29144 1919 29200
rect 0 29142 1919 29144
rect 0 29112 800 29142
rect 1853 29139 1919 29142
rect 38101 29202 38167 29205
rect 39200 29202 40000 29232
rect 38101 29200 40000 29202
rect 38101 29144 38106 29200
rect 38162 29144 40000 29200
rect 38101 29142 40000 29144
rect 38101 29139 38167 29142
rect 39200 29112 40000 29142
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 2221 28794 2287 28797
rect 0 28792 2287 28794
rect 0 28736 2226 28792
rect 2282 28736 2287 28792
rect 0 28734 2287 28736
rect 0 28704 800 28734
rect 2221 28731 2287 28734
rect 37181 28794 37247 28797
rect 39200 28794 40000 28824
rect 37181 28792 40000 28794
rect 37181 28736 37186 28792
rect 37242 28736 40000 28792
rect 37181 28734 40000 28736
rect 37181 28731 37247 28734
rect 39200 28704 40000 28734
rect 0 28386 800 28416
rect 1485 28386 1551 28389
rect 0 28384 1551 28386
rect 0 28328 1490 28384
rect 1546 28328 1551 28384
rect 0 28326 1551 28328
rect 0 28296 800 28326
rect 1485 28323 1551 28326
rect 38009 28386 38075 28389
rect 39200 28386 40000 28416
rect 38009 28384 40000 28386
rect 38009 28328 38014 28384
rect 38070 28328 40000 28384
rect 38009 28326 40000 28328
rect 38009 28323 38075 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 39200 28296 40000 28326
rect 19568 28255 19888 28256
rect 0 27978 800 28008
rect 1853 27978 1919 27981
rect 0 27976 1919 27978
rect 0 27920 1858 27976
rect 1914 27920 1919 27976
rect 0 27918 1919 27920
rect 0 27888 800 27918
rect 1853 27915 1919 27918
rect 37273 27978 37339 27981
rect 39200 27978 40000 28008
rect 37273 27976 40000 27978
rect 37273 27920 37278 27976
rect 37334 27920 40000 27976
rect 37273 27918 40000 27920
rect 37273 27915 37339 27918
rect 39200 27888 40000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27570 800 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 800 27510
rect 2773 27507 2839 27510
rect 37181 27570 37247 27573
rect 39200 27570 40000 27600
rect 37181 27568 40000 27570
rect 37181 27512 37186 27568
rect 37242 27512 40000 27568
rect 37181 27510 40000 27512
rect 37181 27507 37247 27510
rect 39200 27480 40000 27510
rect 19568 27232 19888 27233
rect 0 27162 800 27192
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 1485 27162 1551 27165
rect 0 27160 1551 27162
rect 0 27104 1490 27160
rect 1546 27104 1551 27160
rect 0 27102 1551 27104
rect 0 27072 800 27102
rect 1485 27099 1551 27102
rect 38009 27162 38075 27165
rect 39200 27162 40000 27192
rect 38009 27160 40000 27162
rect 38009 27104 38014 27160
rect 38070 27104 40000 27160
rect 38009 27102 40000 27104
rect 38009 27099 38075 27102
rect 39200 27072 40000 27102
rect 0 26890 800 26920
rect 1853 26890 1919 26893
rect 0 26888 1919 26890
rect 0 26832 1858 26888
rect 1914 26832 1919 26888
rect 0 26830 1919 26832
rect 0 26800 800 26830
rect 1853 26827 1919 26830
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 38009 26618 38075 26621
rect 39200 26618 40000 26648
rect 38009 26616 40000 26618
rect 38009 26560 38014 26616
rect 38070 26560 40000 26616
rect 38009 26558 40000 26560
rect 38009 26555 38075 26558
rect 39200 26528 40000 26558
rect 0 26482 800 26512
rect 2221 26482 2287 26485
rect 0 26480 2287 26482
rect 0 26424 2226 26480
rect 2282 26424 2287 26480
rect 0 26422 2287 26424
rect 0 26392 800 26422
rect 2221 26419 2287 26422
rect 38101 26210 38167 26213
rect 39200 26210 40000 26240
rect 38101 26208 40000 26210
rect 38101 26152 38106 26208
rect 38162 26152 40000 26208
rect 38101 26150 40000 26152
rect 38101 26147 38167 26150
rect 19568 26144 19888 26145
rect 0 26074 800 26104
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 39200 26120 40000 26150
rect 19568 26079 19888 26080
rect 2773 26074 2839 26077
rect 0 26072 2839 26074
rect 0 26016 2778 26072
rect 2834 26016 2839 26072
rect 0 26014 2839 26016
rect 0 25984 800 26014
rect 2773 26011 2839 26014
rect 38009 25802 38075 25805
rect 39200 25802 40000 25832
rect 38009 25800 40000 25802
rect 38009 25744 38014 25800
rect 38070 25744 40000 25800
rect 38009 25742 40000 25744
rect 38009 25739 38075 25742
rect 39200 25712 40000 25742
rect 0 25666 800 25696
rect 1945 25666 2011 25669
rect 0 25664 2011 25666
rect 0 25608 1950 25664
rect 2006 25608 2011 25664
rect 0 25606 2011 25608
rect 0 25576 800 25606
rect 1945 25603 2011 25606
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 38009 25394 38075 25397
rect 39200 25394 40000 25424
rect 38009 25392 40000 25394
rect 38009 25336 38014 25392
rect 38070 25336 40000 25392
rect 38009 25334 40000 25336
rect 38009 25331 38075 25334
rect 39200 25304 40000 25334
rect 0 25258 800 25288
rect 2129 25258 2195 25261
rect 0 25256 2195 25258
rect 0 25200 2134 25256
rect 2190 25200 2195 25256
rect 0 25198 2195 25200
rect 0 25168 800 25198
rect 2129 25195 2195 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 37365 24986 37431 24989
rect 39200 24986 40000 25016
rect 37365 24984 40000 24986
rect 37365 24928 37370 24984
rect 37426 24928 40000 24984
rect 37365 24926 40000 24928
rect 37365 24923 37431 24926
rect 39200 24896 40000 24926
rect 0 24850 800 24880
rect 1485 24850 1551 24853
rect 0 24848 1551 24850
rect 0 24792 1490 24848
rect 1546 24792 1551 24848
rect 0 24790 1551 24792
rect 0 24760 800 24790
rect 1485 24787 1551 24790
rect 38009 24578 38075 24581
rect 39200 24578 40000 24608
rect 38009 24576 40000 24578
rect 38009 24520 38014 24576
rect 38070 24520 40000 24576
rect 38009 24518 40000 24520
rect 38009 24515 38075 24518
rect 4208 24512 4528 24513
rect 0 24442 800 24472
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 39200 24488 40000 24518
rect 34928 24447 35248 24448
rect 1853 24442 1919 24445
rect 0 24440 1919 24442
rect 0 24384 1858 24440
rect 1914 24384 1919 24440
rect 0 24382 1919 24384
rect 0 24352 800 24382
rect 1853 24379 1919 24382
rect 38009 24170 38075 24173
rect 39200 24170 40000 24200
rect 38009 24168 40000 24170
rect 38009 24112 38014 24168
rect 38070 24112 40000 24168
rect 38009 24110 40000 24112
rect 38009 24107 38075 24110
rect 39200 24080 40000 24110
rect 0 24034 800 24064
rect 1393 24034 1459 24037
rect 0 24032 1459 24034
rect 0 23976 1398 24032
rect 1454 23976 1459 24032
rect 0 23974 1459 23976
rect 0 23944 800 23974
rect 1393 23971 1459 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 37365 23762 37431 23765
rect 39200 23762 40000 23792
rect 37365 23760 40000 23762
rect 37365 23704 37370 23760
rect 37426 23704 40000 23760
rect 37365 23702 40000 23704
rect 37365 23699 37431 23702
rect 39200 23672 40000 23702
rect 0 23626 800 23656
rect 1485 23626 1551 23629
rect 0 23624 1551 23626
rect 0 23568 1490 23624
rect 1546 23568 1551 23624
rect 0 23566 1551 23568
rect 0 23536 800 23566
rect 1485 23563 1551 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 38009 23354 38075 23357
rect 39200 23354 40000 23384
rect 38009 23352 40000 23354
rect 38009 23296 38014 23352
rect 38070 23296 40000 23352
rect 38009 23294 40000 23296
rect 38009 23291 38075 23294
rect 39200 23264 40000 23294
rect 0 23218 800 23248
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23128 800 23158
rect 1853 23155 1919 23158
rect 38009 22946 38075 22949
rect 39200 22946 40000 22976
rect 38009 22944 40000 22946
rect 38009 22888 38014 22944
rect 38070 22888 40000 22944
rect 38009 22886 40000 22888
rect 38009 22883 38075 22886
rect 19568 22880 19888 22881
rect 0 22810 800 22840
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 39200 22856 40000 22886
rect 19568 22815 19888 22816
rect 2129 22810 2195 22813
rect 0 22808 2195 22810
rect 0 22752 2134 22808
rect 2190 22752 2195 22808
rect 0 22750 2195 22752
rect 0 22720 800 22750
rect 2129 22747 2195 22750
rect 37365 22538 37431 22541
rect 39200 22538 40000 22568
rect 37365 22536 40000 22538
rect 37365 22480 37370 22536
rect 37426 22480 40000 22536
rect 37365 22478 40000 22480
rect 37365 22475 37431 22478
rect 39200 22448 40000 22478
rect 0 22402 800 22432
rect 1485 22402 1551 22405
rect 0 22400 1551 22402
rect 0 22344 1490 22400
rect 1546 22344 1551 22400
rect 0 22342 1551 22344
rect 0 22312 800 22342
rect 1485 22339 1551 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21994 800 22024
rect 1853 21994 1919 21997
rect 0 21992 1919 21994
rect 0 21936 1858 21992
rect 1914 21936 1919 21992
rect 0 21934 1919 21936
rect 0 21904 800 21934
rect 1853 21931 1919 21934
rect 38009 21994 38075 21997
rect 39200 21994 40000 22024
rect 38009 21992 40000 21994
rect 38009 21936 38014 21992
rect 38070 21936 40000 21992
rect 38009 21934 40000 21936
rect 38009 21931 38075 21934
rect 39200 21904 40000 21934
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 0 21586 800 21616
rect 2773 21586 2839 21589
rect 0 21584 2839 21586
rect 0 21528 2778 21584
rect 2834 21528 2839 21584
rect 0 21526 2839 21528
rect 0 21496 800 21526
rect 2773 21523 2839 21526
rect 38101 21586 38167 21589
rect 39200 21586 40000 21616
rect 38101 21584 40000 21586
rect 38101 21528 38106 21584
rect 38162 21528 40000 21584
rect 38101 21526 40000 21528
rect 38101 21523 38167 21526
rect 39200 21496 40000 21526
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 1485 21178 1551 21181
rect 0 21176 1551 21178
rect 0 21120 1490 21176
rect 1546 21120 1551 21176
rect 0 21118 1551 21120
rect 0 21088 800 21118
rect 1485 21115 1551 21118
rect 37365 21178 37431 21181
rect 39200 21178 40000 21208
rect 37365 21176 40000 21178
rect 37365 21120 37370 21176
rect 37426 21120 40000 21176
rect 37365 21118 40000 21120
rect 37365 21115 37431 21118
rect 39200 21088 40000 21118
rect 0 20770 800 20800
rect 1853 20770 1919 20773
rect 0 20768 1919 20770
rect 0 20712 1858 20768
rect 1914 20712 1919 20768
rect 0 20710 1919 20712
rect 0 20680 800 20710
rect 1853 20707 1919 20710
rect 38009 20770 38075 20773
rect 39200 20770 40000 20800
rect 38009 20768 40000 20770
rect 38009 20712 38014 20768
rect 38070 20712 40000 20768
rect 38009 20710 40000 20712
rect 38009 20707 38075 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 39200 20680 40000 20710
rect 19568 20639 19888 20640
rect 0 20362 800 20392
rect 2129 20362 2195 20365
rect 0 20360 2195 20362
rect 0 20304 2134 20360
rect 2190 20304 2195 20360
rect 0 20302 2195 20304
rect 0 20272 800 20302
rect 2129 20299 2195 20302
rect 38101 20362 38167 20365
rect 39200 20362 40000 20392
rect 38101 20360 40000 20362
rect 38101 20304 38106 20360
rect 38162 20304 40000 20360
rect 38101 20302 40000 20304
rect 38101 20299 38167 20302
rect 39200 20272 40000 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19954 800 19984
rect 1485 19954 1551 19957
rect 0 19952 1551 19954
rect 0 19896 1490 19952
rect 1546 19896 1551 19952
rect 0 19894 1551 19896
rect 0 19864 800 19894
rect 1485 19891 1551 19894
rect 37089 19954 37155 19957
rect 39200 19954 40000 19984
rect 37089 19952 40000 19954
rect 37089 19896 37094 19952
rect 37150 19896 40000 19952
rect 37089 19894 40000 19896
rect 37089 19891 37155 19894
rect 39200 19864 40000 19894
rect 19568 19616 19888 19617
rect 0 19546 800 19576
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 1853 19546 1919 19549
rect 0 19544 1919 19546
rect 0 19488 1858 19544
rect 1914 19488 1919 19544
rect 0 19486 1919 19488
rect 0 19456 800 19486
rect 1853 19483 1919 19486
rect 38009 19546 38075 19549
rect 39200 19546 40000 19576
rect 38009 19544 40000 19546
rect 38009 19488 38014 19544
rect 38070 19488 40000 19544
rect 38009 19486 40000 19488
rect 38009 19483 38075 19486
rect 39200 19456 40000 19486
rect 0 19138 800 19168
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 19048 800 19078
rect 2221 19075 2287 19078
rect 37181 19138 37247 19141
rect 39200 19138 40000 19168
rect 37181 19136 40000 19138
rect 37181 19080 37186 19136
rect 37242 19080 40000 19136
rect 37181 19078 40000 19080
rect 37181 19075 37247 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 39200 19048 40000 19078
rect 34928 19007 35248 19008
rect 0 18730 800 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 800 18670
rect 1485 18667 1551 18670
rect 37181 18730 37247 18733
rect 39200 18730 40000 18760
rect 37181 18728 40000 18730
rect 37181 18672 37186 18728
rect 37242 18672 40000 18728
rect 37181 18670 40000 18672
rect 37181 18667 37247 18670
rect 39200 18640 40000 18670
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 0 18322 800 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 800 18262
rect 1853 18259 1919 18262
rect 38009 18322 38075 18325
rect 39200 18322 40000 18352
rect 38009 18320 40000 18322
rect 38009 18264 38014 18320
rect 38070 18264 40000 18320
rect 38009 18262 40000 18264
rect 38009 18259 38075 18262
rect 39200 18232 40000 18262
rect 4208 17984 4528 17985
rect 0 17914 800 17944
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 2129 17914 2195 17917
rect 0 17912 2195 17914
rect 0 17856 2134 17912
rect 2190 17856 2195 17912
rect 0 17854 2195 17856
rect 0 17824 800 17854
rect 2129 17851 2195 17854
rect 38009 17778 38075 17781
rect 39200 17778 40000 17808
rect 38009 17776 40000 17778
rect 38009 17720 38014 17776
rect 38070 17720 40000 17776
rect 38009 17718 40000 17720
rect 38009 17715 38075 17718
rect 39200 17688 40000 17718
rect 0 17506 800 17536
rect 1485 17506 1551 17509
rect 0 17504 1551 17506
rect 0 17448 1490 17504
rect 1546 17448 1551 17504
rect 0 17446 1551 17448
rect 0 17416 800 17446
rect 1485 17443 1551 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 38101 17370 38167 17373
rect 39200 17370 40000 17400
rect 38101 17368 40000 17370
rect 38101 17312 38106 17368
rect 38162 17312 40000 17368
rect 38101 17310 40000 17312
rect 38101 17307 38167 17310
rect 39200 17280 40000 17310
rect 0 17098 800 17128
rect 2865 17098 2931 17101
rect 0 17096 2931 17098
rect 0 17040 2870 17096
rect 2926 17040 2931 17096
rect 0 17038 2931 17040
rect 0 17008 800 17038
rect 2865 17035 2931 17038
rect 38009 16962 38075 16965
rect 39200 16962 40000 16992
rect 38009 16960 40000 16962
rect 38009 16904 38014 16960
rect 38070 16904 40000 16960
rect 38009 16902 40000 16904
rect 38009 16899 38075 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 39200 16872 40000 16902
rect 34928 16831 35248 16832
rect 0 16690 800 16720
rect 2221 16690 2287 16693
rect 0 16688 2287 16690
rect 0 16632 2226 16688
rect 2282 16632 2287 16688
rect 0 16630 2287 16632
rect 0 16600 800 16630
rect 2221 16627 2287 16630
rect 38009 16554 38075 16557
rect 39200 16554 40000 16584
rect 38009 16552 40000 16554
rect 38009 16496 38014 16552
rect 38070 16496 40000 16552
rect 38009 16494 40000 16496
rect 38009 16491 38075 16494
rect 39200 16464 40000 16494
rect 19568 16352 19888 16353
rect 0 16282 800 16312
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 2773 16282 2839 16285
rect 0 16280 2839 16282
rect 0 16224 2778 16280
rect 2834 16224 2839 16280
rect 0 16222 2839 16224
rect 0 16192 800 16222
rect 2773 16219 2839 16222
rect 37365 16146 37431 16149
rect 39200 16146 40000 16176
rect 37365 16144 40000 16146
rect 37365 16088 37370 16144
rect 37426 16088 40000 16144
rect 37365 16086 40000 16088
rect 37365 16083 37431 16086
rect 39200 16056 40000 16086
rect 0 15874 800 15904
rect 1853 15874 1919 15877
rect 0 15872 1919 15874
rect 0 15816 1858 15872
rect 1914 15816 1919 15872
rect 0 15814 1919 15816
rect 0 15784 800 15814
rect 1853 15811 1919 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 38009 15738 38075 15741
rect 39200 15738 40000 15768
rect 38009 15736 40000 15738
rect 38009 15680 38014 15736
rect 38070 15680 40000 15736
rect 38009 15678 40000 15680
rect 38009 15675 38075 15678
rect 39200 15648 40000 15678
rect 0 15466 800 15496
rect 2221 15466 2287 15469
rect 0 15464 2287 15466
rect 0 15408 2226 15464
rect 2282 15408 2287 15464
rect 0 15406 2287 15408
rect 0 15376 800 15406
rect 2221 15403 2287 15406
rect 37273 15330 37339 15333
rect 39200 15330 40000 15360
rect 37273 15328 40000 15330
rect 37273 15272 37278 15328
rect 37334 15272 40000 15328
rect 37273 15270 40000 15272
rect 37273 15267 37339 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 39200 15240 40000 15270
rect 19568 15199 19888 15200
rect 0 15058 800 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 800 14998
rect 2773 14995 2839 14998
rect 36261 14922 36327 14925
rect 39200 14922 40000 14952
rect 36261 14920 40000 14922
rect 36261 14864 36266 14920
rect 36322 14864 40000 14920
rect 36261 14862 40000 14864
rect 36261 14859 36327 14862
rect 39200 14832 40000 14862
rect 4208 14720 4528 14721
rect 0 14650 800 14680
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 38009 14514 38075 14517
rect 39200 14514 40000 14544
rect 38009 14512 40000 14514
rect 38009 14456 38014 14512
rect 38070 14456 40000 14512
rect 38009 14454 40000 14456
rect 38009 14451 38075 14454
rect 39200 14424 40000 14454
rect 0 14242 800 14272
rect 1393 14242 1459 14245
rect 0 14240 1459 14242
rect 0 14184 1398 14240
rect 1454 14184 1459 14240
rect 0 14182 1459 14184
rect 0 14152 800 14182
rect 1393 14179 1459 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 38009 14106 38075 14109
rect 39200 14106 40000 14136
rect 38009 14104 40000 14106
rect 38009 14048 38014 14104
rect 38070 14048 40000 14104
rect 38009 14046 40000 14048
rect 38009 14043 38075 14046
rect 39200 14016 40000 14046
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 37181 13698 37247 13701
rect 39200 13698 40000 13728
rect 37181 13696 40000 13698
rect 37181 13640 37186 13696
rect 37242 13640 40000 13696
rect 37181 13638 40000 13640
rect 37181 13635 37247 13638
rect 4208 13632 4528 13633
rect 0 13562 800 13592
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 39200 13608 40000 13638
rect 34928 13567 35248 13568
rect 1853 13562 1919 13565
rect 0 13560 1919 13562
rect 0 13504 1858 13560
rect 1914 13504 1919 13560
rect 0 13502 1919 13504
rect 0 13472 800 13502
rect 1853 13499 1919 13502
rect 0 13154 800 13184
rect 2129 13154 2195 13157
rect 0 13152 2195 13154
rect 0 13096 2134 13152
rect 2190 13096 2195 13152
rect 0 13094 2195 13096
rect 0 13064 800 13094
rect 2129 13091 2195 13094
rect 38009 13154 38075 13157
rect 39200 13154 40000 13184
rect 38009 13152 40000 13154
rect 38009 13096 38014 13152
rect 38070 13096 40000 13152
rect 38009 13094 40000 13096
rect 38009 13091 38075 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 39200 13064 40000 13094
rect 19568 13023 19888 13024
rect 0 12746 800 12776
rect 1485 12746 1551 12749
rect 0 12744 1551 12746
rect 0 12688 1490 12744
rect 1546 12688 1551 12744
rect 0 12686 1551 12688
rect 0 12656 800 12686
rect 1485 12683 1551 12686
rect 38009 12746 38075 12749
rect 39200 12746 40000 12776
rect 38009 12744 40000 12746
rect 38009 12688 38014 12744
rect 38070 12688 40000 12744
rect 38009 12686 40000 12688
rect 38009 12683 38075 12686
rect 39200 12656 40000 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 1853 12472 1919 12477
rect 1853 12416 1858 12472
rect 1914 12416 1919 12472
rect 1853 12411 1919 12416
rect 0 12338 800 12368
rect 1856 12338 1916 12411
rect 0 12278 1916 12338
rect 38101 12338 38167 12341
rect 39200 12338 40000 12368
rect 38101 12336 40000 12338
rect 38101 12280 38106 12336
rect 38162 12280 40000 12336
rect 38101 12278 40000 12280
rect 0 12248 800 12278
rect 38101 12275 38167 12278
rect 39200 12248 40000 12278
rect 2037 12202 2103 12205
rect 27797 12202 27863 12205
rect 2037 12200 27863 12202
rect 2037 12144 2042 12200
rect 2098 12144 27802 12200
rect 27858 12144 27863 12200
rect 2037 12142 27863 12144
rect 2037 12139 2103 12142
rect 27797 12139 27863 12142
rect 19568 12000 19888 12001
rect 0 11930 800 11960
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 2129 11930 2195 11933
rect 0 11928 2195 11930
rect 0 11872 2134 11928
rect 2190 11872 2195 11928
rect 0 11870 2195 11872
rect 0 11840 800 11870
rect 2129 11867 2195 11870
rect 38009 11930 38075 11933
rect 39200 11930 40000 11960
rect 38009 11928 40000 11930
rect 38009 11872 38014 11928
rect 38070 11872 40000 11928
rect 38009 11870 40000 11872
rect 38009 11867 38075 11870
rect 39200 11840 40000 11870
rect 0 11522 800 11552
rect 1485 11522 1551 11525
rect 0 11520 1551 11522
rect 0 11464 1490 11520
rect 1546 11464 1551 11520
rect 0 11462 1551 11464
rect 0 11432 800 11462
rect 1485 11459 1551 11462
rect 38009 11522 38075 11525
rect 39200 11522 40000 11552
rect 38009 11520 40000 11522
rect 38009 11464 38014 11520
rect 38070 11464 40000 11520
rect 38009 11462 40000 11464
rect 38009 11459 38075 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 39200 11432 40000 11462
rect 34928 11391 35248 11392
rect 0 11114 800 11144
rect 1853 11114 1919 11117
rect 0 11112 1919 11114
rect 0 11056 1858 11112
rect 1914 11056 1919 11112
rect 0 11054 1919 11056
rect 0 11024 800 11054
rect 1853 11051 1919 11054
rect 2037 11114 2103 11117
rect 27705 11114 27771 11117
rect 2037 11112 27771 11114
rect 2037 11056 2042 11112
rect 2098 11056 27710 11112
rect 27766 11056 27771 11112
rect 2037 11054 27771 11056
rect 2037 11051 2103 11054
rect 27705 11051 27771 11054
rect 37365 11114 37431 11117
rect 39200 11114 40000 11144
rect 37365 11112 40000 11114
rect 37365 11056 37370 11112
rect 37426 11056 40000 11112
rect 37365 11054 40000 11056
rect 37365 11051 37431 11054
rect 39200 11024 40000 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 0 10706 800 10736
rect 2773 10706 2839 10709
rect 0 10704 2839 10706
rect 0 10648 2778 10704
rect 2834 10648 2839 10704
rect 0 10646 2839 10648
rect 0 10616 800 10646
rect 2773 10643 2839 10646
rect 38009 10706 38075 10709
rect 39200 10706 40000 10736
rect 38009 10704 40000 10706
rect 38009 10648 38014 10704
rect 38070 10648 40000 10704
rect 38009 10646 40000 10648
rect 38009 10643 38075 10646
rect 39200 10616 40000 10646
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 38009 10298 38075 10301
rect 39200 10298 40000 10328
rect 38009 10296 40000 10298
rect 38009 10240 38014 10296
rect 38070 10240 40000 10296
rect 38009 10238 40000 10240
rect 38009 10235 38075 10238
rect 39200 10208 40000 10238
rect 0 9890 800 9920
rect 1853 9890 1919 9893
rect 0 9888 1919 9890
rect 0 9832 1858 9888
rect 1914 9832 1919 9888
rect 0 9830 1919 9832
rect 0 9800 800 9830
rect 1853 9827 1919 9830
rect 36537 9890 36603 9893
rect 39200 9890 40000 9920
rect 36537 9888 40000 9890
rect 36537 9832 36542 9888
rect 36598 9832 40000 9888
rect 36537 9830 40000 9832
rect 36537 9827 36603 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 39200 9800 40000 9830
rect 19568 9759 19888 9760
rect 0 9482 800 9512
rect 1393 9482 1459 9485
rect 0 9480 1459 9482
rect 0 9424 1398 9480
rect 1454 9424 1459 9480
rect 0 9422 1459 9424
rect 0 9392 800 9422
rect 1393 9419 1459 9422
rect 38009 9482 38075 9485
rect 39200 9482 40000 9512
rect 38009 9480 40000 9482
rect 38009 9424 38014 9480
rect 38070 9424 40000 9480
rect 38009 9422 40000 9424
rect 38009 9419 38075 9422
rect 39200 9392 40000 9422
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 9074 800 9104
rect 2037 9074 2103 9077
rect 0 9072 2103 9074
rect 0 9016 2042 9072
rect 2098 9016 2103 9072
rect 0 9014 2103 9016
rect 0 8984 800 9014
rect 2037 9011 2103 9014
rect 38101 8938 38167 8941
rect 39200 8938 40000 8968
rect 38101 8936 40000 8938
rect 38101 8880 38106 8936
rect 38162 8880 40000 8936
rect 38101 8878 40000 8880
rect 38101 8875 38167 8878
rect 39200 8848 40000 8878
rect 19568 8736 19888 8737
rect 0 8666 800 8696
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 800 8606
rect 1485 8603 1551 8606
rect 37365 8530 37431 8533
rect 39200 8530 40000 8560
rect 37365 8528 40000 8530
rect 37365 8472 37370 8528
rect 37426 8472 40000 8528
rect 37365 8470 40000 8472
rect 37365 8467 37431 8470
rect 39200 8440 40000 8470
rect 0 8258 800 8288
rect 1853 8258 1919 8261
rect 0 8256 1919 8258
rect 0 8200 1858 8256
rect 1914 8200 1919 8256
rect 0 8198 1919 8200
rect 0 8168 800 8198
rect 1853 8195 1919 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 38009 8122 38075 8125
rect 39200 8122 40000 8152
rect 38009 8120 40000 8122
rect 38009 8064 38014 8120
rect 38070 8064 40000 8120
rect 38009 8062 40000 8064
rect 38009 8059 38075 8062
rect 39200 8032 40000 8062
rect 0 7850 800 7880
rect 1393 7850 1459 7853
rect 0 7848 1459 7850
rect 0 7792 1398 7848
rect 1454 7792 1459 7848
rect 0 7790 1459 7792
rect 0 7760 800 7790
rect 1393 7787 1459 7790
rect 38009 7714 38075 7717
rect 39200 7714 40000 7744
rect 38009 7712 40000 7714
rect 38009 7656 38014 7712
rect 38070 7656 40000 7712
rect 38009 7654 40000 7656
rect 38009 7651 38075 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 39200 7624 40000 7654
rect 19568 7583 19888 7584
rect 0 7442 800 7472
rect 2037 7442 2103 7445
rect 0 7440 2103 7442
rect 0 7384 2042 7440
rect 2098 7384 2103 7440
rect 0 7382 2103 7384
rect 0 7352 800 7382
rect 2037 7379 2103 7382
rect 37365 7306 37431 7309
rect 39200 7306 40000 7336
rect 37365 7304 40000 7306
rect 37365 7248 37370 7304
rect 37426 7248 40000 7304
rect 37365 7246 40000 7248
rect 37365 7243 37431 7246
rect 39200 7216 40000 7246
rect 4208 7104 4528 7105
rect 0 7034 800 7064
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 1485 7034 1551 7037
rect 0 7032 1551 7034
rect 0 6976 1490 7032
rect 1546 6976 1551 7032
rect 0 6974 1551 6976
rect 0 6944 800 6974
rect 1485 6971 1551 6974
rect 38009 6898 38075 6901
rect 39200 6898 40000 6928
rect 38009 6896 40000 6898
rect 38009 6840 38014 6896
rect 38070 6840 40000 6896
rect 38009 6838 40000 6840
rect 38009 6835 38075 6838
rect 39200 6808 40000 6838
rect 0 6626 800 6656
rect 1853 6626 1919 6629
rect 0 6624 1919 6626
rect 0 6568 1858 6624
rect 1914 6568 1919 6624
rect 0 6566 1919 6568
rect 0 6536 800 6566
rect 1853 6563 1919 6566
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 38009 6490 38075 6493
rect 39200 6490 40000 6520
rect 38009 6488 40000 6490
rect 38009 6432 38014 6488
rect 38070 6432 40000 6488
rect 38009 6430 40000 6432
rect 38009 6427 38075 6430
rect 39200 6400 40000 6430
rect 0 6218 800 6248
rect 2129 6218 2195 6221
rect 0 6216 2195 6218
rect 0 6160 2134 6216
rect 2190 6160 2195 6216
rect 0 6158 2195 6160
rect 0 6128 800 6158
rect 2129 6155 2195 6158
rect 38009 6082 38075 6085
rect 39200 6082 40000 6112
rect 38009 6080 40000 6082
rect 38009 6024 38014 6080
rect 38070 6024 40000 6080
rect 38009 6022 40000 6024
rect 38009 6019 38075 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 39200 5992 40000 6022
rect 34928 5951 35248 5952
rect 0 5810 800 5840
rect 2221 5810 2287 5813
rect 0 5808 2287 5810
rect 0 5752 2226 5808
rect 2282 5752 2287 5808
rect 0 5750 2287 5752
rect 0 5720 800 5750
rect 2221 5747 2287 5750
rect 37365 5674 37431 5677
rect 39200 5674 40000 5704
rect 37365 5672 40000 5674
rect 37365 5616 37370 5672
rect 37426 5616 40000 5672
rect 37365 5614 40000 5616
rect 37365 5611 37431 5614
rect 39200 5584 40000 5614
rect 19568 5472 19888 5473
rect 0 5402 800 5432
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 1485 5402 1551 5405
rect 0 5400 1551 5402
rect 0 5344 1490 5400
rect 1546 5344 1551 5400
rect 0 5342 1551 5344
rect 0 5312 800 5342
rect 1485 5339 1551 5342
rect 38009 5266 38075 5269
rect 39200 5266 40000 5296
rect 38009 5264 40000 5266
rect 38009 5208 38014 5264
rect 38070 5208 40000 5264
rect 38009 5206 40000 5208
rect 38009 5203 38075 5206
rect 39200 5176 40000 5206
rect 0 4994 800 5024
rect 1853 4994 1919 4997
rect 0 4992 1919 4994
rect 0 4936 1858 4992
rect 1914 4936 1919 4992
rect 0 4934 1919 4936
rect 0 4904 800 4934
rect 1853 4931 1919 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 38009 4858 38075 4861
rect 39200 4858 40000 4888
rect 38009 4856 40000 4858
rect 38009 4800 38014 4856
rect 38070 4800 40000 4856
rect 38009 4798 40000 4800
rect 38009 4795 38075 4798
rect 39200 4768 40000 4798
rect 0 4586 800 4616
rect 2773 4586 2839 4589
rect 0 4584 2839 4586
rect 0 4528 2778 4584
rect 2834 4528 2839 4584
rect 0 4526 2839 4528
rect 0 4496 800 4526
rect 2773 4523 2839 4526
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 38009 4314 38075 4317
rect 39200 4314 40000 4344
rect 38009 4312 40000 4314
rect 38009 4256 38014 4312
rect 38070 4256 40000 4312
rect 38009 4254 40000 4256
rect 38009 4251 38075 4254
rect 39200 4224 40000 4254
rect 0 4178 800 4208
rect 1853 4178 1919 4181
rect 0 4176 1919 4178
rect 0 4120 1858 4176
rect 1914 4120 1919 4176
rect 0 4118 1919 4120
rect 0 4088 800 4118
rect 1853 4115 1919 4118
rect 3877 4042 3943 4045
rect 29913 4042 29979 4045
rect 3877 4040 29979 4042
rect 3877 3984 3882 4040
rect 3938 3984 29918 4040
rect 29974 3984 29979 4040
rect 3877 3982 29979 3984
rect 3877 3979 3943 3982
rect 29913 3979 29979 3982
rect 36077 3906 36143 3909
rect 39200 3906 40000 3936
rect 36077 3904 40000 3906
rect 36077 3848 36082 3904
rect 36138 3848 40000 3904
rect 36077 3846 40000 3848
rect 36077 3843 36143 3846
rect 4208 3840 4528 3841
rect 0 3770 800 3800
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 39200 3816 40000 3846
rect 34928 3775 35248 3776
rect 1485 3770 1551 3773
rect 0 3768 1551 3770
rect 0 3712 1490 3768
rect 1546 3712 1551 3768
rect 0 3710 1551 3712
rect 0 3680 800 3710
rect 1485 3707 1551 3710
rect 38009 3498 38075 3501
rect 39200 3498 40000 3528
rect 38009 3496 40000 3498
rect 38009 3440 38014 3496
rect 38070 3440 40000 3496
rect 38009 3438 40000 3440
rect 38009 3435 38075 3438
rect 39200 3408 40000 3438
rect 0 3362 800 3392
rect 1853 3362 1919 3365
rect 0 3360 1919 3362
rect 0 3304 1858 3360
rect 1914 3304 1919 3360
rect 0 3302 1919 3304
rect 0 3272 800 3302
rect 1853 3299 1919 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 38009 3090 38075 3093
rect 39200 3090 40000 3120
rect 38009 3088 40000 3090
rect 38009 3032 38014 3088
rect 38070 3032 40000 3088
rect 38009 3030 40000 3032
rect 38009 3027 38075 3030
rect 39200 3000 40000 3030
rect 0 2954 800 2984
rect 3233 2954 3299 2957
rect 0 2952 3299 2954
rect 0 2896 3238 2952
rect 3294 2896 3299 2952
rect 0 2894 3299 2896
rect 0 2864 800 2894
rect 3233 2891 3299 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 37273 2682 37339 2685
rect 39200 2682 40000 2712
rect 37273 2680 40000 2682
rect 37273 2624 37278 2680
rect 37334 2624 40000 2680
rect 37273 2622 40000 2624
rect 37273 2619 37339 2622
rect 39200 2592 40000 2622
rect 0 2546 800 2576
rect 1853 2546 1919 2549
rect 0 2544 1919 2546
rect 0 2488 1858 2544
rect 1914 2488 1919 2544
rect 0 2486 1919 2488
rect 0 2456 800 2486
rect 1853 2483 1919 2486
rect 35249 2274 35315 2277
rect 39200 2274 40000 2304
rect 35249 2272 40000 2274
rect 35249 2216 35254 2272
rect 35310 2216 40000 2272
rect 35249 2214 40000 2216
rect 35249 2211 35315 2214
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 39200 2184 40000 2214
rect 19568 2143 19888 2144
rect 4061 2138 4127 2141
rect 0 2136 4127 2138
rect 0 2080 4066 2136
rect 4122 2080 4127 2136
rect 0 2078 4127 2080
rect 0 2048 800 2078
rect 4061 2075 4127 2078
rect 38101 1866 38167 1869
rect 39200 1866 40000 1896
rect 38101 1864 40000 1866
rect 38101 1808 38106 1864
rect 38162 1808 40000 1864
rect 38101 1806 40000 1808
rect 38101 1803 38167 1806
rect 39200 1776 40000 1806
rect 0 1730 800 1760
rect 2773 1730 2839 1733
rect 0 1728 2839 1730
rect 0 1672 2778 1728
rect 2834 1672 2839 1728
rect 0 1670 2839 1672
rect 0 1640 800 1670
rect 2773 1667 2839 1670
rect 38009 1458 38075 1461
rect 39200 1458 40000 1488
rect 38009 1456 40000 1458
rect 38009 1400 38014 1456
rect 38070 1400 40000 1456
rect 38009 1398 40000 1400
rect 38009 1395 38075 1398
rect 39200 1368 40000 1398
rect 0 1322 800 1352
rect 3049 1322 3115 1325
rect 0 1320 3115 1322
rect 0 1264 3054 1320
rect 3110 1264 3115 1320
rect 0 1262 3115 1264
rect 0 1232 800 1262
rect 3049 1259 3115 1262
rect 35801 1050 35867 1053
rect 39200 1050 40000 1080
rect 35801 1048 40000 1050
rect 35801 992 35806 1048
rect 35862 992 40000 1048
rect 35801 990 40000 992
rect 35801 987 35867 990
rect 39200 960 40000 990
rect 0 914 800 944
rect 3969 914 4035 917
rect 0 912 4035 914
rect 0 856 3974 912
rect 4030 856 4035 912
rect 0 854 4035 856
rect 0 824 800 854
rect 3969 851 4035 854
rect 35709 642 35775 645
rect 39200 642 40000 672
rect 35709 640 40000 642
rect 35709 584 35714 640
rect 35770 584 40000 640
rect 35709 582 40000 584
rect 35709 579 35775 582
rect 39200 552 40000 582
rect 0 506 800 536
rect 3141 506 3207 509
rect 0 504 3207 506
rect 0 448 3146 504
rect 3202 448 3207 504
rect 0 446 3207 448
rect 0 416 800 446
rect 3141 443 3207 446
rect 0 234 800 264
rect 2865 234 2931 237
rect 0 232 2931 234
rect 0 176 2870 232
rect 2926 176 2931 232
rect 0 174 2931 176
rect 0 144 800 174
rect 2865 171 2931 174
rect 35617 234 35683 237
rect 39200 234 40000 264
rect 35617 232 40000 234
rect 35617 176 35622 232
rect 35678 176 40000 232
rect 35617 174 40000 176
rect 35617 171 35683 174
rect 39200 144 40000 174
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1644511149
transform -1 0 32936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1644511149
transform -1 0 33028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1644511149
transform 1 0 34040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1644511149
transform -1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1644511149
transform -1 0 33764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1644511149
transform -1 0 32752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1644511149
transform -1 0 32568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1644511149
transform 1 0 32568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1644511149
transform -1 0 32660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1644511149
transform 1 0 23736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1644511149
transform -1 0 22816 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1644511149
transform -1 0 22080 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__B
timestamp 1644511149
transform -1 0 21068 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__B
timestamp 1644511149
transform -1 0 21068 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__B
timestamp 1644511149
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__B
timestamp 1644511149
transform -1 0 21068 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B
timestamp 1644511149
transform -1 0 22264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1644511149
transform -1 0 30820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1644511149
transform -1 0 31648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__B
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1644511149
transform -1 0 29900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1644511149
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1644511149
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1644511149
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1644511149
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1644511149
transform 1 0 36156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1644511149
transform 1 0 35328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1644511149
transform -1 0 36432 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1644511149
transform -1 0 3496 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 1644511149
transform -1 0 36064 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1644511149
transform -1 0 3496 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1644511149
transform -1 0 4048 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1644511149
transform -1 0 5244 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1644511149
transform -1 0 5060 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__B
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__B
timestamp 1644511149
transform -1 0 23092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__B
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A_N
timestamp 1644511149
transform -1 0 25576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 1644511149
transform -1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1644511149
transform -1 0 27324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1644511149
transform 1 0 27232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1644511149
transform -1 0 27324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1644511149
transform -1 0 26496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1644511149
transform 1 0 26496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1644511149
transform -1 0 27876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1644511149
transform -1 0 27876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1644511149
transform 1 0 27784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1644511149
transform -1 0 28152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1644511149
transform 1 0 28336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1644511149
transform -1 0 28612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1644511149
transform -1 0 29808 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1644511149
transform -1 0 29716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1644511149
transform -1 0 29808 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1644511149
transform 1 0 28152 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1644511149
transform -1 0 29072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1644511149
transform -1 0 29072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1644511149
transform 1 0 27600 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1644511149
transform -1 0 26036 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1644511149
transform -1 0 26496 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1644511149
transform -1 0 26496 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1644511149
transform -1 0 25576 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1644511149
transform -1 0 25300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1644511149
transform -1 0 29900 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1644511149
transform -1 0 29440 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1644511149
transform -1 0 29440 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1644511149
transform -1 0 29532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1644511149
transform -1 0 29900 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A
timestamp 1644511149
transform 1 0 30544 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1644511149
transform 1 0 24472 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__B
timestamp 1644511149
transform 1 0 25484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1644511149
transform -1 0 24104 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__B
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1644511149
transform -1 0 24012 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__B
timestamp 1644511149
transform 1 0 25208 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1644511149
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__B
timestamp 1644511149
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__C
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A1
timestamp 1644511149
transform -1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1644511149
transform -1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A0
timestamp 1644511149
transform -1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__S
timestamp 1644511149
transform 1 0 7544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A0
timestamp 1644511149
transform -1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__S
timestamp 1644511149
transform 1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__B
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A1
timestamp 1644511149
transform -1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1644511149
transform -1 0 25208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A0
timestamp 1644511149
transform -1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__S
timestamp 1644511149
transform -1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A0
timestamp 1644511149
transform -1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__S
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A0
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__S
timestamp 1644511149
transform 1 0 11960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1644511149
transform 1 0 8004 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A0
timestamp 1644511149
transform -1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A0
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A0
timestamp 1644511149
transform 1 0 4968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A0
timestamp 1644511149
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A0
timestamp 1644511149
transform 1 0 4968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1644511149
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A0
timestamp 1644511149
transform 1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1644511149
transform 1 0 8372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A0
timestamp 1644511149
transform 1 0 7912 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A0
timestamp 1644511149
transform 1 0 4968 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__S
timestamp 1644511149
transform -1 0 8740 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__A1
timestamp 1644511149
transform -1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__A2
timestamp 1644511149
transform -1 0 23644 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__B1_N
timestamp 1644511149
transform 1 0 21160 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__A1
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1644511149
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1644511149
transform -1 0 24380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1644511149
transform 1 0 23736 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1644511149
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1644511149
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1644511149
transform 1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1644511149
transform 1 0 4784 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1644511149
transform 1 0 10856 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1644511149
transform 1 0 10488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1644511149
transform 1 0 16836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1644511149
transform 1 0 4508 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1644511149
transform 1 0 9476 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1644511149
transform 1 0 4508 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1644511149
transform 1 0 10856 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1644511149
transform -1 0 18584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1644511149
transform 1 0 10856 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1644511149
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1644511149
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_wb_clk_i_A
timestamp 1644511149
transform -1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_wb_clk_i_A
timestamp 1644511149
transform -1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_wb_clk_i_A
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_wb_clk_i_A
timestamp 1644511149
transform 1 0 15456 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 35512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 34960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 37536 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 36800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 36800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 36800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 37444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 37444 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 37444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 37536 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 36800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 36340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 36800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 37444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 37444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 36892 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 36800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 37444 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 36156 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 35604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 34040 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 36892 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 36800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 36800 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 35604 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 36800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 35972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 36800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 36800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 36800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform -1 0 36340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 4048 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 2300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 2944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 2852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 2944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 2208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 2668 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 2852 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 3312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 2852 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 2852 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 2944 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 3312 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 2944 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 2944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 2668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 2852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 2668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 2300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 2300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1644511149
transform -1 0 2668 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1644511149
transform -1 0 3220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1644511149
transform -1 0 2300 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1644511149
transform -1 0 3404 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1644511149
transform -1 0 2300 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1644511149
transform -1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1644511149
transform -1 0 3404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1644511149
transform -1 0 2668 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1644511149
transform -1 0 2668 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1644511149
transform -1 0 2300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1644511149
transform -1 0 2668 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1644511149
transform -1 0 2300 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1644511149
transform -1 0 3220 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1644511149
transform -1 0 4876 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1644511149
transform -1 0 5428 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1644511149
transform -1 0 5428 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1644511149
transform -1 0 2668 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1644511149
transform -1 0 6532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1644511149
transform -1 0 7084 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1644511149
transform -1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1644511149
transform -1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1644511149
transform -1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1644511149
transform -1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1644511149
transform -1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1644511149
transform -1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1644511149
transform -1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1644511149
transform -1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1644511149
transform -1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1644511149
transform -1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1644511149
transform -1 0 2852 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1644511149
transform -1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1644511149
transform -1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1644511149
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output160_A
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output162_A
timestamp 1644511149
transform -1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output163_A
timestamp 1644511149
transform -1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1644511149
transform 1 0 3312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1644511149
transform -1 0 2852 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output166_A
timestamp 1644511149
transform -1 0 3404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1644511149
transform -1 0 3220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1644511149
transform 1 0 2576 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1644511149
transform -1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1644511149
transform -1 0 2852 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1644511149
transform -1 0 2852 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1644511149
transform -1 0 3404 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1644511149
transform 1 0 3312 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output177_A
timestamp 1644511149
transform -1 0 4600 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1644511149
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output188_A
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output189_A
timestamp 1644511149
transform -1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1644511149
transform -1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1644511149
transform -1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output192_A
timestamp 1644511149
transform -1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_372
timestamp 1644511149
transform 1 0 35328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_380
timestamp 1644511149
transform 1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_86 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_97
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1644511149
transform 1 0 34684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1644511149
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1644511149
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_381
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_31
timestamp 1644511149
transform 1 0 3956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_95
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_102
timestamp 1644511149
transform 1 0 10488 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_124
timestamp 1644511149
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_173
timestamp 1644511149
transform 1 0 17020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_185
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1644511149
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_213
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_225
timestamp 1644511149
transform 1 0 21804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_237
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1644511149
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_256
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_262
timestamp 1644511149
transform 1 0 25208 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_274
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_282
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_294
timestamp 1644511149
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1644511149
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_318
timestamp 1644511149
transform 1 0 30360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_330
timestamp 1644511149
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_342
timestamp 1644511149
transform 1 0 32568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp 1644511149
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1644511149
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_383
timestamp 1644511149
transform 1 0 36340 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_387
timestamp 1644511149
transform 1 0 36708 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1644511149
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_26
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_34
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_59
timestamp 1644511149
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_71
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_83
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_95
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1644511149
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_175
timestamp 1644511149
transform 1 0 17204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1644511149
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1644511149
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_234
timestamp 1644511149
transform 1 0 22632 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_241
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_268
timestamp 1644511149
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_297
timestamp 1644511149
transform 1 0 28428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_303
timestamp 1644511149
transform 1 0 28980 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1644511149
transform 1 0 30360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_347
timestamp 1644511149
transform 1 0 33028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_356
timestamp 1644511149
transform 1 0 33856 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_368
timestamp 1644511149
transform 1 0 34960 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_376
timestamp 1644511149
transform 1 0 35696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1644511149
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_11
timestamp 1644511149
transform 1 0 2116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 1644511149
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_37
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_45
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_61
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_73
timestamp 1644511149
transform 1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1644511149
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_260
timestamp 1644511149
transform 1 0 25024 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_272
timestamp 1644511149
transform 1 0 26128 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_286
timestamp 1644511149
transform 1 0 27416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_295
timestamp 1644511149
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_348
timestamp 1644511149
transform 1 0 33120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_383
timestamp 1644511149
transform 1 0 36340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_393
timestamp 1644511149
transform 1 0 37260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1644511149
transform 1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1644511149
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1644511149
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_315
timestamp 1644511149
transform 1 0 30084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_327
timestamp 1644511149
transform 1 0 31188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_339
timestamp 1644511149
transform 1 0 32292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_351
timestamp 1644511149
transform 1 0 33396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1644511149
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_370
timestamp 1644511149
transform 1 0 35144 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_382
timestamp 1644511149
transform 1 0 36248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_388
timestamp 1644511149
transform 1 0 36800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1644511149
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1644511149
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1644511149
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_120
timestamp 1644511149
transform 1 0 12144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1644511149
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1644511149
transform 1 0 13892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1644511149
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_245
timestamp 1644511149
transform 1 0 23644 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1644511149
transform 1 0 23920 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1644511149
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1644511149
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_353
timestamp 1644511149
transform 1 0 33580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_365
timestamp 1644511149
transform 1 0 34684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_377
timestamp 1644511149
transform 1 0 35788 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1644511149
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_11
timestamp 1644511149
transform 1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_17
timestamp 1644511149
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1644511149
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp 1644511149
transform 1 0 7452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_72
timestamp 1644511149
transform 1 0 7728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1644511149
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_157
timestamp 1644511149
transform 1 0 15548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1644511149
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1644511149
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp 1644511149
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_285
timestamp 1644511149
transform 1 0 27324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_294
timestamp 1644511149
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1644511149
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 1644511149
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_388
timestamp 1644511149
transform 1 0 36800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 1644511149
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1644511149
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1644511149
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1644511149
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp 1644511149
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_73
timestamp 1644511149
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1644511149
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_191
timestamp 1644511149
transform 1 0 18676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_203
timestamp 1644511149
transform 1 0 19780 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_206
timestamp 1644511149
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1644511149
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_323
timestamp 1644511149
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1644511149
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_342
timestamp 1644511149
transform 1 0 32568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1644511149
transform 1 0 33672 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_366
timestamp 1644511149
transform 1 0 34776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_378
timestamp 1644511149
transform 1 0 35880 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_384
timestamp 1644511149
transform 1 0 36432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1644511149
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1644511149
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_200
timestamp 1644511149
transform 1 0 19504 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_222
timestamp 1644511149
transform 1 0 21528 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_234
timestamp 1644511149
transform 1 0 22632 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_246
timestamp 1644511149
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_315
timestamp 1644511149
transform 1 0 30084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_327
timestamp 1644511149
transform 1 0 31188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_339
timestamp 1644511149
transform 1 0 32292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_351
timestamp 1644511149
transform 1 0 33396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_393
timestamp 1644511149
transform 1 0 37260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1644511149
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1644511149
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1644511149
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1644511149
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1644511149
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_286
timestamp 1644511149
transform 1 0 27416 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_298
timestamp 1644511149
transform 1 0 28520 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1644511149
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1644511149
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_357
timestamp 1644511149
transform 1 0 33948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_366
timestamp 1644511149
transform 1 0 34776 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_378
timestamp 1644511149
transform 1 0 35880 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_384
timestamp 1644511149
transform 1 0 36432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1644511149
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_395
timestamp 1644511149
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1644511149
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1644511149
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_52
timestamp 1644511149
transform 1 0 5888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_64
timestamp 1644511149
transform 1 0 6992 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_341
timestamp 1644511149
transform 1 0 32476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_354
timestamp 1644511149
transform 1 0 33672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1644511149
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_385
timestamp 1644511149
transform 1 0 36524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1644511149
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1644511149
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1644511149
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_26
timestamp 1644511149
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_38
timestamp 1644511149
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1644511149
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_255
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_267
timestamp 1644511149
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_283
timestamp 1644511149
transform 1 0 27140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_297
timestamp 1644511149
transform 1 0 28428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_309
timestamp 1644511149
transform 1 0 29532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_313
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1644511149
transform 1 0 31004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_342
timestamp 1644511149
transform 1 0 32568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_350
timestamp 1644511149
transform 1 0 33304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_355
timestamp 1644511149
transform 1 0 33764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_364
timestamp 1644511149
transform 1 0 34592 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_376
timestamp 1644511149
transform 1 0 35696 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_384
timestamp 1644511149
transform 1 0 36432 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1644511149
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1644511149
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1644511149
transform 1 0 9108 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1644511149
transform 1 0 10212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1644511149
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1644511149
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1644511149
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1644511149
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1644511149
transform 1 0 14444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_173
timestamp 1644511149
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_178
timestamp 1644511149
transform 1 0 17480 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1644511149
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_237
timestamp 1644511149
transform 1 0 22908 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_242
timestamp 1644511149
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1644511149
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1644511149
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1644511149
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_317
timestamp 1644511149
transform 1 0 30268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_329
timestamp 1644511149
transform 1 0 31372 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_341
timestamp 1644511149
transform 1 0 32476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_353
timestamp 1644511149
transform 1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1644511149
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_379
timestamp 1644511149
transform 1 0 35972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_386
timestamp 1644511149
transform 1 0 36616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_393
timestamp 1644511149
transform 1 0 37260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1644511149
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1644511149
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1644511149
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_155
timestamp 1644511149
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1644511149
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_200
timestamp 1644511149
transform 1 0 19504 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_212
timestamp 1644511149
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_258
timestamp 1644511149
transform 1 0 24840 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_270
timestamp 1644511149
transform 1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1644511149
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1644511149
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1644511149
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_18
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1644511149
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 1644511149
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1644511149
transform 1 0 10488 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1644511149
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_126
timestamp 1644511149
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1644511149
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1644511149
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_230
timestamp 1644511149
transform 1 0 22264 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1644511149
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1644511149
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_368
timestamp 1644511149
transform 1 0 34960 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_380
timestamp 1644511149
transform 1 0 36064 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_388
timestamp 1644511149
transform 1 0 36800 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1644511149
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_19
timestamp 1644511149
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1644511149
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_85
timestamp 1644511149
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_97
timestamp 1644511149
transform 1 0 10028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_157
timestamp 1644511149
transform 1 0 15548 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_256
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_268
timestamp 1644511149
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1644511149
transform 1 0 32476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_344
timestamp 1644511149
transform 1 0 32752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_356
timestamp 1644511149
transform 1 0 33856 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_368
timestamp 1644511149
transform 1 0 34960 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_380
timestamp 1644511149
transform 1 0 36064 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_384
timestamp 1644511149
transform 1 0 36432 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1644511149
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1644511149
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_7
timestamp 1644511149
transform 1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_14
timestamp 1644511149
transform 1 0 2392 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_20
timestamp 1644511149
transform 1 0 2944 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_38
timestamp 1644511149
transform 1 0 4600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1644511149
transform 1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1644511149
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1644511149
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_148
timestamp 1644511149
transform 1 0 14720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_160
timestamp 1644511149
transform 1 0 15824 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_172
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_184
timestamp 1644511149
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_237
timestamp 1644511149
transform 1 0 22908 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1644511149
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1644511149
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1644511149
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1644511149
transform 1 0 29992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_328
timestamp 1644511149
transform 1 0 31280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_336
timestamp 1644511149
transform 1 0 32016 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_340
timestamp 1644511149
transform 1 0 32384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_349
timestamp 1644511149
transform 1 0 33212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1644511149
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_385
timestamp 1644511149
transform 1 0 36524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_397
timestamp 1644511149
transform 1 0 37628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1644511149
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_11
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_36
timestamp 1644511149
transform 1 0 4416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1644511149
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1644511149
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 1644511149
transform 1 0 14076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1644511149
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1644511149
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1644511149
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_342
timestamp 1644511149
transform 1 0 32568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_351
timestamp 1644511149
transform 1 0 33396 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_363
timestamp 1644511149
transform 1 0 34500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_375
timestamp 1644511149
transform 1 0 35604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1644511149
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1644511149
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1644511149
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1644511149
transform 1 0 25300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_275
timestamp 1644511149
transform 1 0 26404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_287
timestamp 1644511149
transform 1 0 27508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1644511149
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_383
timestamp 1644511149
transform 1 0 36340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_390
timestamp 1644511149
transform 1 0 36984 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_398
timestamp 1644511149
transform 1 0 37720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1644511149
transform 1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1644511149
transform 1 0 2668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_23
timestamp 1644511149
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_35
timestamp 1644511149
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1644511149
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1644511149
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1644511149
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1644511149
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1644511149
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1644511149
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1644511149
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1644511149
transform 1 0 23092 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_245
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_255
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_267
timestamp 1644511149
transform 1 0 25668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_294
timestamp 1644511149
transform 1 0 28152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_306
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_318
timestamp 1644511149
transform 1 0 30360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_343
timestamp 1644511149
transform 1 0 32660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_352
timestamp 1644511149
transform 1 0 33488 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_364
timestamp 1644511149
transform 1 0 34592 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_376
timestamp 1644511149
transform 1 0 35696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_384
timestamp 1644511149
transform 1 0 36432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1644511149
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_396
timestamp 1644511149
transform 1 0 37536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1644511149
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1644511149
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1644511149
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1644511149
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1644511149
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1644511149
transform 1 0 24840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_270
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_278
timestamp 1644511149
transform 1 0 26680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_285
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_293
timestamp 1644511149
transform 1 0 28060 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_313
timestamp 1644511149
transform 1 0 29900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_337
timestamp 1644511149
transform 1 0 32108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_341
timestamp 1644511149
transform 1 0 32476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_344
timestamp 1644511149
transform 1 0 32752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1644511149
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1644511149
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_385
timestamp 1644511149
transform 1 0 36524 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_388
timestamp 1644511149
transform 1 0 36800 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_395
timestamp 1644511149
transform 1 0 37444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_17
timestamp 1644511149
transform 1 0 2668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_23
timestamp 1644511149
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_35
timestamp 1644511149
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1644511149
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_68
timestamp 1644511149
transform 1 0 7360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_80
timestamp 1644511149
transform 1 0 8464 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_92
timestamp 1644511149
transform 1 0 9568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1644511149
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_131
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_143
timestamp 1644511149
transform 1 0 14260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_155
timestamp 1644511149
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_179
timestamp 1644511149
transform 1 0 17572 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_187
timestamp 1644511149
transform 1 0 18308 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_204
timestamp 1644511149
transform 1 0 19872 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_247
timestamp 1644511149
transform 1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_251
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_255
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_345
timestamp 1644511149
transform 1 0 32844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_353
timestamp 1644511149
transform 1 0 33580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_365
timestamp 1644511149
transform 1 0 34684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_381
timestamp 1644511149
transform 1 0 36156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1644511149
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1644511149
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1644511149
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_31
timestamp 1644511149
transform 1 0 3956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_43
timestamp 1644511149
transform 1 0 5060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_55
timestamp 1644511149
transform 1 0 6164 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1644511149
transform 1 0 9108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1644511149
transform 1 0 10212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_118
timestamp 1644511149
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1644511149
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1644511149
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_172
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_383
timestamp 1644511149
transform 1 0 36340 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_395
timestamp 1644511149
transform 1 0 37444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_11
timestamp 1644511149
transform 1 0 2116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1644511149
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_23
timestamp 1644511149
transform 1 0 3220 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_29
timestamp 1644511149
transform 1 0 3772 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_35
timestamp 1644511149
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1644511149
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1644511149
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_85
timestamp 1644511149
transform 1 0 8924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_97
timestamp 1644511149
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1644511149
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_299
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_308
timestamp 1644511149
transform 1 0 29440 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_316
timestamp 1644511149
transform 1 0 30176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_321
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1644511149
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_379
timestamp 1644511149
transform 1 0 35972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1644511149
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1644511149
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1644511149
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1644511149
transform 1 0 4600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1644511149
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1644511149
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_325
timestamp 1644511149
transform 1 0 31004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_337
timestamp 1644511149
transform 1 0 32108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_349
timestamp 1644511149
transform 1 0 33212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1644511149
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_385
timestamp 1644511149
transform 1 0 36524 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_391
timestamp 1644511149
transform 1 0 37076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1644511149
transform 1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1644511149
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_17
timestamp 1644511149
transform 1 0 2668 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_41
timestamp 1644511149
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1644511149
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_77
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_89
timestamp 1644511149
transform 1 0 9292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_101
timestamp 1644511149
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1644511149
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_131
timestamp 1644511149
transform 1 0 13156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_145
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 1644511149
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1644511149
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1644511149
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1644511149
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_299
timestamp 1644511149
transform 1 0 28612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_365
timestamp 1644511149
transform 1 0 34684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_377
timestamp 1644511149
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_395
timestamp 1644511149
transform 1 0 37444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1644511149
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1644511149
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_31
timestamp 1644511149
transform 1 0 3956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_43
timestamp 1644511149
transform 1 0 5060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_55
timestamp 1644511149
transform 1 0 6164 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_67
timestamp 1644511149
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1644511149
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1644511149
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_220
timestamp 1644511149
transform 1 0 21344 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_232
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1644511149
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_281
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_293
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1644511149
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_312
timestamp 1644511149
transform 1 0 29808 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_324
timestamp 1644511149
transform 1 0 30912 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_336
timestamp 1644511149
transform 1 0 32016 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_348
timestamp 1644511149
transform 1 0 33120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1644511149
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_393
timestamp 1644511149
transform 1 0 37260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_396
timestamp 1644511149
transform 1 0 37536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_14
timestamp 1644511149
transform 1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_20
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1644511149
transform 1 0 16928 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1644511149
transform 1 0 19136 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1644511149
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_230
timestamp 1644511149
transform 1 0 22264 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_242
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_254
timestamp 1644511149
transform 1 0 24472 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_266
timestamp 1644511149
transform 1 0 25576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1644511149
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1644511149
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_311
timestamp 1644511149
transform 1 0 29716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_340
timestamp 1644511149
transform 1 0 32384 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_352
timestamp 1644511149
transform 1 0 33488 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_362
timestamp 1644511149
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_374
timestamp 1644511149
transform 1 0 35512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_381
timestamp 1644511149
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1644511149
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_17
timestamp 1644511149
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1644511149
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1644511149
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1644511149
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_279
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_291
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1644511149
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1644511149
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_388
timestamp 1644511149
transform 1 0 36800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_395
timestamp 1644511149
transform 1 0 37444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1644511149
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_19
timestamp 1644511149
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_116
timestamp 1644511149
transform 1 0 11776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_140
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_152
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_239
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_251
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_263
timestamp 1644511149
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1644511149
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_311
timestamp 1644511149
transform 1 0 29716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_320
timestamp 1644511149
transform 1 0 30544 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1644511149
transform 1 0 32660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_355
timestamp 1644511149
transform 1 0 33764 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_367
timestamp 1644511149
transform 1 0 34868 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_377
timestamp 1644511149
transform 1 0 35788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_398
timestamp 1644511149
transform 1 0 37720 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1644511149
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1644511149
transform 1 0 2668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1644511149
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_61
timestamp 1644511149
transform 1 0 6716 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1644511149
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1644511149
transform 1 0 9108 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_99
timestamp 1644511149
transform 1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_104
timestamp 1644511149
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_124
timestamp 1644511149
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_229
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_240
timestamp 1644511149
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_373
timestamp 1644511149
transform 1 0 35420 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_385
timestamp 1644511149
transform 1 0 36524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_394
timestamp 1644511149
transform 1 0 37352 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_398
timestamp 1644511149
transform 1 0 37720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1644511149
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_7
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_14
timestamp 1644511149
transform 1 0 2392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_26
timestamp 1644511149
transform 1 0 3496 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_38
timestamp 1644511149
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1644511149
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1644511149
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_71
timestamp 1644511149
transform 1 0 7636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_83
timestamp 1644511149
transform 1 0 8740 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_95
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1644511149
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1644511149
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1644511149
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_309
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_312
timestamp 1644511149
transform 1 0 29808 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1644511149
transform 1 0 32660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1644511149
transform 1 0 33764 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1644511149
transform 1 0 34868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1644511149
transform 1 0 35972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1644511149
transform 1 0 38180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_11
timestamp 1644511149
transform 1 0 2116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_19
timestamp 1644511149
transform 1 0 2852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1644511149
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_38
timestamp 1644511149
transform 1 0 4600 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_50
timestamp 1644511149
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_62
timestamp 1644511149
transform 1 0 6808 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_67
timestamp 1644511149
transform 1 0 7268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1644511149
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1644511149
transform 1 0 15272 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1644511149
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1644511149
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_240
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_267
timestamp 1644511149
transform 1 0 25668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_385
timestamp 1644511149
transform 1 0 36524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_388
timestamp 1644511149
transform 1 0 36800 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_395
timestamp 1644511149
transform 1 0 37444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1644511149
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_33
timestamp 1644511149
transform 1 0 4140 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_152
timestamp 1644511149
transform 1 0 15088 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1644511149
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_235
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_247
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_265
timestamp 1644511149
transform 1 0 25484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_271
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_302
timestamp 1644511149
transform 1 0 28888 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_314
timestamp 1644511149
transform 1 0 29992 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_326
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1644511149
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1644511149
transform 1 0 38180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1644511149
transform 1 0 2116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_18
timestamp 1644511149
transform 1 0 2760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_167
timestamp 1644511149
transform 1 0 16468 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_173
timestamp 1644511149
transform 1 0 17020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_185
timestamp 1644511149
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1644511149
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1644511149
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_218
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_230
timestamp 1644511149
transform 1 0 22264 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_337
timestamp 1644511149
transform 1 0 32108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_341
timestamp 1644511149
transform 1 0 32476 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1644511149
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_373
timestamp 1644511149
transform 1 0 35420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_381
timestamp 1644511149
transform 1 0 36156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_385
timestamp 1644511149
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_388
timestamp 1644511149
transform 1 0 36800 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_395
timestamp 1644511149
transform 1 0 37444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp 1644511149
transform 1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_19
timestamp 1644511149
transform 1 0 2852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_25
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_37
timestamp 1644511149
transform 1 0 4508 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_49
timestamp 1644511149
transform 1 0 5612 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_89
timestamp 1644511149
transform 1 0 9292 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_248
timestamp 1644511149
transform 1 0 23920 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_256
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_311
timestamp 1644511149
transform 1 0 29716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_320
timestamp 1644511149
transform 1 0 30544 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_365
timestamp 1644511149
transform 1 0 34684 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_377
timestamp 1644511149
transform 1 0 35788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_395
timestamp 1644511149
transform 1 0 37444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1644511149
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_14
timestamp 1644511149
transform 1 0 2392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_20
timestamp 1644511149
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1644511149
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1644511149
transform 1 0 9200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_92
timestamp 1644511149
transform 1 0 9568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_217
timestamp 1644511149
transform 1 0 21068 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_222
timestamp 1644511149
transform 1 0 21528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_228
timestamp 1644511149
transform 1 0 22080 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_317
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_336
timestamp 1644511149
transform 1 0 32016 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_348
timestamp 1644511149
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_369
timestamp 1644511149
transform 1 0 35052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_386
timestamp 1644511149
transform 1 0 36616 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_395
timestamp 1644511149
transform 1 0 37444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_17
timestamp 1644511149
transform 1 0 2668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_309
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_312
timestamp 1644511149
transform 1 0 29808 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_324
timestamp 1644511149
transform 1 0 30912 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_369
timestamp 1644511149
transform 1 0 35052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_374
timestamp 1644511149
transform 1 0 35512 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1644511149
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_395
timestamp 1644511149
transform 1 0 37444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1644511149
transform 1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_6
timestamp 1644511149
transform 1 0 1656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_12
timestamp 1644511149
transform 1 0 2208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp 1644511149
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1644511149
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_145
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_157
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_169
timestamp 1644511149
transform 1 0 16652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_181
timestamp 1644511149
transform 1 0 17756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1644511149
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_288
timestamp 1644511149
transform 1 0 27600 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_300
timestamp 1644511149
transform 1 0 28704 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_314
timestamp 1644511149
transform 1 0 29992 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_326
timestamp 1644511149
transform 1 0 31096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_330
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_334
timestamp 1644511149
transform 1 0 31832 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_346
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 1644511149
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_369
timestamp 1644511149
transform 1 0 35052 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_373
timestamp 1644511149
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_388
timestamp 1644511149
transform 1 0 36800 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1644511149
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_17
timestamp 1644511149
transform 1 0 2668 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1644511149
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1644511149
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_75
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1644511149
transform 1 0 17572 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_199
timestamp 1644511149
transform 1 0 19412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_211
timestamp 1644511149
transform 1 0 20516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1644511149
transform 1 0 24748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1644511149
transform 1 0 25852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1644511149
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_395
timestamp 1644511149
transform 1 0 37444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1644511149
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_14
timestamp 1644511149
transform 1 0 2392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_18
timestamp 1644511149
transform 1 0 2760 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp 1644511149
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_38
timestamp 1644511149
transform 1 0 4600 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1644511149
transform 1 0 5152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_56
timestamp 1644511149
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_60
timestamp 1644511149
transform 1 0 6624 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_70
timestamp 1644511149
transform 1 0 7544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1644511149
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_176
timestamp 1644511149
transform 1 0 17296 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1644511149
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_236
timestamp 1644511149
transform 1 0 22816 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_273
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1644511149
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1644511149
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_329
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_388
timestamp 1644511149
transform 1 0 36800 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_395
timestamp 1644511149
transform 1 0 37444 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1644511149
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_11
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_33
timestamp 1644511149
transform 1 0 4140 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_178
timestamp 1644511149
transform 1 0 17480 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_190
timestamp 1644511149
transform 1 0 18584 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1644511149
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1644511149
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_242
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_254
timestamp 1644511149
transform 1 0 24472 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_266
timestamp 1644511149
transform 1 0 25576 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1644511149
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_284
timestamp 1644511149
transform 1 0 27232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_296
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_304
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_313
timestamp 1644511149
transform 1 0 29900 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_325
timestamp 1644511149
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1644511149
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_369
timestamp 1644511149
transform 1 0 35052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_374
timestamp 1644511149
transform 1 0 35512 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_380
timestamp 1644511149
transform 1 0 36064 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1644511149
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1644511149
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_31
timestamp 1644511149
transform 1 0 3956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_43
timestamp 1644511149
transform 1 0 5060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_55
timestamp 1644511149
transform 1 0 6164 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1644511149
transform 1 0 7176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp 1644511149
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_117
timestamp 1644511149
transform 1 0 11868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_127
timestamp 1644511149
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_241
timestamp 1644511149
transform 1 0 23276 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_314
timestamp 1644511149
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_329
timestamp 1644511149
transform 1 0 31372 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_341
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_353
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 1644511149
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1644511149
transform 1 0 35328 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_384
timestamp 1644511149
transform 1 0 36432 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_392
timestamp 1644511149
transform 1 0 37168 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_396
timestamp 1644511149
transform 1 0 37536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1644511149
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_19
timestamp 1644511149
transform 1 0 2852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_25
timestamp 1644511149
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_37
timestamp 1644511149
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1644511149
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_132
timestamp 1644511149
transform 1 0 13248 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_144
timestamp 1644511149
transform 1 0 14352 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_156
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_265
timestamp 1644511149
transform 1 0 25484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1644511149
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1644511149
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1644511149
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1644511149
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1644511149
transform 1 0 9108 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1644511149
transform 1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_111
timestamp 1644511149
transform 1 0 11316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_120
timestamp 1644511149
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1644511149
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1644511149
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1644511149
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_18
timestamp 1644511149
transform 1 0 2760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_24
timestamp 1644511149
transform 1 0 3312 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_36
timestamp 1644511149
transform 1 0 4416 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 1644511149
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_179
timestamp 1644511149
transform 1 0 17572 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_199
timestamp 1644511149
transform 1 0 19412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_211
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_289
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_294
timestamp 1644511149
transform 1 0 28152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_306
timestamp 1644511149
transform 1 0 29256 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_318
timestamp 1644511149
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1644511149
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_380
timestamp 1644511149
transform 1 0 36064 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_398
timestamp 1644511149
transform 1 0 37720 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1644511149
transform 1 0 38456 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_7
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_13
timestamp 1644511149
transform 1 0 2300 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1644511149
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1644511149
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1644511149
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_226
timestamp 1644511149
transform 1 0 21896 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1644511149
transform 1 0 26036 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_280
timestamp 1644511149
transform 1 0 26864 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_292
timestamp 1644511149
transform 1 0 27968 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_385
timestamp 1644511149
transform 1 0 36524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_388
timestamp 1644511149
transform 1 0 36800 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_395
timestamp 1644511149
transform 1 0 37444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1644511149
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_19
timestamp 1644511149
transform 1 0 2852 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_25
timestamp 1644511149
transform 1 0 3404 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_37
timestamp 1644511149
transform 1 0 4508 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_49
timestamp 1644511149
transform 1 0 5612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_286
timestamp 1644511149
transform 1 0 27416 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_295
timestamp 1644511149
transform 1 0 28244 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_307
timestamp 1644511149
transform 1 0 29348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_319
timestamp 1644511149
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1644511149
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_369
timestamp 1644511149
transform 1 0 35052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_376
timestamp 1644511149
transform 1 0 35696 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_398
timestamp 1644511149
transform 1 0 37720 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1644511149
transform 1 0 38456 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_11
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_385
timestamp 1644511149
transform 1 0 36524 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_388
timestamp 1644511149
transform 1 0 36800 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_395
timestamp 1644511149
transform 1 0 37444 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_13
timestamp 1644511149
transform 1 0 2300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_19
timestamp 1644511149
transform 1 0 2852 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_25
timestamp 1644511149
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_37
timestamp 1644511149
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1644511149
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_286
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_292
timestamp 1644511149
transform 1 0 27968 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_296
timestamp 1644511149
transform 1 0 28336 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_308
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_320
timestamp 1644511149
transform 1 0 30544 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_386
timestamp 1644511149
transform 1 0 36616 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_395
timestamp 1644511149
transform 1 0 37444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_17
timestamp 1644511149
transform 1 0 2668 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_25
timestamp 1644511149
transform 1 0 3404 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_61
timestamp 1644511149
transform 1 0 6716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1644511149
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1644511149
transform 1 0 9108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1644511149
transform 1 0 10212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_111
timestamp 1644511149
transform 1 0 11316 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_126
timestamp 1644511149
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1644511149
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1644511149
transform 1 0 16560 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_226
timestamp 1644511149
transform 1 0 21896 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_238
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1644511149
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_353
timestamp 1644511149
transform 1 0 33580 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1644511149
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_373
timestamp 1644511149
transform 1 0 35420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_378
timestamp 1644511149
transform 1 0 35880 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_384
timestamp 1644511149
transform 1 0 36432 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_395
timestamp 1644511149
transform 1 0 37444 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1644511149
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_7
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_20
timestamp 1644511149
transform 1 0 2944 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_26
timestamp 1644511149
transform 1 0 3496 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_38
timestamp 1644511149
transform 1 0 4600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1644511149
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_65
timestamp 1644511149
transform 1 0 7084 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_77
timestamp 1644511149
transform 1 0 8188 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_83
timestamp 1644511149
transform 1 0 8740 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_95
timestamp 1644511149
transform 1 0 9844 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_103
timestamp 1644511149
transform 1 0 10580 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_130
timestamp 1644511149
transform 1 0 13064 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_142
timestamp 1644511149
transform 1 0 14168 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_154
timestamp 1644511149
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1644511149
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1644511149
transform 1 0 16928 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1644511149
transform 1 0 19136 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_208
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_216
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_230
timestamp 1644511149
transform 1 0 22264 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_238
timestamp 1644511149
transform 1 0 23000 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_284
timestamp 1644511149
transform 1 0 27232 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_290
timestamp 1644511149
transform 1 0 27784 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_302
timestamp 1644511149
transform 1 0 28888 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_314
timestamp 1644511149
transform 1 0 29992 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_326
timestamp 1644511149
transform 1 0 31096 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1644511149
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_377
timestamp 1644511149
transform 1 0 35788 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_383
timestamp 1644511149
transform 1 0 36340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1644511149
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_11
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_17
timestamp 1644511149
transform 1 0 2668 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1644511149
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_72
timestamp 1644511149
transform 1 0 7728 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_115
timestamp 1644511149
transform 1 0 11684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_119
timestamp 1644511149
transform 1 0 12052 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_131
timestamp 1644511149
transform 1 0 13156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_184
timestamp 1644511149
transform 1 0 18032 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1644511149
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_217
timestamp 1644511149
transform 1 0 21068 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_226
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_234
timestamp 1644511149
transform 1 0 22632 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1644511149
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_261
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_266
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_275
timestamp 1644511149
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_290
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_302
timestamp 1644511149
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_353
timestamp 1644511149
transform 1 0 33580 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_358
timestamp 1644511149
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_395
timestamp 1644511149
transform 1 0 37444 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1644511149
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_13
timestamp 1644511149
transform 1 0 2300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_20
timestamp 1644511149
transform 1 0 2944 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_26
timestamp 1644511149
transform 1 0 3496 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_38
timestamp 1644511149
transform 1 0 4600 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_50
timestamp 1644511149
transform 1 0 5704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_263
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1644511149
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_301
timestamp 1644511149
transform 1 0 28796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_307
timestamp 1644511149
transform 1 0 29348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_313
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_325
timestamp 1644511149
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1644511149
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_399
timestamp 1644511149
transform 1 0 37812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_11
timestamp 1644511149
transform 1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_18
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_284
timestamp 1644511149
transform 1 0 27232 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_296
timestamp 1644511149
transform 1 0 28336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_374
timestamp 1644511149
transform 1 0 35512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_380
timestamp 1644511149
transform 1 0 36064 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_386
timestamp 1644511149
transform 1 0 36616 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_396
timestamp 1644511149
transform 1 0 37536 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_340
timestamp 1644511149
transform 1 0 32384 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_352
timestamp 1644511149
transform 1 0 33488 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_364
timestamp 1644511149
transform 1 0 34592 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_376
timestamp 1644511149
transform 1 0 35696 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1644511149
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_395
timestamp 1644511149
transform 1 0 37444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_11
timestamp 1644511149
transform 1 0 2116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_17
timestamp 1644511149
transform 1 0 2668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1644511149
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_353
timestamp 1644511149
transform 1 0 33580 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_374
timestamp 1644511149
transform 1 0 35512 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_388
timestamp 1644511149
transform 1 0 36800 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_395
timestamp 1644511149
transform 1 0 37444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_11
timestamp 1644511149
transform 1 0 2116 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_20
timestamp 1644511149
transform 1 0 2944 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_26
timestamp 1644511149
transform 1 0 3496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_32
timestamp 1644511149
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_44
timestamp 1644511149
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_308
timestamp 1644511149
transform 1 0 29440 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_340
timestamp 1644511149
transform 1 0 32384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_352
timestamp 1644511149
transform 1 0 33488 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_364
timestamp 1644511149
transform 1 0 34592 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_376
timestamp 1644511149
transform 1 0 35696 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_384
timestamp 1644511149
transform 1 0 36432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_399
timestamp 1644511149
transform 1 0 37812 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_19
timestamp 1644511149
transform 1 0 2852 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1644511149
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1644511149
transform 1 0 4048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_38
timestamp 1644511149
transform 1 0 4600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_50
timestamp 1644511149
transform 1 0 5704 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_62
timestamp 1644511149
transform 1 0 6808 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_74
timestamp 1644511149
transform 1 0 7912 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1644511149
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_261
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_273
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_285
timestamp 1644511149
transform 1 0 27324 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1644511149
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_375
timestamp 1644511149
transform 1 0 35604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_381
timestamp 1644511149
transform 1 0 36156 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_388
timestamp 1644511149
transform 1 0 36800 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_395
timestamp 1644511149
transform 1 0 37444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_11
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_23
timestamp 1644511149
transform 1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_37
timestamp 1644511149
transform 1 0 4508 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_213
timestamp 1644511149
transform 1 0 20700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_227
timestamp 1644511149
transform 1 0 21988 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_239
timestamp 1644511149
transform 1 0 23092 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_247
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_250
timestamp 1644511149
transform 1 0 24104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_259
timestamp 1644511149
transform 1 0 24932 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_267
timestamp 1644511149
transform 1 0 25668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_271
timestamp 1644511149
transform 1 0 26036 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_275
timestamp 1644511149
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_309
timestamp 1644511149
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1644511149
transform 1 0 30360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1644511149
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_348
timestamp 1644511149
transform 1 0 33120 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_360
timestamp 1644511149
transform 1 0 34224 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_372
timestamp 1644511149
transform 1 0 35328 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_375
timestamp 1644511149
transform 1 0 35604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_379
timestamp 1644511149
transform 1 0 35972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_386
timestamp 1644511149
transform 1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_395
timestamp 1644511149
transform 1 0 37444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_11
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_32
timestamp 1644511149
transform 1 0 4048 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_39
timestamp 1644511149
transform 1 0 4692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_45
timestamp 1644511149
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_57
timestamp 1644511149
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_69
timestamp 1644511149
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1644511149
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_224
timestamp 1644511149
transform 1 0 21712 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1644511149
transform 1 0 23092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_256
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_269
timestamp 1644511149
transform 1 0 25852 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_273
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_280
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_292
timestamp 1644511149
transform 1 0 27968 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_318
timestamp 1644511149
transform 1 0 30360 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1644511149
transform 1 0 31188 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_339
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_349
timestamp 1644511149
transform 1 0 33212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_356
timestamp 1644511149
transform 1 0 33856 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_369
timestamp 1644511149
transform 1 0 35052 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_373
timestamp 1644511149
transform 1 0 35420 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_383
timestamp 1644511149
transform 1 0 36340 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_11
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_35
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_41
timestamp 1644511149
transform 1 0 4876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1644511149
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_258
timestamp 1644511149
transform 1 0 24840 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_264
timestamp 1644511149
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_313
timestamp 1644511149
transform 1 0 29900 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_319
timestamp 1644511149
transform 1 0 30452 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1644511149
transform 1 0 30728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1644511149
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_355
timestamp 1644511149
transform 1 0 33764 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_358
timestamp 1644511149
transform 1 0 34040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_365
timestamp 1644511149
transform 1 0 34684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_383
timestamp 1644511149
transform 1 0 36340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1644511149
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_19
timestamp 1644511149
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_33
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_47
timestamp 1644511149
transform 1 0 5428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1644511149
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_59
timestamp 1644511149
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_181
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1644511149
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_355
timestamp 1644511149
transform 1 0 33764 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_372
timestamp 1644511149
transform 1 0 35328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_380
timestamp 1644511149
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_388
timestamp 1644511149
transform 1 0 36800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _190_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _191_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _192_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _193_
timestamp 1644511149
transform 1 0 32752 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _194_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _195_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _196_
timestamp 1644511149
transform 1 0 33396 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1644511149
transform -1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _198_
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1644511149
transform -1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1644511149
transform -1 0 36800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _202_
timestamp 1644511149
transform 1 0 34132 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1644511149
transform -1 0 36892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1644511149
transform -1 0 32384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1644511149
transform 1 0 32752 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1644511149
transform -1 0 34960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1644511149
transform 1 0 32936 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1644511149
transform -1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _209_
timestamp 1644511149
transform 1 0 33120 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1644511149
transform -1 0 36984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _211_
timestamp 1644511149
transform 1 0 33028 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1644511149
transform -1 0 37536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _213_
timestamp 1644511149
transform 1 0 33120 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1644511149
transform -1 0 36800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1644511149
transform -1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 1644511149
transform 1 0 20884 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _217_
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _218_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _219_
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _220_
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _221_
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _222_
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _223_
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _225_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1644511149
transform -1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1644511149
transform -1 0 25208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _229_
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1644511149
transform -1 0 26496 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _231_
timestamp 1644511149
transform 1 0 23184 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1644511149
transform -1 0 26588 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _233_
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1644511149
transform -1 0 27232 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _235_
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1644511149
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _237_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _238_
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _239_
timestamp 1644511149
transform 1 0 23000 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _240_
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _241_
timestamp 1644511149
transform 1 0 23092 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _242_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _243_
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _245_
timestamp 1644511149
transform 1 0 22908 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 1644511149
transform 1 0 21252 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1644511149
transform -1 0 36800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _248_
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1644511149
transform -1 0 33120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _250_
timestamp 1644511149
transform 1 0 31188 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1644511149
transform -1 0 33580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _252_
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1644511149
transform -1 0 36800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _254_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _255_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 1644511149
transform -1 0 30268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _257_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 30360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _259_
timestamp 1644511149
transform -1 0 30360 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _261_
timestamp 1644511149
transform -1 0 30084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _263_
timestamp 1644511149
transform -1 0 30084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1644511149
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _265_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1644511149
transform -1 0 24564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 1644511149
transform -1 0 24564 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _268_
timestamp 1644511149
transform -1 0 23368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _269_
timestamp 1644511149
transform -1 0 24840 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _270_
timestamp 1644511149
transform -1 0 23736 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _271_
timestamp 1644511149
transform -1 0 24656 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _272_
timestamp 1644511149
transform -1 0 23368 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _273_
timestamp 1644511149
transform -1 0 25300 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _274_
timestamp 1644511149
transform -1 0 24564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _275_
timestamp 1644511149
transform -1 0 24840 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _276_
timestamp 1644511149
transform -1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1644511149
transform -1 0 35788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1644511149
transform -1 0 37720 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _279_
timestamp 1644511149
transform -1 0 36432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _280_
timestamp 1644511149
transform -1 0 36524 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _281_
timestamp 1644511149
transform -1 0 34684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _282_
timestamp 1644511149
transform -1 0 36156 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1644511149
transform -1 0 34408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _284_
timestamp 1644511149
transform -1 0 37720 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _285_
timestamp 1644511149
transform -1 0 35420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _286_
timestamp 1644511149
transform -1 0 37352 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _287_
timestamp 1644511149
transform -1 0 35788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1644511149
transform -1 0 35788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _289_
timestamp 1644511149
transform -1 0 36156 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _290_
timestamp 1644511149
transform -1 0 34684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 1644511149
transform -1 0 36616 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _292_
timestamp 1644511149
transform -1 0 35052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _293_
timestamp 1644511149
transform -1 0 36800 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _294_
timestamp 1644511149
transform -1 0 35052 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _295_
timestamp 1644511149
transform -1 0 36800 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _296_
timestamp 1644511149
transform -1 0 35512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _297_
timestamp 1644511149
transform -1 0 36616 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _298_
timestamp 1644511149
transform -1 0 35328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1644511149
transform -1 0 35880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _300_
timestamp 1644511149
transform -1 0 37720 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _301_
timestamp 1644511149
transform -1 0 36064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _302_
timestamp 1644511149
transform -1 0 37720 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _303_
timestamp 1644511149
transform -1 0 35696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _304_
timestamp 1644511149
transform -1 0 36616 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _305_
timestamp 1644511149
transform -1 0 34040 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _306_
timestamp 1644511149
transform -1 0 36340 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _307_
timestamp 1644511149
transform -1 0 34040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _308_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1644511149
transform 1 0 2668 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1644511149
transform -1 0 35512 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _311_
timestamp 1644511149
transform -1 0 35512 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _312_
timestamp 1644511149
transform -1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _313_
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1644511149
transform 1 0 2668 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _315_
timestamp 1644511149
transform -1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1644511149
transform 1 0 2944 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _317_
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _319_
timestamp 1644511149
transform 1 0 35788 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _321_
timestamp 1644511149
transform -1 0 21712 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform -1 0 4508 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp 1644511149
transform -1 0 22540 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform 1 0 4416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _325_
timestamp 1644511149
transform -1 0 20884 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1644511149
transform -1 0 4048 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _327_
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _328_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _329_
timestamp 1644511149
transform 1 0 27508 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _330_
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1644511149
transform -1 0 36708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _332_
timestamp 1644511149
transform 1 0 27784 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1644511149
transform -1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _334_
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1644511149
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _336_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1644511149
transform -1 0 37260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _338_
timestamp 1644511149
transform -1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1644511149
transform -1 0 27324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _340_
timestamp 1644511149
transform 1 0 28244 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1644511149
transform -1 0 36800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _342_
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1644511149
transform -1 0 37260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _344_
timestamp 1644511149
transform 1 0 28336 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1644511149
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _346_
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1644511149
transform -1 0 36340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _348_
timestamp 1644511149
transform 1 0 28152 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1644511149
transform -1 0 29900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1644511149
transform -1 0 29164 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _351_
timestamp 1644511149
transform 1 0 28980 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1644511149
transform -1 0 30636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _353_
timestamp 1644511149
transform 1 0 29256 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1644511149
transform -1 0 31004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1644511149
transform -1 0 32384 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _357_
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1644511149
transform -1 0 32660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _359_
timestamp 1644511149
transform 1 0 30176 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _360_
timestamp 1644511149
transform -1 0 32660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _361_
timestamp 1644511149
transform -1 0 28980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _362_
timestamp 1644511149
transform 1 0 30084 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _363_
timestamp 1644511149
transform -1 0 32476 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _364_
timestamp 1644511149
transform 1 0 29808 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _365_
timestamp 1644511149
transform -1 0 32016 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _366_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1644511149
transform -1 0 31832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _368_
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1644511149
transform -1 0 31740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _370_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1644511149
transform -1 0 31372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _373_
timestamp 1644511149
transform 1 0 26404 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp 1644511149
transform -1 0 28152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _375_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _376_
timestamp 1644511149
transform -1 0 28244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _377_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1644511149
transform -1 0 28336 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _379_
timestamp 1644511149
transform 1 0 25944 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1644511149
transform -1 0 27784 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _381_
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _382_
timestamp 1644511149
transform -1 0 27232 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1644511149
transform -1 0 29348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _384_
timestamp 1644511149
transform 1 0 29808 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1644511149
transform -1 0 32384 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _386_
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _387_
timestamp 1644511149
transform -1 0 32384 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _388_
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1644511149
transform -1 0 33120 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _390_
timestamp 1644511149
transform 1 0 29900 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _391_
timestamp 1644511149
transform -1 0 33212 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _392_
timestamp 1644511149
transform 1 0 30728 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _393_
timestamp 1644511149
transform -1 0 33856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _394_
timestamp 1644511149
transform 1 0 25024 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1644511149
transform -1 0 26864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp 1644511149
transform 1 0 24472 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1644511149
transform -1 0 26220 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _398_
timestamp 1644511149
transform 1 0 24380 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1644511149
transform -1 0 26404 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _400_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3036 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _401_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 15456 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _402_
timestamp 1644511149
transform 1 0 15824 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _403_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 1644511149
transform -1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1644511149
transform -1 0 18676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1644511149
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _407_
timestamp 1644511149
transform -1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _408_
timestamp 1644511149
transform -1 0 8372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1644511149
transform -1 0 7820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1644511149
transform -1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _412_
timestamp 1644511149
transform -1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _414_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _415_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25024 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1644511149
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _417_
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1644511149
transform -1 0 9844 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp 1644511149
transform -1 0 10488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1644511149
transform 1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _421_
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1644511149
transform -1 0 13340 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _423_
timestamp 1644511149
transform -1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _424_
timestamp 1644511149
transform -1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1644511149
transform -1 0 3312 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1644511149
transform -1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1644511149
transform -1 0 8188 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1644511149
transform -1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _430_
timestamp 1644511149
transform 1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp 1644511149
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1644511149
transform -1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _435_
timestamp 1644511149
transform 1 0 12788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1644511149
transform 1 0 11684 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1644511149
transform -1 0 11960 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _438_
timestamp 1644511149
transform -1 0 16928 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1644511149
transform -1 0 17572 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _440_
timestamp 1644511149
transform 1 0 16652 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _441_
timestamp 1644511149
transform -1 0 16928 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _442_
timestamp 1644511149
transform 1 0 11408 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _443_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _444_
timestamp 1644511149
transform -1 0 15272 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1644511149
transform -1 0 15088 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _446_
timestamp 1644511149
transform -1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1644511149
transform 1 0 6808 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1644511149
transform -1 0 7268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _450_
timestamp 1644511149
transform 1 0 2944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _451_
timestamp 1644511149
transform -1 0 8280 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _452_
timestamp 1644511149
transform -1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _454_
timestamp 1644511149
transform -1 0 7176 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _456_
timestamp 1644511149
transform 1 0 2852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _457_
timestamp 1644511149
transform -1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1644511149
transform -1 0 17480 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1644511149
transform -1 0 17296 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp 1644511149
transform 1 0 11960 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _461_
timestamp 1644511149
transform -1 0 12144 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1644511149
transform -1 0 16836 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _463_
timestamp 1644511149
transform -1 0 17480 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1644511149
transform -1 0 16560 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _465_
timestamp 1644511149
transform -1 0 16928 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1644511149
transform 1 0 11868 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp 1644511149
transform 1 0 11776 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1644511149
transform 1 0 7360 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1644511149
transform 1 0 7452 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _470_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _471_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _472_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _473_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1644511149
transform 1 0 20056 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _475_
timestamp 1644511149
transform 1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _476_
timestamp 1644511149
transform 1 0 14812 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _477_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _478_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24288 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _479_
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _480_
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _481_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _482_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _483_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _484_
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _485_
timestamp 1644511149
transform 1 0 6900 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _486_
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1644511149
transform 1 0 11684 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1644511149
transform 1 0 18400 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1644511149
transform 1 0 11040 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1644511149
transform -1 0 16468 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1644511149
transform 1 0 6900 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1644511149
transform 1 0 6992 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1644511149
transform 1 0 2668 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1644511149
transform 1 0 17940 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1644511149
transform 1 0 11776 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1644511149
transform 1 0 16560 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1644511149
transform 1 0 11592 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1644511149
transform 1 0 6992 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1644511149
transform -1 0 17020 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1644511149
transform -1 0 20884 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _505_
timestamp 1644511149
transform 1 0 36984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1644511149
transform -1 0 9660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1644511149
transform -1 0 9660 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform -1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 37168 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform -1 0 37444 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 37168 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 37168 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 37168 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 37168 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 37168 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 37904 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 37444 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 35880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform -1 0 37444 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 37168 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 37904 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 37260 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 37168 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 37168 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 36524 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform -1 0 35420 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform -1 0 34684 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1644511149
transform 1 0 37260 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 37168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 37260 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 36340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 37168 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 37904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 37168 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform -1 0 36156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform -1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1644511149
transform -1 0 2300 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform -1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1644511149
transform -1 0 2300 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform -1 0 2392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform -1 0 2760 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform -1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform -1 0 2392 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1644511149
transform -1 0 2300 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform -1 0 2760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform -1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform -1 0 2300 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1644511149
transform -1 0 2300 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform -1 0 2392 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform -1 0 2760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform -1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform -1 0 2760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform -1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform -1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform -1 0 2300 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1644511149
transform 1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input91
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input93
timestamp 1644511149
transform -1 0 2300 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1644511149
transform -1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1644511149
transform -1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1644511149
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 37812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 37812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 37812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 37812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 37812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 37812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 37812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 37812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 37812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 37812 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 37812 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 37812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 37812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 37812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 37812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 37812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1644511149
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1644511149
transform 1 0 37812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1644511149
transform 1 0 37812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1644511149
transform 1 0 37812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1644511149
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1644511149
transform 1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1644511149
transform 1 0 37812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1644511149
transform 1 0 37812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1644511149
transform 1 0 37076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform 1 0 37812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 37812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform 1 0 37076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 37812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 37812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 36432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 35696 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 34960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 35052 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform 1 0 33856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform 1 0 37812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform 1 0 37812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 37812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform 1 0 37812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform 1 0 37076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform -1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform -1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform -1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform -1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform -1 0 2852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform -1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform -1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform -1 0 2852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform -1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform -1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform -1 0 2484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform -1 0 2852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform -1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform -1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform -1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform -1 0 3036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform -1 0 2852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform -1 0 2852 0 -1 3264
box -38 -48 406 592
<< labels >>
rlabel metal3 s 39200 1368 40000 1488 6 peripheralBus_address[0]
port 0 nsew signal tristate
rlabel metal3 s 39200 15648 40000 15768 6 peripheralBus_address[10]
port 1 nsew signal tristate
rlabel metal3 s 39200 16872 40000 16992 6 peripheralBus_address[11]
port 2 nsew signal tristate
rlabel metal3 s 39200 18232 40000 18352 6 peripheralBus_address[12]
port 3 nsew signal tristate
rlabel metal3 s 39200 19456 40000 19576 6 peripheralBus_address[13]
port 4 nsew signal tristate
rlabel metal3 s 39200 20680 40000 20800 6 peripheralBus_address[14]
port 5 nsew signal tristate
rlabel metal3 s 39200 21904 40000 22024 6 peripheralBus_address[15]
port 6 nsew signal tristate
rlabel metal3 s 39200 23264 40000 23384 6 peripheralBus_address[16]
port 7 nsew signal tristate
rlabel metal3 s 39200 24488 40000 24608 6 peripheralBus_address[17]
port 8 nsew signal tristate
rlabel metal3 s 39200 25712 40000 25832 6 peripheralBus_address[18]
port 9 nsew signal tristate
rlabel metal3 s 39200 27072 40000 27192 6 peripheralBus_address[19]
port 10 nsew signal tristate
rlabel metal3 s 39200 3000 40000 3120 6 peripheralBus_address[1]
port 11 nsew signal tristate
rlabel metal3 s 39200 28296 40000 28416 6 peripheralBus_address[20]
port 12 nsew signal tristate
rlabel metal3 s 39200 29520 40000 29640 6 peripheralBus_address[21]
port 13 nsew signal tristate
rlabel metal3 s 39200 30744 40000 30864 6 peripheralBus_address[22]
port 14 nsew signal tristate
rlabel metal3 s 39200 32104 40000 32224 6 peripheralBus_address[23]
port 15 nsew signal tristate
rlabel metal3 s 39200 4768 40000 4888 6 peripheralBus_address[2]
port 16 nsew signal tristate
rlabel metal3 s 39200 6400 40000 6520 6 peripheralBus_address[3]
port 17 nsew signal tristate
rlabel metal3 s 39200 8032 40000 8152 6 peripheralBus_address[4]
port 18 nsew signal tristate
rlabel metal3 s 39200 9392 40000 9512 6 peripheralBus_address[5]
port 19 nsew signal tristate
rlabel metal3 s 39200 10616 40000 10736 6 peripheralBus_address[6]
port 20 nsew signal tristate
rlabel metal3 s 39200 11840 40000 11960 6 peripheralBus_address[7]
port 21 nsew signal tristate
rlabel metal3 s 39200 13064 40000 13184 6 peripheralBus_address[8]
port 22 nsew signal tristate
rlabel metal3 s 39200 14424 40000 14544 6 peripheralBus_address[9]
port 23 nsew signal tristate
rlabel metal3 s 39200 144 40000 264 6 peripheralBus_busy
port 24 nsew signal input
rlabel metal3 s 39200 1776 40000 1896 6 peripheralBus_byteSelect[0]
port 25 nsew signal tristate
rlabel metal3 s 39200 3408 40000 3528 6 peripheralBus_byteSelect[1]
port 26 nsew signal tristate
rlabel metal3 s 39200 5176 40000 5296 6 peripheralBus_byteSelect[2]
port 27 nsew signal tristate
rlabel metal3 s 39200 6808 40000 6928 6 peripheralBus_byteSelect[3]
port 28 nsew signal tristate
rlabel metal3 s 39200 2184 40000 2304 6 peripheralBus_dataRead[0]
port 29 nsew signal input
rlabel metal3 s 39200 16056 40000 16176 6 peripheralBus_dataRead[10]
port 30 nsew signal input
rlabel metal3 s 39200 17280 40000 17400 6 peripheralBus_dataRead[11]
port 31 nsew signal input
rlabel metal3 s 39200 18640 40000 18760 6 peripheralBus_dataRead[12]
port 32 nsew signal input
rlabel metal3 s 39200 19864 40000 19984 6 peripheralBus_dataRead[13]
port 33 nsew signal input
rlabel metal3 s 39200 21088 40000 21208 6 peripheralBus_dataRead[14]
port 34 nsew signal input
rlabel metal3 s 39200 22448 40000 22568 6 peripheralBus_dataRead[15]
port 35 nsew signal input
rlabel metal3 s 39200 23672 40000 23792 6 peripheralBus_dataRead[16]
port 36 nsew signal input
rlabel metal3 s 39200 24896 40000 25016 6 peripheralBus_dataRead[17]
port 37 nsew signal input
rlabel metal3 s 39200 26120 40000 26240 6 peripheralBus_dataRead[18]
port 38 nsew signal input
rlabel metal3 s 39200 27480 40000 27600 6 peripheralBus_dataRead[19]
port 39 nsew signal input
rlabel metal3 s 39200 3816 40000 3936 6 peripheralBus_dataRead[1]
port 40 nsew signal input
rlabel metal3 s 39200 28704 40000 28824 6 peripheralBus_dataRead[20]
port 41 nsew signal input
rlabel metal3 s 39200 29928 40000 30048 6 peripheralBus_dataRead[21]
port 42 nsew signal input
rlabel metal3 s 39200 31288 40000 31408 6 peripheralBus_dataRead[22]
port 43 nsew signal input
rlabel metal3 s 39200 32512 40000 32632 6 peripheralBus_dataRead[23]
port 44 nsew signal input
rlabel metal3 s 39200 33328 40000 33448 6 peripheralBus_dataRead[24]
port 45 nsew signal input
rlabel metal3 s 39200 34144 40000 34264 6 peripheralBus_dataRead[25]
port 46 nsew signal input
rlabel metal3 s 39200 34960 40000 35080 6 peripheralBus_dataRead[26]
port 47 nsew signal input
rlabel metal3 s 39200 35912 40000 36032 6 peripheralBus_dataRead[27]
port 48 nsew signal input
rlabel metal3 s 39200 36728 40000 36848 6 peripheralBus_dataRead[28]
port 49 nsew signal input
rlabel metal3 s 39200 37544 40000 37664 6 peripheralBus_dataRead[29]
port 50 nsew signal input
rlabel metal3 s 39200 5584 40000 5704 6 peripheralBus_dataRead[2]
port 51 nsew signal input
rlabel metal3 s 39200 38360 40000 38480 6 peripheralBus_dataRead[30]
port 52 nsew signal input
rlabel metal3 s 39200 39176 40000 39296 6 peripheralBus_dataRead[31]
port 53 nsew signal input
rlabel metal3 s 39200 7216 40000 7336 6 peripheralBus_dataRead[3]
port 54 nsew signal input
rlabel metal3 s 39200 8440 40000 8560 6 peripheralBus_dataRead[4]
port 55 nsew signal input
rlabel metal3 s 39200 9800 40000 9920 6 peripheralBus_dataRead[5]
port 56 nsew signal input
rlabel metal3 s 39200 11024 40000 11144 6 peripheralBus_dataRead[6]
port 57 nsew signal input
rlabel metal3 s 39200 12248 40000 12368 6 peripheralBus_dataRead[7]
port 58 nsew signal input
rlabel metal3 s 39200 13608 40000 13728 6 peripheralBus_dataRead[8]
port 59 nsew signal input
rlabel metal3 s 39200 14832 40000 14952 6 peripheralBus_dataRead[9]
port 60 nsew signal input
rlabel metal3 s 39200 2592 40000 2712 6 peripheralBus_dataWrite[0]
port 61 nsew signal tristate
rlabel metal3 s 39200 16464 40000 16584 6 peripheralBus_dataWrite[10]
port 62 nsew signal tristate
rlabel metal3 s 39200 17688 40000 17808 6 peripheralBus_dataWrite[11]
port 63 nsew signal tristate
rlabel metal3 s 39200 19048 40000 19168 6 peripheralBus_dataWrite[12]
port 64 nsew signal tristate
rlabel metal3 s 39200 20272 40000 20392 6 peripheralBus_dataWrite[13]
port 65 nsew signal tristate
rlabel metal3 s 39200 21496 40000 21616 6 peripheralBus_dataWrite[14]
port 66 nsew signal tristate
rlabel metal3 s 39200 22856 40000 22976 6 peripheralBus_dataWrite[15]
port 67 nsew signal tristate
rlabel metal3 s 39200 24080 40000 24200 6 peripheralBus_dataWrite[16]
port 68 nsew signal tristate
rlabel metal3 s 39200 25304 40000 25424 6 peripheralBus_dataWrite[17]
port 69 nsew signal tristate
rlabel metal3 s 39200 26528 40000 26648 6 peripheralBus_dataWrite[18]
port 70 nsew signal tristate
rlabel metal3 s 39200 27888 40000 28008 6 peripheralBus_dataWrite[19]
port 71 nsew signal tristate
rlabel metal3 s 39200 4224 40000 4344 6 peripheralBus_dataWrite[1]
port 72 nsew signal tristate
rlabel metal3 s 39200 29112 40000 29232 6 peripheralBus_dataWrite[20]
port 73 nsew signal tristate
rlabel metal3 s 39200 30336 40000 30456 6 peripheralBus_dataWrite[21]
port 74 nsew signal tristate
rlabel metal3 s 39200 31696 40000 31816 6 peripheralBus_dataWrite[22]
port 75 nsew signal tristate
rlabel metal3 s 39200 32920 40000 33040 6 peripheralBus_dataWrite[23]
port 76 nsew signal tristate
rlabel metal3 s 39200 33736 40000 33856 6 peripheralBus_dataWrite[24]
port 77 nsew signal tristate
rlabel metal3 s 39200 34552 40000 34672 6 peripheralBus_dataWrite[25]
port 78 nsew signal tristate
rlabel metal3 s 39200 35368 40000 35488 6 peripheralBus_dataWrite[26]
port 79 nsew signal tristate
rlabel metal3 s 39200 36320 40000 36440 6 peripheralBus_dataWrite[27]
port 80 nsew signal tristate
rlabel metal3 s 39200 37136 40000 37256 6 peripheralBus_dataWrite[28]
port 81 nsew signal tristate
rlabel metal3 s 39200 37952 40000 38072 6 peripheralBus_dataWrite[29]
port 82 nsew signal tristate
rlabel metal3 s 39200 5992 40000 6112 6 peripheralBus_dataWrite[2]
port 83 nsew signal tristate
rlabel metal3 s 39200 38768 40000 38888 6 peripheralBus_dataWrite[30]
port 84 nsew signal tristate
rlabel metal3 s 39200 39584 40000 39704 6 peripheralBus_dataWrite[31]
port 85 nsew signal tristate
rlabel metal3 s 39200 7624 40000 7744 6 peripheralBus_dataWrite[3]
port 86 nsew signal tristate
rlabel metal3 s 39200 8848 40000 8968 6 peripheralBus_dataWrite[4]
port 87 nsew signal tristate
rlabel metal3 s 39200 10208 40000 10328 6 peripheralBus_dataWrite[5]
port 88 nsew signal tristate
rlabel metal3 s 39200 11432 40000 11552 6 peripheralBus_dataWrite[6]
port 89 nsew signal tristate
rlabel metal3 s 39200 12656 40000 12776 6 peripheralBus_dataWrite[7]
port 90 nsew signal tristate
rlabel metal3 s 39200 14016 40000 14136 6 peripheralBus_dataWrite[8]
port 91 nsew signal tristate
rlabel metal3 s 39200 15240 40000 15360 6 peripheralBus_dataWrite[9]
port 92 nsew signal tristate
rlabel metal3 s 39200 552 40000 672 6 peripheralBus_oe
port 93 nsew signal tristate
rlabel metal3 s 39200 960 40000 1080 6 peripheralBus_we
port 94 nsew signal tristate
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 95 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 95 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 96 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 97 nsew signal tristate
rlabel metal3 s 0 2864 800 2984 6 wb_adr_i[0]
port 98 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 wb_adr_i[10]
port 99 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 wb_adr_i[11]
port 100 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[12]
port 101 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[13]
port 102 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[14]
port 103 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[15]
port 104 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 wb_adr_i[16]
port 105 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wb_adr_i[17]
port 106 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 wb_adr_i[18]
port 107 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wb_adr_i[19]
port 108 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 wb_adr_i[1]
port 109 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 wb_adr_i[20]
port 110 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 wb_adr_i[21]
port 111 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 wb_adr_i[22]
port 112 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 wb_adr_i[23]
port 113 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wb_adr_i[2]
port 114 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wb_adr_i[3]
port 115 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 wb_adr_i[4]
port 116 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_adr_i[5]
port 117 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_adr_i[6]
port 118 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_adr_i[7]
port 119 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wb_adr_i[8]
port 120 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wb_adr_i[9]
port 121 nsew signal input
rlabel metal3 s 0 416 800 536 6 wb_clk_i
port 122 nsew signal input
rlabel metal3 s 0 824 800 944 6 wb_cyc_i
port 123 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 wb_data_i[0]
port 124 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wb_data_i[10]
port 125 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 wb_data_i[11]
port 126 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[12]
port 127 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[13]
port 128 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[14]
port 129 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[15]
port 130 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wb_data_i[16]
port 131 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 wb_data_i[17]
port 132 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wb_data_i[18]
port 133 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wb_data_i[19]
port 134 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 wb_data_i[1]
port 135 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_data_i[20]
port 136 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_data_i[21]
port 137 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_data_i[22]
port 138 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 wb_data_i[23]
port 139 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 wb_data_i[24]
port 140 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 wb_data_i[25]
port 141 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 wb_data_i[26]
port 142 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 wb_data_i[27]
port 143 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 wb_data_i[28]
port 144 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 wb_data_i[29]
port 145 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 wb_data_i[2]
port 146 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 wb_data_i[30]
port 147 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 wb_data_i[31]
port 148 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wb_data_i[3]
port 149 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_data_i[4]
port 150 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 wb_data_i[5]
port 151 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wb_data_i[6]
port 152 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 wb_data_i[7]
port 153 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wb_data_i[8]
port 154 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wb_data_i[9]
port 155 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 wb_data_o[0]
port 156 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 wb_data_o[10]
port 157 nsew signal tristate
rlabel metal3 s 0 18640 800 18760 6 wb_data_o[11]
port 158 nsew signal tristate
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[12]
port 159 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[13]
port 160 nsew signal tristate
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[14]
port 161 nsew signal tristate
rlabel metal3 s 0 23536 800 23656 6 wb_data_o[15]
port 162 nsew signal tristate
rlabel metal3 s 0 24760 800 24880 6 wb_data_o[16]
port 163 nsew signal tristate
rlabel metal3 s 0 25984 800 26104 6 wb_data_o[17]
port 164 nsew signal tristate
rlabel metal3 s 0 27072 800 27192 6 wb_data_o[18]
port 165 nsew signal tristate
rlabel metal3 s 0 28296 800 28416 6 wb_data_o[19]
port 166 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 wb_data_o[1]
port 167 nsew signal tristate
rlabel metal3 s 0 29520 800 29640 6 wb_data_o[20]
port 168 nsew signal tristate
rlabel metal3 s 0 30744 800 30864 6 wb_data_o[21]
port 169 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 wb_data_o[22]
port 170 nsew signal tristate
rlabel metal3 s 0 33192 800 33312 6 wb_data_o[23]
port 171 nsew signal tristate
rlabel metal3 s 0 34008 800 34128 6 wb_data_o[24]
port 172 nsew signal tristate
rlabel metal3 s 0 34824 800 34944 6 wb_data_o[25]
port 173 nsew signal tristate
rlabel metal3 s 0 35640 800 35760 6 wb_data_o[26]
port 174 nsew signal tristate
rlabel metal3 s 0 36456 800 36576 6 wb_data_o[27]
port 175 nsew signal tristate
rlabel metal3 s 0 37272 800 37392 6 wb_data_o[28]
port 176 nsew signal tristate
rlabel metal3 s 0 38088 800 38208 6 wb_data_o[29]
port 177 nsew signal tristate
rlabel metal3 s 0 6944 800 7064 6 wb_data_o[2]
port 178 nsew signal tristate
rlabel metal3 s 0 38904 800 39024 6 wb_data_o[30]
port 179 nsew signal tristate
rlabel metal3 s 0 39720 800 39840 6 wb_data_o[31]
port 180 nsew signal tristate
rlabel metal3 s 0 8576 800 8696 6 wb_data_o[3]
port 181 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 wb_data_o[4]
port 182 nsew signal tristate
rlabel metal3 s 0 11432 800 11552 6 wb_data_o[5]
port 183 nsew signal tristate
rlabel metal3 s 0 12656 800 12776 6 wb_data_o[6]
port 184 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 wb_data_o[7]
port 185 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 wb_data_o[8]
port 186 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 wb_data_o[9]
port 187 nsew signal tristate
rlabel metal3 s 0 1232 800 1352 6 wb_rst_i
port 188 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wb_sel_i[0]
port 189 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 wb_sel_i[1]
port 190 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wb_sel_i[2]
port 191 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 wb_sel_i[3]
port 192 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 wb_stall_o
port 193 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 wb_stb_i
port 194 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wb_we_i
port 195 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
