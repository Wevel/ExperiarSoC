magic
tech sky130A
magscale 1 2
timestamp 1651272821
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 38824 37584
<< metal2 >>
rect 9954 39200 10010 40000
rect 29918 39200 29974 40000
<< obsm2 >>
rect 1398 39144 9898 39681
rect 10066 39144 29862 39681
rect 30030 39144 38162 39681
rect 1398 303 38162 39144
<< metal3 >>
rect 0 39584 800 39704
rect 0 38904 800 39024
rect 0 38224 800 38344
rect 39200 37816 40000 37936
rect 0 37544 800 37664
rect 0 36864 800 36984
rect 0 36184 800 36304
rect 0 35504 800 35624
rect 0 34824 800 34944
rect 0 34144 800 34264
rect 39200 33872 40000 33992
rect 0 33464 800 33584
rect 0 32784 800 32904
rect 0 32104 800 32224
rect 0 31424 800 31544
rect 0 30744 800 30864
rect 0 30064 800 30184
rect 39200 29792 40000 29912
rect 0 29384 800 29504
rect 0 28704 800 28824
rect 0 28024 800 28144
rect 0 27344 800 27464
rect 0 26664 800 26784
rect 0 25984 800 26104
rect 39200 25848 40000 25968
rect 0 25304 800 25424
rect 0 24624 800 24744
rect 0 23944 800 24064
rect 0 23264 800 23384
rect 0 22584 800 22704
rect 0 21904 800 22024
rect 39200 21904 40000 22024
rect 0 21224 800 21344
rect 0 20544 800 20664
rect 0 19864 800 19984
rect 0 19184 800 19304
rect 0 18504 800 18624
rect 0 17824 800 17944
rect 39200 17824 40000 17944
rect 0 17144 800 17264
rect 0 16464 800 16584
rect 0 15784 800 15904
rect 0 15104 800 15224
rect 0 14424 800 14544
rect 0 13744 800 13864
rect 39200 13880 40000 14000
rect 0 13064 800 13184
rect 0 12384 800 12504
rect 0 11704 800 11824
rect 0 11024 800 11144
rect 0 10344 800 10464
rect 0 9664 800 9784
rect 39200 9800 40000 9920
rect 0 8984 800 9104
rect 0 8304 800 8424
rect 0 7624 800 7744
rect 0 6944 800 7064
rect 0 6264 800 6384
rect 39200 5856 40000 5976
rect 0 5584 800 5704
rect 0 4904 800 5024
rect 0 4224 800 4344
rect 0 3544 800 3664
rect 0 2864 800 2984
rect 0 2184 800 2304
rect 39200 1912 40000 2032
rect 0 1504 800 1624
rect 0 824 800 944
rect 0 280 800 400
<< obsm3 >>
rect 880 39504 39200 39677
rect 800 39104 39200 39504
rect 880 38824 39200 39104
rect 800 38424 39200 38824
rect 880 38144 39200 38424
rect 800 38016 39200 38144
rect 800 37744 39120 38016
rect 880 37736 39120 37744
rect 880 37464 39200 37736
rect 800 37064 39200 37464
rect 880 36784 39200 37064
rect 800 36384 39200 36784
rect 880 36104 39200 36384
rect 800 35704 39200 36104
rect 880 35424 39200 35704
rect 800 35024 39200 35424
rect 880 34744 39200 35024
rect 800 34344 39200 34744
rect 880 34072 39200 34344
rect 880 34064 39120 34072
rect 800 33792 39120 34064
rect 800 33664 39200 33792
rect 880 33384 39200 33664
rect 800 32984 39200 33384
rect 880 32704 39200 32984
rect 800 32304 39200 32704
rect 880 32024 39200 32304
rect 800 31624 39200 32024
rect 880 31344 39200 31624
rect 800 30944 39200 31344
rect 880 30664 39200 30944
rect 800 30264 39200 30664
rect 880 29992 39200 30264
rect 880 29984 39120 29992
rect 800 29712 39120 29984
rect 800 29584 39200 29712
rect 880 29304 39200 29584
rect 800 28904 39200 29304
rect 880 28624 39200 28904
rect 800 28224 39200 28624
rect 880 27944 39200 28224
rect 800 27544 39200 27944
rect 880 27264 39200 27544
rect 800 26864 39200 27264
rect 880 26584 39200 26864
rect 800 26184 39200 26584
rect 880 26048 39200 26184
rect 880 25904 39120 26048
rect 800 25768 39120 25904
rect 800 25504 39200 25768
rect 880 25224 39200 25504
rect 800 24824 39200 25224
rect 880 24544 39200 24824
rect 800 24144 39200 24544
rect 880 23864 39200 24144
rect 800 23464 39200 23864
rect 880 23184 39200 23464
rect 800 22784 39200 23184
rect 880 22504 39200 22784
rect 800 22104 39200 22504
rect 880 21824 39120 22104
rect 800 21424 39200 21824
rect 880 21144 39200 21424
rect 800 20744 39200 21144
rect 880 20464 39200 20744
rect 800 20064 39200 20464
rect 880 19784 39200 20064
rect 800 19384 39200 19784
rect 880 19104 39200 19384
rect 800 18704 39200 19104
rect 880 18424 39200 18704
rect 800 18024 39200 18424
rect 880 17744 39120 18024
rect 800 17344 39200 17744
rect 880 17064 39200 17344
rect 800 16664 39200 17064
rect 880 16384 39200 16664
rect 800 15984 39200 16384
rect 880 15704 39200 15984
rect 800 15304 39200 15704
rect 880 15024 39200 15304
rect 800 14624 39200 15024
rect 880 14344 39200 14624
rect 800 14080 39200 14344
rect 800 13944 39120 14080
rect 880 13800 39120 13944
rect 880 13664 39200 13800
rect 800 13264 39200 13664
rect 880 12984 39200 13264
rect 800 12584 39200 12984
rect 880 12304 39200 12584
rect 800 11904 39200 12304
rect 880 11624 39200 11904
rect 800 11224 39200 11624
rect 880 10944 39200 11224
rect 800 10544 39200 10944
rect 880 10264 39200 10544
rect 800 10000 39200 10264
rect 800 9864 39120 10000
rect 880 9720 39120 9864
rect 880 9584 39200 9720
rect 800 9184 39200 9584
rect 880 8904 39200 9184
rect 800 8504 39200 8904
rect 880 8224 39200 8504
rect 800 7824 39200 8224
rect 880 7544 39200 7824
rect 800 7144 39200 7544
rect 880 6864 39200 7144
rect 800 6464 39200 6864
rect 880 6184 39200 6464
rect 800 6056 39200 6184
rect 800 5784 39120 6056
rect 880 5776 39120 5784
rect 880 5504 39200 5776
rect 800 5104 39200 5504
rect 880 4824 39200 5104
rect 800 4424 39200 4824
rect 880 4144 39200 4424
rect 800 3744 39200 4144
rect 880 3464 39200 3744
rect 800 3064 39200 3464
rect 880 2784 39200 3064
rect 800 2384 39200 2784
rect 880 2112 39200 2384
rect 880 2104 39120 2112
rect 800 1832 39120 2104
rect 800 1704 39200 1832
rect 880 1424 39200 1704
rect 800 1024 39200 1424
rect 880 744 39200 1024
rect 800 480 39200 744
rect 880 307 39200 480
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal2 s 9954 39200 10010 40000 6 clk
port 1 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 peripheralBus_address[0]
port 2 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 peripheralBus_address[10]
port 3 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 peripheralBus_address[11]
port 4 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 peripheralBus_address[12]
port 5 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 peripheralBus_address[13]
port 6 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 peripheralBus_address[14]
port 7 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 peripheralBus_address[15]
port 8 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 peripheralBus_address[16]
port 9 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 peripheralBus_address[17]
port 10 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 peripheralBus_address[18]
port 11 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 peripheralBus_address[19]
port 12 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 peripheralBus_address[1]
port 13 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 peripheralBus_address[20]
port 14 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 peripheralBus_address[21]
port 15 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 peripheralBus_address[22]
port 16 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 peripheralBus_address[23]
port 17 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 peripheralBus_address[2]
port 18 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 peripheralBus_address[3]
port 19 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 peripheralBus_address[4]
port 20 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 peripheralBus_address[5]
port 21 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 peripheralBus_address[6]
port 22 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 peripheralBus_address[7]
port 23 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 peripheralBus_address[8]
port 24 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 peripheralBus_address[9]
port 25 nsew signal input
rlabel metal3 s 0 280 800 400 6 peripheralBus_busy
port 26 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 peripheralBus_data[0]
port 27 nsew signal bidirectional
rlabel metal3 s 0 16464 800 16584 6 peripheralBus_data[10]
port 28 nsew signal bidirectional
rlabel metal3 s 0 17824 800 17944 6 peripheralBus_data[11]
port 29 nsew signal bidirectional
rlabel metal3 s 0 19184 800 19304 6 peripheralBus_data[12]
port 30 nsew signal bidirectional
rlabel metal3 s 0 20544 800 20664 6 peripheralBus_data[13]
port 31 nsew signal bidirectional
rlabel metal3 s 0 21904 800 22024 6 peripheralBus_data[14]
port 32 nsew signal bidirectional
rlabel metal3 s 0 23264 800 23384 6 peripheralBus_data[15]
port 33 nsew signal bidirectional
rlabel metal3 s 0 24624 800 24744 6 peripheralBus_data[16]
port 34 nsew signal bidirectional
rlabel metal3 s 0 25984 800 26104 6 peripheralBus_data[17]
port 35 nsew signal bidirectional
rlabel metal3 s 0 27344 800 27464 6 peripheralBus_data[18]
port 36 nsew signal bidirectional
rlabel metal3 s 0 28704 800 28824 6 peripheralBus_data[19]
port 37 nsew signal bidirectional
rlabel metal3 s 0 4224 800 4344 6 peripheralBus_data[1]
port 38 nsew signal bidirectional
rlabel metal3 s 0 30064 800 30184 6 peripheralBus_data[20]
port 39 nsew signal bidirectional
rlabel metal3 s 0 31424 800 31544 6 peripheralBus_data[21]
port 40 nsew signal bidirectional
rlabel metal3 s 0 32784 800 32904 6 peripheralBus_data[22]
port 41 nsew signal bidirectional
rlabel metal3 s 0 34144 800 34264 6 peripheralBus_data[23]
port 42 nsew signal bidirectional
rlabel metal3 s 0 34824 800 34944 6 peripheralBus_data[24]
port 43 nsew signal bidirectional
rlabel metal3 s 0 35504 800 35624 6 peripheralBus_data[25]
port 44 nsew signal bidirectional
rlabel metal3 s 0 36184 800 36304 6 peripheralBus_data[26]
port 45 nsew signal bidirectional
rlabel metal3 s 0 36864 800 36984 6 peripheralBus_data[27]
port 46 nsew signal bidirectional
rlabel metal3 s 0 37544 800 37664 6 peripheralBus_data[28]
port 47 nsew signal bidirectional
rlabel metal3 s 0 38224 800 38344 6 peripheralBus_data[29]
port 48 nsew signal bidirectional
rlabel metal3 s 0 5584 800 5704 6 peripheralBus_data[2]
port 49 nsew signal bidirectional
rlabel metal3 s 0 38904 800 39024 6 peripheralBus_data[30]
port 50 nsew signal bidirectional
rlabel metal3 s 0 39584 800 39704 6 peripheralBus_data[31]
port 51 nsew signal bidirectional
rlabel metal3 s 0 6944 800 7064 6 peripheralBus_data[3]
port 52 nsew signal bidirectional
rlabel metal3 s 0 8304 800 8424 6 peripheralBus_data[4]
port 53 nsew signal bidirectional
rlabel metal3 s 0 9664 800 9784 6 peripheralBus_data[5]
port 54 nsew signal bidirectional
rlabel metal3 s 0 11024 800 11144 6 peripheralBus_data[6]
port 55 nsew signal bidirectional
rlabel metal3 s 0 12384 800 12504 6 peripheralBus_data[7]
port 56 nsew signal bidirectional
rlabel metal3 s 0 13744 800 13864 6 peripheralBus_data[8]
port 57 nsew signal bidirectional
rlabel metal3 s 0 15104 800 15224 6 peripheralBus_data[9]
port 58 nsew signal bidirectional
rlabel metal3 s 0 824 800 944 6 peripheralBus_oe
port 59 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 peripheralBus_we
port 60 nsew signal input
rlabel metal2 s 29918 39200 29974 40000 6 rst
port 61 nsew signal input
rlabel metal3 s 39200 1912 40000 2032 6 spi_clk[0]
port 62 nsew signal output
rlabel metal3 s 39200 21904 40000 22024 6 spi_clk[1]
port 63 nsew signal output
rlabel metal3 s 39200 5856 40000 5976 6 spi_cs[0]
port 64 nsew signal output
rlabel metal3 s 39200 25848 40000 25968 6 spi_cs[1]
port 65 nsew signal output
rlabel metal3 s 39200 9800 40000 9920 6 spi_en[0]
port 66 nsew signal output
rlabel metal3 s 39200 29792 40000 29912 6 spi_en[1]
port 67 nsew signal output
rlabel metal3 s 39200 13880 40000 14000 6 spi_miso[0]
port 68 nsew signal input
rlabel metal3 s 39200 33872 40000 33992 6 spi_miso[1]
port 69 nsew signal input
rlabel metal3 s 39200 17824 40000 17944 6 spi_mosi[0]
port 70 nsew signal output
rlabel metal3 s 39200 37816 40000 37936 6 spi_mosi[1]
port 71 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 72 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 72 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 73 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2495006
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_SPI/runs/Peripheral_SPI/results/finishing/SPI.magic.gds
string GDS_START 264836
<< end >>

