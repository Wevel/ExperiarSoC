magic
tech sky130A
magscale 1 2
timestamp 1654262689
<< obsli1 >>
rect 1104 2159 118864 187697
<< obsm1 >>
rect 14 1844 119218 187808
<< metal2 >>
rect 754 189200 810 190000
rect 2226 189200 2282 190000
rect 3790 189200 3846 190000
rect 5354 189200 5410 190000
rect 6918 189200 6974 190000
rect 8482 189200 8538 190000
rect 10046 189200 10102 190000
rect 11610 189200 11666 190000
rect 13174 189200 13230 190000
rect 14738 189200 14794 190000
rect 16302 189200 16358 190000
rect 17866 189200 17922 190000
rect 19430 189200 19486 190000
rect 20994 189200 21050 190000
rect 22558 189200 22614 190000
rect 24122 189200 24178 190000
rect 25594 189200 25650 190000
rect 27158 189200 27214 190000
rect 28722 189200 28778 190000
rect 30286 189200 30342 190000
rect 31850 189200 31906 190000
rect 33414 189200 33470 190000
rect 34978 189200 35034 190000
rect 36542 189200 36598 190000
rect 38106 189200 38162 190000
rect 39670 189200 39726 190000
rect 41234 189200 41290 190000
rect 42798 189200 42854 190000
rect 44362 189200 44418 190000
rect 45926 189200 45982 190000
rect 47490 189200 47546 190000
rect 48962 189200 49018 190000
rect 50526 189200 50582 190000
rect 52090 189200 52146 190000
rect 53654 189200 53710 190000
rect 55218 189200 55274 190000
rect 56782 189200 56838 190000
rect 58346 189200 58402 190000
rect 59910 189200 59966 190000
rect 61474 189200 61530 190000
rect 63038 189200 63094 190000
rect 64602 189200 64658 190000
rect 66166 189200 66222 190000
rect 67730 189200 67786 190000
rect 69294 189200 69350 190000
rect 70858 189200 70914 190000
rect 72422 189200 72478 190000
rect 73894 189200 73950 190000
rect 75458 189200 75514 190000
rect 77022 189200 77078 190000
rect 78586 189200 78642 190000
rect 80150 189200 80206 190000
rect 81714 189200 81770 190000
rect 83278 189200 83334 190000
rect 84842 189200 84898 190000
rect 86406 189200 86462 190000
rect 87970 189200 88026 190000
rect 89534 189200 89590 190000
rect 91098 189200 91154 190000
rect 92662 189200 92718 190000
rect 94226 189200 94282 190000
rect 95790 189200 95846 190000
rect 97262 189200 97318 190000
rect 98826 189200 98882 190000
rect 100390 189200 100446 190000
rect 101954 189200 102010 190000
rect 103518 189200 103574 190000
rect 105082 189200 105138 190000
rect 106646 189200 106702 190000
rect 108210 189200 108266 190000
rect 109774 189200 109830 190000
rect 111338 189200 111394 190000
rect 112902 189200 112958 190000
rect 114466 189200 114522 190000
rect 116030 189200 116086 190000
rect 117594 189200 117650 190000
rect 119158 189200 119214 190000
rect 938 0 994 800
rect 2870 0 2926 800
rect 4802 0 4858 800
rect 6826 0 6882 800
rect 8758 0 8814 800
rect 10690 0 10746 800
rect 12714 0 12770 800
rect 14646 0 14702 800
rect 16670 0 16726 800
rect 18602 0 18658 800
rect 20534 0 20590 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28446 0 28502 800
rect 30378 0 30434 800
rect 32402 0 32458 800
rect 34334 0 34390 800
rect 36266 0 36322 800
rect 38290 0 38346 800
rect 40222 0 40278 800
rect 42154 0 42210 800
rect 44178 0 44234 800
rect 46110 0 46166 800
rect 48134 0 48190 800
rect 50066 0 50122 800
rect 51998 0 52054 800
rect 54022 0 54078 800
rect 55954 0 56010 800
rect 57886 0 57942 800
rect 59910 0 59966 800
rect 61842 0 61898 800
rect 63866 0 63922 800
rect 65798 0 65854 800
rect 67730 0 67786 800
rect 69754 0 69810 800
rect 71686 0 71742 800
rect 73618 0 73674 800
rect 75642 0 75698 800
rect 77574 0 77630 800
rect 79598 0 79654 800
rect 81530 0 81586 800
rect 83462 0 83518 800
rect 85486 0 85542 800
rect 87418 0 87474 800
rect 89350 0 89406 800
rect 91374 0 91430 800
rect 93306 0 93362 800
rect 95330 0 95386 800
rect 97262 0 97318 800
rect 99194 0 99250 800
rect 101218 0 101274 800
rect 103150 0 103206 800
rect 105082 0 105138 800
rect 107106 0 107162 800
rect 109038 0 109094 800
rect 111062 0 111118 800
rect 112994 0 113050 800
rect 114926 0 114982 800
rect 116950 0 117006 800
rect 118882 0 118938 800
<< obsm2 >>
rect 20 189144 698 189258
rect 866 189144 2170 189258
rect 2338 189144 3734 189258
rect 3902 189144 5298 189258
rect 5466 189144 6862 189258
rect 7030 189144 8426 189258
rect 8594 189144 9990 189258
rect 10158 189144 11554 189258
rect 11722 189144 13118 189258
rect 13286 189144 14682 189258
rect 14850 189144 16246 189258
rect 16414 189144 17810 189258
rect 17978 189144 19374 189258
rect 19542 189144 20938 189258
rect 21106 189144 22502 189258
rect 22670 189144 24066 189258
rect 24234 189144 25538 189258
rect 25706 189144 27102 189258
rect 27270 189144 28666 189258
rect 28834 189144 30230 189258
rect 30398 189144 31794 189258
rect 31962 189144 33358 189258
rect 33526 189144 34922 189258
rect 35090 189144 36486 189258
rect 36654 189144 38050 189258
rect 38218 189144 39614 189258
rect 39782 189144 41178 189258
rect 41346 189144 42742 189258
rect 42910 189144 44306 189258
rect 44474 189144 45870 189258
rect 46038 189144 47434 189258
rect 47602 189144 48906 189258
rect 49074 189144 50470 189258
rect 50638 189144 52034 189258
rect 52202 189144 53598 189258
rect 53766 189144 55162 189258
rect 55330 189144 56726 189258
rect 56894 189144 58290 189258
rect 58458 189144 59854 189258
rect 60022 189144 61418 189258
rect 61586 189144 62982 189258
rect 63150 189144 64546 189258
rect 64714 189144 66110 189258
rect 66278 189144 67674 189258
rect 67842 189144 69238 189258
rect 69406 189144 70802 189258
rect 70970 189144 72366 189258
rect 72534 189144 73838 189258
rect 74006 189144 75402 189258
rect 75570 189144 76966 189258
rect 77134 189144 78530 189258
rect 78698 189144 80094 189258
rect 80262 189144 81658 189258
rect 81826 189144 83222 189258
rect 83390 189144 84786 189258
rect 84954 189144 86350 189258
rect 86518 189144 87914 189258
rect 88082 189144 89478 189258
rect 89646 189144 91042 189258
rect 91210 189144 92606 189258
rect 92774 189144 94170 189258
rect 94338 189144 95734 189258
rect 95902 189144 97206 189258
rect 97374 189144 98770 189258
rect 98938 189144 100334 189258
rect 100502 189144 101898 189258
rect 102066 189144 103462 189258
rect 103630 189144 105026 189258
rect 105194 189144 106590 189258
rect 106758 189144 108154 189258
rect 108322 189144 109718 189258
rect 109886 189144 111282 189258
rect 111450 189144 112846 189258
rect 113014 189144 114410 189258
rect 114578 189144 115974 189258
rect 116142 189144 117538 189258
rect 117706 189144 119102 189258
rect 20 856 119212 189144
rect 20 800 882 856
rect 1050 800 2814 856
rect 2982 800 4746 856
rect 4914 800 6770 856
rect 6938 800 8702 856
rect 8870 800 10634 856
rect 10802 800 12658 856
rect 12826 800 14590 856
rect 14758 800 16614 856
rect 16782 800 18546 856
rect 18714 800 20478 856
rect 20646 800 22502 856
rect 22670 800 24434 856
rect 24602 800 26366 856
rect 26534 800 28390 856
rect 28558 800 30322 856
rect 30490 800 32346 856
rect 32514 800 34278 856
rect 34446 800 36210 856
rect 36378 800 38234 856
rect 38402 800 40166 856
rect 40334 800 42098 856
rect 42266 800 44122 856
rect 44290 800 46054 856
rect 46222 800 48078 856
rect 48246 800 50010 856
rect 50178 800 51942 856
rect 52110 800 53966 856
rect 54134 800 55898 856
rect 56066 800 57830 856
rect 57998 800 59854 856
rect 60022 800 61786 856
rect 61954 800 63810 856
rect 63978 800 65742 856
rect 65910 800 67674 856
rect 67842 800 69698 856
rect 69866 800 71630 856
rect 71798 800 73562 856
rect 73730 800 75586 856
rect 75754 800 77518 856
rect 77686 800 79542 856
rect 79710 800 81474 856
rect 81642 800 83406 856
rect 83574 800 85430 856
rect 85598 800 87362 856
rect 87530 800 89294 856
rect 89462 800 91318 856
rect 91486 800 93250 856
rect 93418 800 95274 856
rect 95442 800 97206 856
rect 97374 800 99138 856
rect 99306 800 101162 856
rect 101330 800 103094 856
rect 103262 800 105026 856
rect 105194 800 107050 856
rect 107218 800 108982 856
rect 109150 800 111006 856
rect 111174 800 112938 856
rect 113106 800 114870 856
rect 115038 800 116894 856
rect 117062 800 118826 856
rect 118994 800 119212 856
<< metal3 >>
rect 0 188912 800 189032
rect 0 187144 800 187264
rect 0 185240 800 185360
rect 0 183472 800 183592
rect 0 181568 800 181688
rect 0 179800 800 179920
rect 0 177896 800 178016
rect 0 176128 800 176248
rect 0 174360 800 174480
rect 119200 174088 120000 174208
rect 0 172456 800 172576
rect 0 170688 800 170808
rect 0 168784 800 168904
rect 0 167016 800 167136
rect 0 165112 800 165232
rect 0 163344 800 163464
rect 0 161576 800 161696
rect 0 159672 800 159792
rect 0 157904 800 158024
rect 0 156000 800 156120
rect 0 154232 800 154352
rect 0 152328 800 152448
rect 0 150560 800 150680
rect 0 148792 800 148912
rect 0 146888 800 147008
rect 0 145120 800 145240
rect 0 143216 800 143336
rect 119200 142400 120000 142520
rect 0 141448 800 141568
rect 0 139544 800 139664
rect 0 137776 800 137896
rect 0 136008 800 136128
rect 0 134104 800 134224
rect 0 132336 800 132456
rect 0 130432 800 130552
rect 0 128664 800 128784
rect 0 126760 800 126880
rect 0 124992 800 125112
rect 0 123088 800 123208
rect 0 121320 800 121440
rect 0 119552 800 119672
rect 0 117648 800 117768
rect 0 115880 800 116000
rect 0 113976 800 114096
rect 0 112208 800 112328
rect 119200 110712 120000 110832
rect 0 110304 800 110424
rect 0 108536 800 108656
rect 0 106768 800 106888
rect 0 104864 800 104984
rect 0 103096 800 103216
rect 0 101192 800 101312
rect 0 99424 800 99544
rect 0 97520 800 97640
rect 0 95752 800 95872
rect 0 93984 800 94104
rect 0 92080 800 92200
rect 0 90312 800 90432
rect 0 88408 800 88528
rect 0 86640 800 86760
rect 0 84736 800 84856
rect 0 82968 800 83088
rect 0 81200 800 81320
rect 0 79296 800 79416
rect 119200 79024 120000 79144
rect 0 77528 800 77648
rect 0 75624 800 75744
rect 0 73856 800 73976
rect 0 71952 800 72072
rect 0 70184 800 70304
rect 0 68416 800 68536
rect 0 66512 800 66632
rect 0 64744 800 64864
rect 0 62840 800 62960
rect 0 61072 800 61192
rect 0 59168 800 59288
rect 0 57400 800 57520
rect 0 55496 800 55616
rect 0 53728 800 53848
rect 0 51960 800 52080
rect 0 50056 800 50176
rect 0 48288 800 48408
rect 119200 47336 120000 47456
rect 0 46384 800 46504
rect 0 44616 800 44736
rect 0 42712 800 42832
rect 0 40944 800 41064
rect 0 39176 800 39296
rect 0 37272 800 37392
rect 0 35504 800 35624
rect 0 33600 800 33720
rect 0 31832 800 31952
rect 0 29928 800 30048
rect 0 28160 800 28280
rect 0 26392 800 26512
rect 0 24488 800 24608
rect 0 22720 800 22840
rect 0 20816 800 20936
rect 0 19048 800 19168
rect 0 17144 800 17264
rect 119200 15784 120000 15904
rect 0 15376 800 15496
rect 0 13608 800 13728
rect 0 11704 800 11824
rect 0 9936 800 10056
rect 0 8032 800 8152
rect 0 6264 800 6384
rect 0 4360 800 4480
rect 0 2592 800 2712
rect 0 824 800 944
<< obsm3 >>
rect 880 188832 119200 189005
rect 800 187344 119200 188832
rect 880 187064 119200 187344
rect 800 185440 119200 187064
rect 880 185160 119200 185440
rect 800 183672 119200 185160
rect 880 183392 119200 183672
rect 800 181768 119200 183392
rect 880 181488 119200 181768
rect 800 180000 119200 181488
rect 880 179720 119200 180000
rect 800 178096 119200 179720
rect 880 177816 119200 178096
rect 800 176328 119200 177816
rect 880 176048 119200 176328
rect 800 174560 119200 176048
rect 880 174288 119200 174560
rect 880 174280 119120 174288
rect 800 174008 119120 174280
rect 800 172656 119200 174008
rect 880 172376 119200 172656
rect 800 170888 119200 172376
rect 880 170608 119200 170888
rect 800 168984 119200 170608
rect 880 168704 119200 168984
rect 800 167216 119200 168704
rect 880 166936 119200 167216
rect 800 165312 119200 166936
rect 880 165032 119200 165312
rect 800 163544 119200 165032
rect 880 163264 119200 163544
rect 800 161776 119200 163264
rect 880 161496 119200 161776
rect 800 159872 119200 161496
rect 880 159592 119200 159872
rect 800 158104 119200 159592
rect 880 157824 119200 158104
rect 800 156200 119200 157824
rect 880 155920 119200 156200
rect 800 154432 119200 155920
rect 880 154152 119200 154432
rect 800 152528 119200 154152
rect 880 152248 119200 152528
rect 800 150760 119200 152248
rect 880 150480 119200 150760
rect 800 148992 119200 150480
rect 880 148712 119200 148992
rect 800 147088 119200 148712
rect 880 146808 119200 147088
rect 800 145320 119200 146808
rect 880 145040 119200 145320
rect 800 143416 119200 145040
rect 880 143136 119200 143416
rect 800 142600 119200 143136
rect 800 142320 119120 142600
rect 800 141648 119200 142320
rect 880 141368 119200 141648
rect 800 139744 119200 141368
rect 880 139464 119200 139744
rect 800 137976 119200 139464
rect 880 137696 119200 137976
rect 800 136208 119200 137696
rect 880 135928 119200 136208
rect 800 134304 119200 135928
rect 880 134024 119200 134304
rect 800 132536 119200 134024
rect 880 132256 119200 132536
rect 800 130632 119200 132256
rect 880 130352 119200 130632
rect 800 128864 119200 130352
rect 880 128584 119200 128864
rect 800 126960 119200 128584
rect 880 126680 119200 126960
rect 800 125192 119200 126680
rect 880 124912 119200 125192
rect 800 123288 119200 124912
rect 880 123008 119200 123288
rect 800 121520 119200 123008
rect 880 121240 119200 121520
rect 800 119752 119200 121240
rect 880 119472 119200 119752
rect 800 117848 119200 119472
rect 880 117568 119200 117848
rect 800 116080 119200 117568
rect 880 115800 119200 116080
rect 800 114176 119200 115800
rect 880 113896 119200 114176
rect 800 112408 119200 113896
rect 880 112128 119200 112408
rect 800 110912 119200 112128
rect 800 110632 119120 110912
rect 800 110504 119200 110632
rect 880 110224 119200 110504
rect 800 108736 119200 110224
rect 880 108456 119200 108736
rect 800 106968 119200 108456
rect 880 106688 119200 106968
rect 800 105064 119200 106688
rect 880 104784 119200 105064
rect 800 103296 119200 104784
rect 880 103016 119200 103296
rect 800 101392 119200 103016
rect 880 101112 119200 101392
rect 800 99624 119200 101112
rect 880 99344 119200 99624
rect 800 97720 119200 99344
rect 880 97440 119200 97720
rect 800 95952 119200 97440
rect 880 95672 119200 95952
rect 800 94184 119200 95672
rect 880 93904 119200 94184
rect 800 92280 119200 93904
rect 880 92000 119200 92280
rect 800 90512 119200 92000
rect 880 90232 119200 90512
rect 800 88608 119200 90232
rect 880 88328 119200 88608
rect 800 86840 119200 88328
rect 880 86560 119200 86840
rect 800 84936 119200 86560
rect 880 84656 119200 84936
rect 800 83168 119200 84656
rect 880 82888 119200 83168
rect 800 81400 119200 82888
rect 880 81120 119200 81400
rect 800 79496 119200 81120
rect 880 79224 119200 79496
rect 880 79216 119120 79224
rect 800 78944 119120 79216
rect 800 77728 119200 78944
rect 880 77448 119200 77728
rect 800 75824 119200 77448
rect 880 75544 119200 75824
rect 800 74056 119200 75544
rect 880 73776 119200 74056
rect 800 72152 119200 73776
rect 880 71872 119200 72152
rect 800 70384 119200 71872
rect 880 70104 119200 70384
rect 800 68616 119200 70104
rect 880 68336 119200 68616
rect 800 66712 119200 68336
rect 880 66432 119200 66712
rect 800 64944 119200 66432
rect 880 64664 119200 64944
rect 800 63040 119200 64664
rect 880 62760 119200 63040
rect 800 61272 119200 62760
rect 880 60992 119200 61272
rect 800 59368 119200 60992
rect 880 59088 119200 59368
rect 800 57600 119200 59088
rect 880 57320 119200 57600
rect 800 55696 119200 57320
rect 880 55416 119200 55696
rect 800 53928 119200 55416
rect 880 53648 119200 53928
rect 800 52160 119200 53648
rect 880 51880 119200 52160
rect 800 50256 119200 51880
rect 880 49976 119200 50256
rect 800 48488 119200 49976
rect 880 48208 119200 48488
rect 800 47536 119200 48208
rect 800 47256 119120 47536
rect 800 46584 119200 47256
rect 880 46304 119200 46584
rect 800 44816 119200 46304
rect 880 44536 119200 44816
rect 800 42912 119200 44536
rect 880 42632 119200 42912
rect 800 41144 119200 42632
rect 880 40864 119200 41144
rect 800 39376 119200 40864
rect 880 39096 119200 39376
rect 800 37472 119200 39096
rect 880 37192 119200 37472
rect 800 35704 119200 37192
rect 880 35424 119200 35704
rect 800 33800 119200 35424
rect 880 33520 119200 33800
rect 800 32032 119200 33520
rect 880 31752 119200 32032
rect 800 30128 119200 31752
rect 880 29848 119200 30128
rect 800 28360 119200 29848
rect 880 28080 119200 28360
rect 800 26592 119200 28080
rect 880 26312 119200 26592
rect 800 24688 119200 26312
rect 880 24408 119200 24688
rect 800 22920 119200 24408
rect 880 22640 119200 22920
rect 800 21016 119200 22640
rect 880 20736 119200 21016
rect 800 19248 119200 20736
rect 880 18968 119200 19248
rect 800 17344 119200 18968
rect 880 17064 119200 17344
rect 800 15984 119200 17064
rect 800 15704 119120 15984
rect 800 15576 119200 15704
rect 880 15296 119200 15576
rect 800 13808 119200 15296
rect 880 13528 119200 13808
rect 800 11904 119200 13528
rect 880 11624 119200 11904
rect 800 10136 119200 11624
rect 880 9856 119200 10136
rect 800 8232 119200 9856
rect 880 7952 119200 8232
rect 800 6464 119200 7952
rect 880 6184 119200 6464
rect 800 4560 119200 6184
rect 880 4280 119200 4560
rect 800 2792 119200 4280
rect 880 2512 119200 2792
rect 800 1024 119200 2512
rect 880 851 119200 1024
<< metal4 >>
rect 4208 2128 4528 187728
rect 19568 2128 19888 187728
rect 34928 2128 35248 187728
rect 50288 2128 50608 187728
rect 65648 2128 65968 187728
rect 81008 2128 81328 187728
rect 96368 2128 96688 187728
rect 111728 2128 112048 187728
<< obsm4 >>
rect 1899 2619 4128 186829
rect 4608 2619 19488 186829
rect 19968 2619 34848 186829
rect 35328 2619 50208 186829
rect 50688 2619 65568 186829
rect 66048 2619 80928 186829
rect 81408 2619 96288 186829
rect 96768 2619 111648 186829
rect 112128 2619 116045 186829
<< labels >>
rlabel metal2 s 79598 0 79654 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 754 189200 810 190000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 16302 189200 16358 190000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 17866 189200 17922 190000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 19430 189200 19486 190000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 20994 189200 21050 190000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 22558 189200 22614 190000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 24122 189200 24178 190000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 25594 189200 25650 190000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 27158 189200 27214 190000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 28722 189200 28778 190000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 30286 189200 30342 190000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2226 189200 2282 190000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 31850 189200 31906 190000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 33414 189200 33470 190000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 34978 189200 35034 190000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 36542 189200 36598 190000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 38106 189200 38162 190000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 39670 189200 39726 190000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 41234 189200 41290 190000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 42798 189200 42854 190000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 44362 189200 44418 190000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 45926 189200 45982 190000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 3790 189200 3846 190000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 47490 189200 47546 190000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 48962 189200 49018 190000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 50526 189200 50582 190000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 52090 189200 52146 190000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 53654 189200 53710 190000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 55218 189200 55274 190000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 56782 189200 56838 190000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 58346 189200 58402 190000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 5354 189200 5410 190000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 6918 189200 6974 190000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 8482 189200 8538 190000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 10046 189200 10102 190000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 11610 189200 11666 190000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 13174 189200 13230 190000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 14738 189200 14794 190000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 938 0 994 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 59910 189200 59966 190000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 75458 189200 75514 190000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 77022 189200 77078 190000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 78586 189200 78642 190000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 80150 189200 80206 190000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 81714 189200 81770 190000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 83278 189200 83334 190000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 84842 189200 84898 190000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 86406 189200 86462 190000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 87970 189200 88026 190000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 89534 189200 89590 190000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 61474 189200 61530 190000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 91098 189200 91154 190000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 92662 189200 92718 190000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 94226 189200 94282 190000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 95790 189200 95846 190000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 97262 189200 97318 190000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 98826 189200 98882 190000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 100390 189200 100446 190000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 101954 189200 102010 190000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 103518 189200 103574 190000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 105082 189200 105138 190000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 63038 189200 63094 190000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 106646 189200 106702 190000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 108210 189200 108266 190000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 109774 189200 109830 190000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 111338 189200 111394 190000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 112902 189200 112958 190000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 114466 189200 114522 190000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 116030 189200 116086 190000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 117594 189200 117650 190000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 64602 189200 64658 190000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 66166 189200 66222 190000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 67730 189200 67786 190000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 69294 189200 69350 190000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 70858 189200 70914 190000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 72422 189200 72478 190000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 73894 189200 73950 190000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 79024 120000 79144 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 110712 120000 110832 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 142400 120000 142520 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 174088 120000 174208 6 jtag_tms
port 128 nsew signal output
rlabel metal2 s 119158 189200 119214 190000 6 peripheral_irq[0]
port 129 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 peripheral_irq[1]
port 130 nsew signal output
rlabel metal3 s 0 183472 800 183592 6 peripheral_irq[2]
port 131 nsew signal output
rlabel metal3 s 0 185240 800 185360 6 peripheral_irq[3]
port 132 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 peripheral_irq[4]
port 133 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 peripheral_irq[5]
port 134 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 peripheral_irq[6]
port 135 nsew signal output
rlabel metal3 s 0 187144 800 187264 6 peripheral_irq[7]
port 136 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 peripheral_irq[8]
port 137 nsew signal output
rlabel metal3 s 0 188912 800 189032 6 peripheral_irq[9]
port 138 nsew signal output
rlabel metal3 s 119200 15784 120000 15904 6 probe_blink[0]
port 139 nsew signal output
rlabel metal3 s 119200 47336 120000 47456 6 probe_blink[1]
port 140 nsew signal output
rlabel metal4 s 4208 2128 4528 187728 6 vccd1
port 141 nsew power input
rlabel metal4 s 34928 2128 35248 187728 6 vccd1
port 141 nsew power input
rlabel metal4 s 65648 2128 65968 187728 6 vccd1
port 141 nsew power input
rlabel metal4 s 96368 2128 96688 187728 6 vccd1
port 141 nsew power input
rlabel metal2 s 99194 0 99250 800 6 vga_b[0]
port 142 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 vga_b[1]
port 143 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 vga_g[0]
port 144 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 vga_g[1]
port 145 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 vga_hsync
port 146 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 vga_r[0]
port 147 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 vga_r[1]
port 148 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 vga_vsync
port 149 nsew signal input
rlabel metal4 s 19568 2128 19888 187728 6 vssd1
port 150 nsew ground input
rlabel metal4 s 50288 2128 50608 187728 6 vssd1
port 150 nsew ground input
rlabel metal4 s 81008 2128 81328 187728 6 vssd1
port 150 nsew ground input
rlabel metal4 s 111728 2128 112048 187728 6 vssd1
port 150 nsew ground input
rlabel metal3 s 0 824 800 944 6 wb_ack_o
port 151 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 wb_adr_i[0]
port 152 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wb_adr_i[10]
port 153 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 wb_adr_i[11]
port 154 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 wb_adr_i[12]
port 155 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 wb_adr_i[13]
port 156 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 wb_adr_i[14]
port 157 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 wb_adr_i[15]
port 158 nsew signal input
rlabel metal3 s 0 110304 800 110424 6 wb_adr_i[16]
port 159 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 wb_adr_i[17]
port 160 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 wb_adr_i[18]
port 161 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 wb_adr_i[19]
port 162 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[1]
port 163 nsew signal input
rlabel metal3 s 0 132336 800 132456 6 wb_adr_i[20]
port 164 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 wb_adr_i[21]
port 165 nsew signal input
rlabel metal3 s 0 143216 800 143336 6 wb_adr_i[22]
port 166 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 wb_adr_i[23]
port 167 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 wb_adr_i[2]
port 168 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 wb_adr_i[3]
port 169 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 wb_adr_i[4]
port 170 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 wb_adr_i[5]
port 171 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 wb_adr_i[6]
port 172 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 wb_adr_i[7]
port 173 nsew signal input
rlabel metal3 s 0 66512 800 66632 6 wb_adr_i[8]
port 174 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wb_adr_i[9]
port 175 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wb_clk_i
port 176 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wb_cyc_i
port 177 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wb_data_i[0]
port 178 nsew signal input
rlabel metal3 s 0 79296 800 79416 6 wb_data_i[10]
port 179 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 wb_data_i[11]
port 180 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 wb_data_i[12]
port 181 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 wb_data_i[13]
port 182 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 wb_data_i[14]
port 183 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 wb_data_i[15]
port 184 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 wb_data_i[16]
port 185 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 wb_data_i[17]
port 186 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 wb_data_i[18]
port 187 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 wb_data_i[19]
port 188 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[1]
port 189 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 wb_data_i[20]
port 190 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 wb_data_i[21]
port 191 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 wb_data_i[22]
port 192 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 wb_data_i[23]
port 193 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 wb_data_i[24]
port 194 nsew signal input
rlabel metal3 s 0 157904 800 158024 6 wb_data_i[25]
port 195 nsew signal input
rlabel metal3 s 0 161576 800 161696 6 wb_data_i[26]
port 196 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 wb_data_i[27]
port 197 nsew signal input
rlabel metal3 s 0 168784 800 168904 6 wb_data_i[28]
port 198 nsew signal input
rlabel metal3 s 0 172456 800 172576 6 wb_data_i[29]
port 199 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 wb_data_i[2]
port 200 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 wb_data_i[30]
port 201 nsew signal input
rlabel metal3 s 0 179800 800 179920 6 wb_data_i[31]
port 202 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 wb_data_i[3]
port 203 nsew signal input
rlabel metal3 s 0 46384 800 46504 6 wb_data_i[4]
port 204 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 wb_data_i[5]
port 205 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 wb_data_i[6]
port 206 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 wb_data_i[7]
port 207 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 wb_data_i[8]
port 208 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 wb_data_i[9]
port 209 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_data_o[0]
port 210 nsew signal output
rlabel metal3 s 0 81200 800 81320 6 wb_data_o[10]
port 211 nsew signal output
rlabel metal3 s 0 86640 800 86760 6 wb_data_o[11]
port 212 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 wb_data_o[12]
port 213 nsew signal output
rlabel metal3 s 0 97520 800 97640 6 wb_data_o[13]
port 214 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 wb_data_o[14]
port 215 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 wb_data_o[15]
port 216 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 wb_data_o[16]
port 217 nsew signal output
rlabel metal3 s 0 119552 800 119672 6 wb_data_o[17]
port 218 nsew signal output
rlabel metal3 s 0 124992 800 125112 6 wb_data_o[18]
port 219 nsew signal output
rlabel metal3 s 0 130432 800 130552 6 wb_data_o[19]
port 220 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 wb_data_o[1]
port 221 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 wb_data_o[20]
port 222 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 wb_data_o[21]
port 223 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 wb_data_o[22]
port 224 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 wb_data_o[23]
port 225 nsew signal output
rlabel metal3 s 0 156000 800 156120 6 wb_data_o[24]
port 226 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 wb_data_o[25]
port 227 nsew signal output
rlabel metal3 s 0 163344 800 163464 6 wb_data_o[26]
port 228 nsew signal output
rlabel metal3 s 0 167016 800 167136 6 wb_data_o[27]
port 229 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 wb_data_o[28]
port 230 nsew signal output
rlabel metal3 s 0 174360 800 174480 6 wb_data_o[29]
port 231 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 wb_data_o[2]
port 232 nsew signal output
rlabel metal3 s 0 177896 800 178016 6 wb_data_o[30]
port 233 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 wb_data_o[31]
port 234 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 wb_data_o[3]
port 235 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 wb_data_o[4]
port 236 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 wb_data_o[5]
port 237 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 wb_data_o[6]
port 238 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 wb_data_o[7]
port 239 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 wb_data_o[8]
port 240 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 wb_data_o[9]
port 241 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 wb_error_o
port 242 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 wb_rst_i
port 243 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 wb_sel_i[0]
port 244 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 wb_sel_i[1]
port 245 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 wb_sel_i[2]
port 246 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 wb_sel_i[3]
port 247 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 wb_stall_o
port 248 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 wb_stb_i
port 249 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wb_we_i
port 250 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 190000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 68718910
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/finishing/Peripherals.magic.gds
string GDS_START 1263966
<< end >>

